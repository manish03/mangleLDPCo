//`include "GF2_LDPC_fgallag_0x0000e_assign_inc.sv"
//always_comb begin
              I9d96959b6b7fd9b9e978d3f23959e9e1['h00000] = 
          (!fgallag_sel['h0000e]) ? 
                       I1f3af771a6bf6da6d9e448fb87a2d186['h00000] : //%
                       I1f3af771a6bf6da6d9e448fb87a2d186['h00001] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00001] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00002] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00002] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00004] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00003] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00006] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00004] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00008] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00005] =  I1f3af771a6bf6da6d9e448fb87a2d186['h0000a] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00006] =  I1f3af771a6bf6da6d9e448fb87a2d186['h0000c] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00007] =  I1f3af771a6bf6da6d9e448fb87a2d186['h0000e] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00008] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00010] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h00009] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00012] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h0000a] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00014] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h0000b] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00016] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h0000c] =  I1f3af771a6bf6da6d9e448fb87a2d186['h00018] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h0000d] =  I1f3af771a6bf6da6d9e448fb87a2d186['h0001a] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h0000e] =  I1f3af771a6bf6da6d9e448fb87a2d186['h0001c] ;
//end
//always_comb begin // 
               I9d96959b6b7fd9b9e978d3f23959e9e1['h0000f] =  I1f3af771a6bf6da6d9e448fb87a2d186['h0001e] ;
//end
