 reg  ['h7f:0] [$clog2('h7000+1)-1:0] Ibbc4b022828a232d4b3d3eccc478fd3f ;
