 reg  ['h1fff:0] [$clog2('h7000+1)-1:0] Ifcca41d795dde8a35d1654b9520c92e7 ;
