//`include "GF2_LDPC_fgallag_0x0000f_assign_inc.sv"
//always_comb begin
              Ice223344c1d41676e20d7b2668ccff71['h00000] = 
          (!fgallag_sel['h0000f]) ? 
                       I9d96959b6b7fd9b9e978d3f23959e9e1['h00000] : //%
                       I9d96959b6b7fd9b9e978d3f23959e9e1['h00001] ;
//end
//always_comb begin // 
               Ice223344c1d41676e20d7b2668ccff71['h00001] =  I9d96959b6b7fd9b9e978d3f23959e9e1['h00002] ;
//end
//always_comb begin // 
               Ice223344c1d41676e20d7b2668ccff71['h00002] =  I9d96959b6b7fd9b9e978d3f23959e9e1['h00004] ;
//end
//always_comb begin // 
               Ice223344c1d41676e20d7b2668ccff71['h00003] =  I9d96959b6b7fd9b9e978d3f23959e9e1['h00006] ;
//end
//always_comb begin // 
               Ice223344c1d41676e20d7b2668ccff71['h00004] =  I9d96959b6b7fd9b9e978d3f23959e9e1['h00008] ;
//end
//always_comb begin // 
               Ice223344c1d41676e20d7b2668ccff71['h00005] =  I9d96959b6b7fd9b9e978d3f23959e9e1['h0000a] ;
//end
//always_comb begin // 
               Ice223344c1d41676e20d7b2668ccff71['h00006] =  I9d96959b6b7fd9b9e978d3f23959e9e1['h0000c] ;
//end
//always_comb begin // 
               Ice223344c1d41676e20d7b2668ccff71['h00007] =  I9d96959b6b7fd9b9e978d3f23959e9e1['h0000e] ;
//end
