 reg  ['h1:0] [$clog2('h7000+1)-1:0] I34f69b29975fc71eeee92e6ac4210723 ;
