              I480377e3a6fbaf775422573d801193be = 
          (!flogtanh_sel[5]) ? 
                       I148a2b6bf6253f900182125f4f086010: 
                       I23d8325c203e2a9e4118ea94210effa0;
              I21550e4abf93f66dbb624e2fa12724ae = 
          (!flogtanh_sel[5]) ? 
                       I9cdc23307c28dd846a7981b6a1b8552e: 
                       I2b9e2a2b9bea3cdd0c7b48f864254aa8;
              I1399556483c51f8d866cc756d4d485f5 = 
          (!flogtanh_sel[5]) ? 
                       I0da340314517b5042829528ed7621d8f: 
                       I4edefd1be2348543f0e11dbce5623271;
              I98c3b475d2c5967e0fea09dd872baf38 = 
          (!flogtanh_sel[5]) ? 
                       I8315a1e97dcb0458031c17b029afac99: 
                       I2b91900229ffbdfcd6ff7f127546ea17;
              I7850d8a8e92d9764f664675c922eca89 = 
          (!flogtanh_sel[5]) ? 
                       I551b47851eee1b096612760b461e8207: 
                       I273b2b9c28034900d30631a61f1aecc7;
              Ib55eb35fe60a4878bffecac46af4d0d6 = 
          (!flogtanh_sel[5]) ? 
                       I641d4634620bb210a64564be02fa920f: 
                       Ib0f8bb863f94f35f2c880323f8793565;
