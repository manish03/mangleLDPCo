`include "fgallag/GF2_LDPC_fgallag.sv.1"
`include "fgallag/GF2_LDPC_fgallag.sv.2"
