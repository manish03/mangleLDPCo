//`include "GF2_LDPC_fgallag_0x00011_assign_inc.sv"
//always_comb begin
              Id639acb3a3eafcec248bdf33943866f07fefacf8e1d90896c6a07bb83a1177a8['h00000] = 
          (!fgallag_sel['h00011]) ? 
                       Ia5096e066539b84a69d699a447597782df45e307c461c4dec11d6ed88887b470['h00000] : //%
                       Ia5096e066539b84a69d699a447597782df45e307c461c4dec11d6ed88887b470['h00001] ;
//end
//always_comb begin // 
               Id639acb3a3eafcec248bdf33943866f07fefacf8e1d90896c6a07bb83a1177a8['h00001] =  Ia5096e066539b84a69d699a447597782df45e307c461c4dec11d6ed88887b470['h00002] ;
//end
