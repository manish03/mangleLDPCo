 reg  ['h3ffff:0] [$clog2('h7000+1)-1:0] Ic8af899784d96b1bcae05a6728ce00582b2cfa841431ae64ece6892ed315cb91 ;
