reg [fgallag_WDTH -1:0] Ib215a1b985e00121a1c48cf2ddae939a, I2e449260cbba5283dbe9d183eaa3006b;
reg [fgallag_WDTH -1:0] I0d9537bea5895773b487fb385690c92c, Ie43af039b1e5b11fe91210b644a1a31e;
reg [fgallag_WDTH -1:0] I287708a4c364df837b06049357518409, Iebddca10e7f7c3688d5011f147ffcd4a;
reg [fgallag_WDTH -1:0] I9e69bf6d258b709d9706052822d9ae16, I93b9a635a3e05192ad53b6e264275aa9;
reg [fgallag_WDTH -1:0] I0d187ebb6dbedda971b33ceebb6f17eb, Ie3012c652b244e53fc44455982b5eefa;
reg [fgallag_WDTH -1:0] I83ab1426707044dca3ed926493081311, Ie287c2f7d9779d50be27d3d5a9de6a33;
reg [fgallag_WDTH -1:0] Ib402ea81f3ba6d26feac26905f0c5edc, Ia9327a6a37a1de7dbf3839eafb5d941e;
reg [fgallag_WDTH -1:0] I457501e8372fe81287f139beeaad0452, I47705f99ef5cb6172811f4046484597c;
reg [fgallag_WDTH -1:0] I6f3ecf6c401215c1242c6d31cb4158d7, Ie1c96dc77190cd04130a400e869a5abd;
reg [fgallag_WDTH -1:0] Ia439d59ddaa34c9a8dec425ac4f7aca1, Iafcc3b17af5dbd70300172c2e2742206;
reg [fgallag_WDTH -1:0] I11a9a93502a123a616205de5969bd5c8, I47731679e4d0f87f9d19934c25f2bdcb;
reg [fgallag_WDTH -1:0] I346c6ffdb07c9d7a5939fcd142871ef8, I9608c445e266884a86508e3ea3a53853;
reg [fgallag_WDTH -1:0] I20fa0bb8e0dc75902328a349f0dca139, I0fb3749641e7b5675524cd796ef4127c;
reg [fgallag_WDTH -1:0] Idb4bf6de8f078619ea6dcb51d8f7d329, Id5b6b690dc055c374a44fb1ecfd54198;
reg [fgallag_WDTH -1:0] I8d2f1e18f0064f50176caa84061bf7ec, I6ae44809304b38046cc0afb4317a3f43;
reg [fgallag_WDTH -1:0] Ic48ab17819fe5de2326e4fcb0a1e84c2, I3ef49ef515a84b68f7bff1fbc0f05be7;
reg [fgallag_WDTH -1:0] If7332a4a9a6924d2fcbd0af70ecc0d1b, I62939bc5509a6ca4278bedb7be3f4534;
reg [fgallag_WDTH -1:0] I65a8d4181ad1817636600b816f41158b, Ieaaab9e41c6a940e06ce877c3e6faebc;
reg [fgallag_WDTH -1:0] I746285d851cff1339ce0b99930415c2b, Iadf3bdeaff4bc193443ef22aef0ad7b7;
reg [fgallag_WDTH -1:0] I3305daafd6c3dc6ceb95673b361f0480, Ic65a2079483506c24674715cc402a81b;
reg [fgallag_WDTH -1:0] I68babd78d3c2b1d6a064b25a3abd690e, Ia7641d441a79bfea63ba407052928bc5;
reg [fgallag_WDTH -1:0] I9e7d989a414d752920fd69ac7c23ca38, I299c542d09419d0998b59bf1f184a78a;
reg [fgallag_WDTH -1:0] Ibf1b1639efba4277e759d747abe85e6b, I8aa5ad4f2f437be64a88554e6dfc3c6b;
reg [fgallag_WDTH -1:0] If67570ab71fa30823c9fe1277f35c1fe, Iaf0980a21e4ee5e842a5b6db664264f6;
reg [fgallag_WDTH -1:0] Ia660cf2aa760392654bbc61cb60d9920, I80df82d24c9507274353efb085b46fda;
reg [fgallag_WDTH -1:0] I2bf7c2dabc30d2207f04e0f6970f2287, I1db5a382bb7c2317716c3137fd10d07c;
reg [fgallag_WDTH -1:0] I75c6cf6f3378e1377047d467a7e827f7, Icb748243d2a5f8cc86c44566e1732232;
reg [fgallag_WDTH -1:0] Ic3dacf077252960c863e8ec1a880f313, I90a0c6bd80d2357d7b865f61a18ae13b;
reg [fgallag_WDTH -1:0] I781a85002cfeb3038120fe37047710bc, I16af13e02ee36dbcdeab785596175a3c;
reg [fgallag_WDTH -1:0] I0e8936dc5acf0e7c165d76a8b58f2765, Id0e47470fba20bc467a05d0dd09bf560;
reg [fgallag_WDTH -1:0] I24b498fb5b12c3d4a5c7c9e36be4baf7, I944adac3cc097911cde333e806fa004c;
reg [fgallag_WDTH -1:0] Id33f743a90e9f61fd4267c72442a98fa, I3292848fc7b015c9900b92b702ba7be9;
reg [fgallag_WDTH -1:0] I6423dda227b49522f0d8d79fbfe32ecb, Ie09561c5bcd6107bd956faddcdddc89c;
reg [fgallag_WDTH -1:0] I6d8b1a2ff9d9d4a659ddd018a5ce1ebb, I7e8791674daae63eda82adbe6b3e9819;
reg [fgallag_WDTH -1:0] I591484046d2f6f71badbd09db2dd16bc, I4274fedf54de3b2a34285844c7a34519;
reg [fgallag_WDTH -1:0] Ibd503cf61b9c2e244852302f6ecbfb49, I4fae388e04252b896bd4e9c527a8c0af;
reg [fgallag_WDTH -1:0] I42c86c7d63e8f622277ad4cd492dd142, Ia3c4f467d029cc1ea1c0993e0d314978;
reg [fgallag_WDTH -1:0] I480e64694b2be630cf58cb8d35e978eb, Iba2915482c44bda3566df7c23e109ec8;
reg [fgallag_WDTH -1:0] I0b029a353bcf76708510cbd17e96da2a, I38fe32f3f6de6ff9c3fcb5644ac3eb66;
reg [fgallag_WDTH -1:0] I8d0c242b4c0b43f6d1f3796ae1a1be58, Ie4c4245a318c6b4c8f55c678837c5d02;
reg [fgallag_WDTH -1:0] I71e27087daf4bc19fb7e5851935a31e9, If54d6a9d910097237f3e20059257bf57;
reg [fgallag_WDTH -1:0] Ieff0a4b462cd624e967db20434f0452d, I7f2473ad5dc2bcdf35ccdce4bc5fafef;
reg [fgallag_WDTH -1:0] I835c19cffb04dfb43ef7c362c7a9cea0, I16027735edf5e40e34bd73920ae40fb7;
reg [fgallag_WDTH -1:0] Ic506210a4fc9ec0b663ed4a364951fbf, Ie1f37173af26d46bb2948c7675bb491a;
reg [fgallag_WDTH -1:0] I409f55664c78aaefc044bebb7177392a, Ib819132b8eb007862e294bb775a7cd3b;
reg [fgallag_WDTH -1:0] I9477257b731d59c02213efd459153ea3, Icfd0596c8f143d0536c06d827bc30018;
reg I4da12bc20380296febc560ba65f58a8e ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I2e449260cbba5283dbe9d183eaa3006b <= 'h0;
 Ie43af039b1e5b11fe91210b644a1a31e <= 'h0;
 Iebddca10e7f7c3688d5011f147ffcd4a <= 'h0;
 I93b9a635a3e05192ad53b6e264275aa9 <= 'h0;
 Ie3012c652b244e53fc44455982b5eefa <= 'h0;
 Ie287c2f7d9779d50be27d3d5a9de6a33 <= 'h0;
 Ia9327a6a37a1de7dbf3839eafb5d941e <= 'h0;
 I47705f99ef5cb6172811f4046484597c <= 'h0;
 Ie1c96dc77190cd04130a400e869a5abd <= 'h0;
 Iafcc3b17af5dbd70300172c2e2742206 <= 'h0;
 I47731679e4d0f87f9d19934c25f2bdcb <= 'h0;
 I9608c445e266884a86508e3ea3a53853 <= 'h0;
 I0fb3749641e7b5675524cd796ef4127c <= 'h0;
 Id5b6b690dc055c374a44fb1ecfd54198 <= 'h0;
 I6ae44809304b38046cc0afb4317a3f43 <= 'h0;
 I3ef49ef515a84b68f7bff1fbc0f05be7 <= 'h0;
 I62939bc5509a6ca4278bedb7be3f4534 <= 'h0;
 Ieaaab9e41c6a940e06ce877c3e6faebc <= 'h0;
 Iadf3bdeaff4bc193443ef22aef0ad7b7 <= 'h0;
 Ic65a2079483506c24674715cc402a81b <= 'h0;
 Ia7641d441a79bfea63ba407052928bc5 <= 'h0;
 I299c542d09419d0998b59bf1f184a78a <= 'h0;
 I8aa5ad4f2f437be64a88554e6dfc3c6b <= 'h0;
 Iaf0980a21e4ee5e842a5b6db664264f6 <= 'h0;
 I80df82d24c9507274353efb085b46fda <= 'h0;
 I1db5a382bb7c2317716c3137fd10d07c <= 'h0;
 Icb748243d2a5f8cc86c44566e1732232 <= 'h0;
 I90a0c6bd80d2357d7b865f61a18ae13b <= 'h0;
 I16af13e02ee36dbcdeab785596175a3c <= 'h0;
 Id0e47470fba20bc467a05d0dd09bf560 <= 'h0;
 I944adac3cc097911cde333e806fa004c <= 'h0;
 I3292848fc7b015c9900b92b702ba7be9 <= 'h0;
 Ie09561c5bcd6107bd956faddcdddc89c <= 'h0;
 I7e8791674daae63eda82adbe6b3e9819 <= 'h0;
 I4274fedf54de3b2a34285844c7a34519 <= 'h0;
 I4fae388e04252b896bd4e9c527a8c0af <= 'h0;
 Ia3c4f467d029cc1ea1c0993e0d314978 <= 'h0;
 Iba2915482c44bda3566df7c23e109ec8 <= 'h0;
 I38fe32f3f6de6ff9c3fcb5644ac3eb66 <= 'h0;
 Ie4c4245a318c6b4c8f55c678837c5d02 <= 'h0;
 If54d6a9d910097237f3e20059257bf57 <= 'h0;
 I7f2473ad5dc2bcdf35ccdce4bc5fafef <= 'h0;
 I16027735edf5e40e34bd73920ae40fb7 <= 'h0;
 Ie1f37173af26d46bb2948c7675bb491a <= 'h0;
 Ib819132b8eb007862e294bb775a7cd3b <= 'h0;
 Icfd0596c8f143d0536c06d827bc30018 <= 'h0;
 I4da12bc20380296febc560ba65f58a8e <= 'h0;
end
else
begin
 I2e449260cbba5283dbe9d183eaa3006b <=  Ib215a1b985e00121a1c48cf2ddae939a;
 Ie43af039b1e5b11fe91210b644a1a31e <=  I0d9537bea5895773b487fb385690c92c;
 Iebddca10e7f7c3688d5011f147ffcd4a <=  I287708a4c364df837b06049357518409;
 I93b9a635a3e05192ad53b6e264275aa9 <=  I9e69bf6d258b709d9706052822d9ae16;
 Ie3012c652b244e53fc44455982b5eefa <=  I0d187ebb6dbedda971b33ceebb6f17eb;
 Ie287c2f7d9779d50be27d3d5a9de6a33 <=  I83ab1426707044dca3ed926493081311;
 Ia9327a6a37a1de7dbf3839eafb5d941e <=  Ib402ea81f3ba6d26feac26905f0c5edc;
 I47705f99ef5cb6172811f4046484597c <=  I457501e8372fe81287f139beeaad0452;
 Ie1c96dc77190cd04130a400e869a5abd <=  I6f3ecf6c401215c1242c6d31cb4158d7;
 Iafcc3b17af5dbd70300172c2e2742206 <=  Ia439d59ddaa34c9a8dec425ac4f7aca1;
 I47731679e4d0f87f9d19934c25f2bdcb <=  I11a9a93502a123a616205de5969bd5c8;
 I9608c445e266884a86508e3ea3a53853 <=  I346c6ffdb07c9d7a5939fcd142871ef8;
 I0fb3749641e7b5675524cd796ef4127c <=  I20fa0bb8e0dc75902328a349f0dca139;
 Id5b6b690dc055c374a44fb1ecfd54198 <=  Idb4bf6de8f078619ea6dcb51d8f7d329;
 I6ae44809304b38046cc0afb4317a3f43 <=  I8d2f1e18f0064f50176caa84061bf7ec;
 I3ef49ef515a84b68f7bff1fbc0f05be7 <=  Ic48ab17819fe5de2326e4fcb0a1e84c2;
 I62939bc5509a6ca4278bedb7be3f4534 <=  If7332a4a9a6924d2fcbd0af70ecc0d1b;
 Ieaaab9e41c6a940e06ce877c3e6faebc <=  I65a8d4181ad1817636600b816f41158b;
 Iadf3bdeaff4bc193443ef22aef0ad7b7 <=  I746285d851cff1339ce0b99930415c2b;
 Ic65a2079483506c24674715cc402a81b <=  I3305daafd6c3dc6ceb95673b361f0480;
 Ia7641d441a79bfea63ba407052928bc5 <=  I68babd78d3c2b1d6a064b25a3abd690e;
 I299c542d09419d0998b59bf1f184a78a <=  I9e7d989a414d752920fd69ac7c23ca38;
 I8aa5ad4f2f437be64a88554e6dfc3c6b <=  Ibf1b1639efba4277e759d747abe85e6b;
 Iaf0980a21e4ee5e842a5b6db664264f6 <=  If67570ab71fa30823c9fe1277f35c1fe;
 I80df82d24c9507274353efb085b46fda <=  Ia660cf2aa760392654bbc61cb60d9920;
 I1db5a382bb7c2317716c3137fd10d07c <=  I2bf7c2dabc30d2207f04e0f6970f2287;
 Icb748243d2a5f8cc86c44566e1732232 <=  I75c6cf6f3378e1377047d467a7e827f7;
 I90a0c6bd80d2357d7b865f61a18ae13b <=  Ic3dacf077252960c863e8ec1a880f313;
 I16af13e02ee36dbcdeab785596175a3c <=  I781a85002cfeb3038120fe37047710bc;
 Id0e47470fba20bc467a05d0dd09bf560 <=  I0e8936dc5acf0e7c165d76a8b58f2765;
 I944adac3cc097911cde333e806fa004c <=  I24b498fb5b12c3d4a5c7c9e36be4baf7;
 I3292848fc7b015c9900b92b702ba7be9 <=  Id33f743a90e9f61fd4267c72442a98fa;
 Ie09561c5bcd6107bd956faddcdddc89c <=  I6423dda227b49522f0d8d79fbfe32ecb;
 I7e8791674daae63eda82adbe6b3e9819 <=  I6d8b1a2ff9d9d4a659ddd018a5ce1ebb;
 I4274fedf54de3b2a34285844c7a34519 <=  I591484046d2f6f71badbd09db2dd16bc;
 I4fae388e04252b896bd4e9c527a8c0af <=  Ibd503cf61b9c2e244852302f6ecbfb49;
 Ia3c4f467d029cc1ea1c0993e0d314978 <=  I42c86c7d63e8f622277ad4cd492dd142;
 Iba2915482c44bda3566df7c23e109ec8 <=  I480e64694b2be630cf58cb8d35e978eb;
 I38fe32f3f6de6ff9c3fcb5644ac3eb66 <=  I0b029a353bcf76708510cbd17e96da2a;
 Ie4c4245a318c6b4c8f55c678837c5d02 <=  I8d0c242b4c0b43f6d1f3796ae1a1be58;
 If54d6a9d910097237f3e20059257bf57 <=  I71e27087daf4bc19fb7e5851935a31e9;
 I7f2473ad5dc2bcdf35ccdce4bc5fafef <=  Ieff0a4b462cd624e967db20434f0452d;
 I16027735edf5e40e34bd73920ae40fb7 <=  I835c19cffb04dfb43ef7c362c7a9cea0;
 Ie1f37173af26d46bb2948c7675bb491a <=  Ic506210a4fc9ec0b663ed4a364951fbf;
 Ib819132b8eb007862e294bb775a7cd3b <=  I409f55664c78aaefc044bebb7177392a;
 Icfd0596c8f143d0536c06d827bc30018 <=  I9477257b731d59c02213efd459153ea3;
 I4da12bc20380296febc560ba65f58a8e <=  If379a89ad17fd061bf987e29aa713945;
end
