 reg  ['h3ffff:0] [$clog2('h7000+1)-1:0] I390047da02f7900e98c63675c9b8e3ed ;
