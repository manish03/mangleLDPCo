//`include "GF2_LDPC_fgallag_0x00012_assign_inc.sv"
//always_comb begin
              Ib10d67e2c07b1438e202f7b58974fa8e94cfa1651476e39e36cd90f61705d1c2['h00000] = 
          (!fgallag_sel['h00012]) ? 
                       Id639acb3a3eafcec248bdf33943866f07fefacf8e1d90896c6a07bb83a1177a8['h00000] : //%
                       Id639acb3a3eafcec248bdf33943866f07fefacf8e1d90896c6a07bb83a1177a8['h00001] ;
//end
