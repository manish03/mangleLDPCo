//`include "GF2_LDPC_flogtanh_0x00012_assign_inc.sv"
//always_comb begin
              I5edb7954620e8b8032a9ad41b528b90c9fbed81d94a9becd64145bb694902376['h00000] = 
          (!flogtanh_sel['h00012]) ? 
                       I1e92c8d19105281ae50f051d46adab55b63f3805ee886a8045e61a0f72842ab4['h00000] : //%
                       I1e92c8d19105281ae50f051d46adab55b63f3805ee886a8045e61a0f72842ab4['h00001] ;
//end
