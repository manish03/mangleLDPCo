 reg  ['h1f:0] [$clog2('h7000+1)-1:0] Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d ;
