//`include "GF2_LDPC_flogtanh_0x00011_assign_inc.sv"
//always_comb begin
              I1e92c8d19105281ae50f051d46adab55b63f3805ee886a8045e61a0f72842ab4['h00000] = 
          (!flogtanh_sel['h00011]) ? 
                       I3bcb7ea9f76eac891526e809fd382eaceb4a8f0a204c5ca7f391e7ffd9b7808f['h00000] : //%
                       I3bcb7ea9f76eac891526e809fd382eaceb4a8f0a204c5ca7f391e7ffd9b7808f['h00001] ;
//end
//always_comb begin // 
               I1e92c8d19105281ae50f051d46adab55b63f3805ee886a8045e61a0f72842ab4['h00001] =  I3bcb7ea9f76eac891526e809fd382eaceb4a8f0a204c5ca7f391e7ffd9b7808f['h00002] ;
//end
