              I9752ae2367e1a6c6f7352ea46ab95440 = 
          (!flogtanh_sel[0]) ? 
                       I371284eed470112cb89e1d361a9d40f7: 
                       If0fb2e90431d89d99912918f83036f4c;
              I798dac490a694c8373633de0ebc4a72f = 
          (!flogtanh_sel[0]) ? 
                       I0ee915f21334d38c75f0207e3b052a69: 
                       Icf5a9bd712d310ac17eb2354f884a237;
              I071022266cc4a3e5b31bfa3e084079d7 = 
          (!flogtanh_sel[0]) ? 
                       I3222cf2f98878be3f453560ddb3dc43c: 
                       I2dd9e89f2842e748c1574ad0e7f4dba9;
              Ie1307d4ee93e9125654b49ccf5ead6b1 = 
          (!flogtanh_sel[0]) ? 
                       I667adc16c92bec8f413a1a9bbfc41ce5: 
                       Ie6aa50a44574542826b78fed7d77b76f;
              I880d7d200dbb730929b87b4936abb6b7 = 
          (!flogtanh_sel[0]) ? 
                       Ie97072fa52f483bbd89f019c21152cdf: 
                       I47f153e1cecaa77f1e6e6f07c0220557;
              Ib692b0f0a9bd1601ef72ea3f12452a6a = 
          (!flogtanh_sel[0]) ? 
                       I1b9dcfaf144b48a64b990e5b020d4a02: 
                       Ie32d4bd927d02e547850331db8028177;
              I697f7ccafe006697dd1aa6298a1cd9b7 = 
          (!flogtanh_sel[0]) ? 
                       I0988db7ca497541e372131a0b0e8075e: 
                       Id13b5577b8baa586fedd34d4aab9d9c5;
              I81006820f7f068a2ea7f42564c53345a = 
          (!flogtanh_sel[0]) ? 
                       Iedd0e0f6ee682a131d4f14c4762ea0eb: 
                       I875d7c55914414298f0fbec0b345c92e;
              Ic2dcdead9d2a2f6575fdec1ba1a2833c = 
          (!flogtanh_sel[0]) ? 
                       Ide64c9647c7898867e0d036e9ff95f6e: 
                       Ied6ccabb348ed7e20567011e027c86ad;
              I88648891ecdf43525247de0259c99cb6 = 
          (!flogtanh_sel[0]) ? 
                       Id030b072054c623c7aac5c571d052951: 
                       Ice55fb2e506accf518b4aa18298d017e;
              Ic4cfab074168cc1d247169480fdd03f6 = 
          (!flogtanh_sel[0]) ? 
                       I07a0167dcdfc76612e1b0da251337a7b: 
                       I045e08f48738d395af2b79f25af73732;
              I49b23654497581d82ca47a35e429a6ed = 
          (!flogtanh_sel[0]) ? 
                       I7df57f27a880fe45f78c108f8faba963: 
                       I60204c1d3a96524bbbdf715f95f08fe4;
              I8f05a4f32582e13de9003ea0651b5e9f = 
          (!flogtanh_sel[0]) ? 
                       Id5b9ae91dc900060caffff2520236f66: 
                       I861fe9da6d004ce3998ab54a8c0d62af;
              I317fe175f4bc5b04ed6b72d871974ef9 = 
          (!flogtanh_sel[0]) ? 
                       I95caae0432aeadc0cbe279f9d6f9062b: 
                       Ic9c3b015d5830bf4834a435eba89caa5;
              If84908bb6f231e3fad7d0f4cbab882de = 
          (!flogtanh_sel[0]) ? 
                       I6e18dd1a579e09b80ac113fe85b483b4: 
                       I51c1c8e8df14396c5c77b5013531a84f;
              I4f761cecb0e8b5c1bdab0e913cf3a798 = 
          (!flogtanh_sel[0]) ? 
                       Ie8f75e8e020d43f6a357b5175047c254: 
                       Ie762d8aa151448cbaa0d005a3c01572a;
              Iaf08740a169f6f62bddfde35939f0e54 = 
          (!flogtanh_sel[0]) ? 
                       I293b32c043e20d6baab178319dd1e2f6: 
                       I200aae813b664e02075eeefbc3b4450d;
              I6577387fa85776dd6899c8b6fe15d202 = 
          (!flogtanh_sel[0]) ? 
                       I006264bde45d8df078ef711c221ff387: 
                       I9200a0071528b14dc52e92082768ca97;
              Ib6958647f2dd08482fe95961b7f8dd09 = 
          (!flogtanh_sel[0]) ? 
                       I55761decd7043b4dc82737b9d6ef6e7d: 
                       I4f51d114002bdfd69a31f95c2fa5234c;
              I9ae8ddd960f78a4b6fcf14c9247a8ae5 = 
          (!flogtanh_sel[0]) ? 
                       I796cb71b28957405c10015a2ab7124c6: 
                       Ic85bacce5db48b4dd3f626749f6effa8;
              I7cef29b33735fd849743c3f06a82cba9 = 
          (!flogtanh_sel[0]) ? 
                       I2a508066cf0e07bbe8a91f276fbb3078: 
                       I85913ae95fcd63de45030d583846b1d6;
              I0cc3d5d926f4c45056afe4e02d652768 = 
          (!flogtanh_sel[0]) ? 
                       I971cff06a60916ea3e136b397d4c620b: 
                       I2c363f7abf62c9026d0b0dfe5a51207a;
              I1660f9dcac2e19e275df76b02173f49e = 
          (!flogtanh_sel[0]) ? 
                       Ia5043b0c8ee086c66e683eb115a75484: 
                       I6b7b63ea23c5b4f3c597f121284cd2da;
              I5c3b87e1908cc3d152b01573f7a87f2e = 
          (!flogtanh_sel[0]) ? 
                       I3cf82abadcee2faa1849d0a9a45b051e: 
                       I8b42f5455dd8f6323d7a4e28c0eaa1a9;
              I302648ef72470338675f108cfc2936b0 = 
          (!flogtanh_sel[0]) ? 
                       I608597017b046d92b77226999df90600: 
                       Ia39b908f8d6b63777376ca560cd0cc8d;
              I6e11ba6fced3ffc0d8f8003bf04bdfbf = 
          (!flogtanh_sel[0]) ? 
                       I87ad38ab473927df7c0bd69c6b4b4c5e: 
                       I8e70752f74ecdbe95a7b33ca264d4589;
              Ia73537a3f8f0321742cdd459d952f4af = 
          (!flogtanh_sel[0]) ? 
                       I6e768e27a3f1804919e3f83c050e19ba: 
                       I2285f424ef2b8b2041267c1652155ad0;
              I297ad7a97cf35acb5bfd1d0612044c49 = 
          (!flogtanh_sel[0]) ? 
                       Ibc5b97632aab1e763ac51f8d18edc792: 
                       Ic4a0165bd71d9e586fdc66c824e45224;
              I712af4b1f576a39d2d96aff81da4863a = 
          (!flogtanh_sel[0]) ? 
                       I40de7aeac837276e7b3f0c4b29ce5eca: 
                       I024a746142e5ff074724f92af62f3bd3;
              I4a7d547601279634b9aaa30a51fbf741 = 
          (!flogtanh_sel[0]) ? 
                       I1e54f934fa92e681472d03199991f0b2: 
                       I8cabd17b81e99a86fc8704aaaae629a3;
              Icec463cb0767bf054a74408bc41536b8 = 
          (!flogtanh_sel[0]) ? 
                       I54c1bf986182c83540d950762048a5e3: 
                       Ia5fbeb5be349b8088a749e25a9e6e416;
              I1ac433e960367e2ca78597357deb20a5 = 
          (!flogtanh_sel[0]) ? 
                       I987b220a4729d14e9fc97b57867436e4: 
                       I7f1d9309d3053256134130574b970425;
               I7ca1e2fa8fc3e66fb6e747f2e0808e00 =  I9fd9d5a2a3a34b532bad740b16ce66fb ;
              Id8930a77f5475a80411dfae4698cdfd8 = 
          (!flogtanh_sel[0]) ? 
                       Ia08c041d1aacfbbd1f8d7980923b9b05: 
                       I6805a2f26b1e51f7ac0087e6829b3c5c;
              Ifc5cdac396efc12756b713195f9fd57a = 
          (!flogtanh_sel[0]) ? 
                       Icc11f9d183454b33624bd411710342a0: 
                       I18f145bedd3864fcebd983f9533a5877;
              I504e5446ead186c601225c6664e047c8 = 
          (!flogtanh_sel[0]) ? 
                       Ifa25d4c9ccc3efd1af4e711d3c32e9c5: 
                       I5bbf8f01c5ddaa02516dde3867ec3d78;
              I8d9b55049a74bde1fdf26004008679a6 = 
          (!flogtanh_sel[0]) ? 
                       I3f8fe2d052a6df20dfaac6f88d4fff8a: 
                       I9fbf9bcb6022bb550bc2dbd52f20d05f;
              I155a7cee8b9f8b4d03f59ecde58fde8a = 
          (!flogtanh_sel[0]) ? 
                       Iacd71ce5854c85450463a0a45ebc6a2d: 
                       Id7c1a8f42cc90b7846105cd103b07228;
               I9cd50d02d3f7a189b5e70907ec8d1e73 =  Ic6d94b59cd6f4c7765463694c9fbae3c ;
              I04a06a7a7af3891b0d53b95f24954344 = 
          (!flogtanh_sel[0]) ? 
                       I760f9ff7bc594c98e71080485cc1a082: 
                       Idb9be12ba6807752b0c36f4cc18843cb;
              I21ea05b8f1be5a38bf4a4251644c370c = 
          (!flogtanh_sel[0]) ? 
                       I192119ad6ad1396dd6fd1fab6e4c4cca: 
                       Ib4c62a865f79eaa2aa5fbd12860f2e80;
              I89b558f53cd3391108aaee100bb68698 = 
          (!flogtanh_sel[0]) ? 
                       I5fb195f29a4e02620d2cca6e7f2a8fa0: 
                       I41b4d1d3d5ae22c8fe4f1e0fe20ccac7;
               I0b5cdc03696628bcb061aa2113444e50 =  Ib2afa3be272607c236cbd5410a88e8c2 ;
               I4293b2867a22e5f63df2ee4c19c88f79 =  Ic27ed0f98cad254a72ade8253ccc01d2 ;
               I966aa14cea82d7fd5872c135f0bbab70 =  I6f83f4d8681a17b7e700a38a78917822 ;
               Id87f3e498747081eddc52a1fb671838d =  I8297012f23a474aa863c56e6ab9f77f4 ;
              Iabb62eea1f75ca64312cbb047714b9ca = 
          (!flogtanh_sel[0]) ? 
                       I4d60a4630a93dbf6460fc525f16fb69b: 
                       If6a1f518420fbc246e2524469689a5e7;
               Ie231dafa87260c19f1ac9c33085b94f4 =  I48c55cdc6c1e3bb5e36a5451cb43c5a9 ;
               Ief8246918e80c45898a4c38d0d5c3cbb =  I0d302535ee6928ed74d7b456efaf01e6 ;
               I574b308a0fd88d3f211b2acd576a3efb =  I7a43154a62ef625844cda08b1dfc9c79 ;
               I8b32db6febf453df9d355666241b9a80 =  I51393ac63dc5f8c0898ffa6dd59ee183 ;
               I7066424a4d00d757a4a0af28b0d95166 =  Ibf76adf5511e851727200f4fd60bf34b ;
              Ifc4d0343efb2e2f499cc6d8e37591f48 = 
          (!flogtanh_sel[0]) ? 
                       I2b42badcbe3d18d033edbd6d4663fac6: 
                       I72450aa2c2f2f501a5465f008e95ba4f;
              I1600115eb31dadcd5e87696ca1a34fbd = 
          (!flogtanh_sel[0]) ? 
                       Ib802f2c9c1265a47e5acfc419034488d: 
                       Idb28449172f54add7ac6fd1287543a5b;
               I5dce546007aab5da05bbd33b54ee3dba =  I6b33174bb2786da0ba9ba988a96aa5bf ;
               I6a5b90479676374b60fa668a358b852c =  Ia0e39ef7db11ff2f95f50e6a912e945e ;
               Ieb0c46dc3852312024e2bf158d159f20 =  I994e4d13d16c12025cb60205b8f7559f ;
              I56080da8b243334ef8414a095477c286 = 
          (!flogtanh_sel[0]) ? 
                       Id1e6e9ac8ddad3aedd347aee9f615d9f: 
                       I5a6da3732e0f265ad95269f5a629c1e8;
               I661a66590947450472c1cc6b8dc9239b =  If8773fa380ec5c1199794d4128d443f1 ;
               Ie56fe9b766c784f90771d1335e397e99 =  Iedcc3a589dba858f1193b1be582db24b ;
              Icaa6152af5f6bed3d595d51767c9ec49 = 
          (!flogtanh_sel[0]) ? 
                       I267e058f7db05744d80df6b52be83475: 
                       I5e121581d8a5f81fc84da2fa982d8fd6;
               I99bddf2f101ab41147b2849d22bd8e0c =  I51f875fbf103d8b8093d73279f127843 ;
              I5ef97e1962a901d1e6557c0dfcae036e = 
          (!flogtanh_sel[0]) ? 
                       Ie0e816b57f511fc0479210deebbd9fc1: 
                       Ia7673dc1d477d486371935040ff7dce9;
               I3e1118befba3c769deb7bbf9d1875d00 =  I7df5c4ad52bf35d254a4a14771a28fe7 ;
               I435152993799746e1f967343ce1b106f =  Icb740a93e2adc0a9f18ac25d0c5d018c ;
               I9e10d71db16be96b3087a3a584a5b55b =  Iab732884bb2d4b1781e31c7a1c109000 ;
               Ic943175727986874531ace57f5697df3 =  I3bb2f03bf7d2f7480187062b45c6fdd9 ;
               I18d1d32d1e58254b964c670e0d83c119 =  I1732bcc59b7bad3d08b232d099fdefdc ;
               I96b27127bbc15301b57d83982260853b =  I886251a3307e5fe20788c8e947f4ef37 ;
               I12d97a28ef39f26eb4996aa2f1d9eafb =  I9f2ba5b0600c5eb81cef40d0822d0aea ;
               Iddafd4529ad594eda9835e76efa116bb =  I2e8c68a51f1f1f4e413897791a6823a0 ;
               Ice9aeaff41b923556b30553d8b42da47 =  Id32b88b33bfbcf79ff0a10d447f69619 ;
              I33e7dfa55b2d2ac83a8f57797fcd68db = 
          (!flogtanh_sel[0]) ? 
                       I53c239961c5745db892194a0a62b5d57: 
                       I0ffed4dfc4e97bb477647e5eab3a18f3;
               I5c3dedd601ffa33d7b649b2c08df54e6 =  I46fcaa5311cc831199bb4a5a3dba797e ;
               I1660ea57c727ecd6e71a4e9c4c288b45 =  Id0ca109680ce0cb6603139baeebac59f ;
               I1c9e513f7524f52e24e7e80807a18ac6 =  I873254d95f4a9976acf9210228365521 ;
               I3d1372ff9b830f5eeb50c4e47d322cf7 =  I50e26d2184d04613f297357308e7c91e ;
              I69460735237cd5bd0f26254f6f32e357 = 
          (!flogtanh_sel[0]) ? 
                       Ibf3a99967d7cbab53676fed78da28eb8: 
                       Ifb6cf60f578b5a5dd0c27da72408cbce;
               Iac63249f3101e957234cb4efee5f6771 =  I000bdba9ccdb068a02fd37d2991675b6 ;
               I769cf83f4404ee0d85e6c13b7d0c737b =  Ic36cb86884806afb677ac8fb42aead36 ;
              Ieff66b38feb970b4ab3006fb31e5cce3 = 
          (!flogtanh_sel[0]) ? 
                       I96373fc8bdf40551ef8206b4ba38cd98: 
                       I7b8a50810f6a4c27a23c82330707c4b6;
               Ifbef84b3392347c7e0e52e232d26f9bd =  Id84a4cc9f82244c2357edc537824eb30 ;
               I13989f78ab3eab13b7f0619fb0386e3d =  I33d92c1bdacf71fa60865f1741288cdf ;
              I61af8fbc53b6f763a8b77012fb56be23 = 
          (!flogtanh_sel[0]) ? 
                       I51bc583f480542f3f95241643bb39eee: 
                       I35539407bedb7d43642e952787216ce6;
               Id0969f699976b1041d15d62912a04b5f =  Ifa78beaa6ae7a7a32f4886a14e4d1532 ;
               I3be47f6dae15615b1b6b0cb52bb8cd5a =  Ie87c6bd3452b53ef57df5f420f351434 ;
               Iabe728226ae671218667d92139083a4c =  I8b947b6c3139066fbd5873d5b818183e ;
               I49d60f1269fcc5a98196ac391823ca1a =  I4c3bda40c1fe5dbacee1829e0d60bcab ;
               Ic88cdb92bf89df187d801b480c7c2770 =  Iae9c6245aa98b5758df6d57f8c33ab31 ;
               I60a972d5f2465dd5f9c3665eee4cffc2 =  I413a7fe2255064627ed283d35d910de4 ;
               Iaafcf98c2c079884e32f2bd70972e5b3 =  I61ce1d41fa5221c01f7e9571965eb3fe ;
               I3c4a90a70e7cfe814427262cae88e2a6 =  Ic854870518bb942314f6269c6833ff5a ;
               I7eb2363c8fe8f49f839b59df19165aab =  I4576ad4e2708a5635d93b304f1f10677 ;
               I60bf9f27a86ec731795d79b656e2229c =  I04e75fe6916169cea741152b9fc6600b ;
               I8d4fa08cc0155e81bb2ce4ab9a39df4a =  I11555ad63e8caa81cb02dd9264668a3d ;
              Ie21b4ae619493ef57536508645aa29bb = 
          (!flogtanh_sel[0]) ? 
                       I21a1b05b4e659507fc3ff2077e7d2e8d: 
                       I5af0b1d227ed007db9cd98d8a93b89a6;
               I854fac49e7921a59773ab612181b9569 =  If9bdb9270926fe47e645cea702bf7775 ;
               I20a9b10f04d9eeca6058889d5c930294 =  I500e2c4d34270abc5a6f51cec578a7b5 ;
               I122fde74534a82953b1a5a476e2e8151 =  Id7d81b33ad4bd7ae9df6a69b8e1e3351 ;
               Ia535aa71b5100fd37cb15ba1612d2d52 =  I614d496a5262a7f6ebd9a2d078ad30ac ;
               I8b588d7b4605f968fd007ed894b4ee68 =  I0ce07744582a47bf9cfcbdb2776a04c3 ;
               I88d97aa0544a09e2a0df10ec0a57ea54 =  I6c2a048243ceddc9e31b7a37f74eeac1 ;
               I81cb66f14210612d88911543c3517731 =  If32b0bc17ee8e3a95335b09550f05167 ;
               Ibd10299291ec40ff247b816be64f07ec =  Ib8528ee13f669ca3b7d0fddcc4fe697c ;
               I3e4ecb5c8164f70ca4b16eb004cb276c =  I2ff4fa27b4aef5cca03eff8bb129a9eb ;
               Id5e6fca7b1cebfd4f2caf7465fb678fa =  Ib731ae113881b22a9abea15970d8c906 ;
               I58a570689c10954778a3e3ded8d4f9b4 =  I5f2f0073edbf2de118fb329b9d2f6d2c ;
              I0a8dea5e3f82d6954d294cf3c3c858d2 = 
          (!flogtanh_sel[0]) ? 
                       Ib3f304bc897f97659a51764e156f4002: 
                       I02c642372452e4dc5069ceb96098ff71;
               I9aea2a89a8d17d14da2fccad570cfc7d =  Ie6a18db9c01142eb719b8426919a114d ;
               I8b661503122504ce012fe534dad9c394 =  I94c6e4bc6b9ec661a6d76814aafa1e74 ;
               Ib9a8e5b5096d6c5ed5cc315a5899b8d5 =  If22f0f17b0156ee153508c5e4c9742ff ;
               Iebf5cd787ff1d73dfbe4e52cfbaffc14 =  Iaefac912d485b61e57075ddb0212fc55 ;
               I4096de17c18f5e0af8d288bc6887c6cb =  I805cf823cf1cc902fe63131647d582c5 ;
               I949e53f68343283236a519295c606cc2 =  I68941b5c1b03152c7425aa0a1e347385 ;
               Id9fc0dbdd3cd0709ef28238589312443 =  I49597f093b8baac9c769fce82f7ad0d3 ;
              Idf5ff15e65f46f3b569ef0d634cd5819 = 
          (!flogtanh_sel[0]) ? 
                       I87fcfc6fe1957f42e271128cfa0be7e0: 
                       I37b6525d09e5cd2be4f64b64d380cf06;
               I3d70051f81db3db896a8455dda9f0022 =  Ib915a0bb2acae5abe82646277a50f211 ;
               I737715c7b75b324dca40210b708166ac =  Ib8ef3c757de68cd0afc90a6786286248 ;
               I3deb95e95d3308de220901f8fe6d2ee4 =  Id59e1e3a73e7db64fd4808fed9e3e173 ;
               I5e7775e3bc484bed7a57f04b0cd7ccca =  I097da986a541504f1f641404c1749e43 ;
               Ic557aa69aa946711cc39627fe6133f87 =  Ib834d61619c282eb6994727f4b1fe2dd ;
               I004142a2c8e12e72c3ac4a439b281fcc =  Ib815852a6d56c5ea21f7a23acb120f3b ;
               Ia112b4cab1631793a8cc6291027c616c =  Ifdff70e8ea00c64f13abd0d6da5bc11e ;
               I3d3a0cda05e77a00523ea3f4aae38d82 =  I303191eabaa2211774eb1341a7ce1d32 ;
               I723f34fa0b35af4e77fbecc65d2ca88b =  I4fa399fc2e70ae442ef421db22b5ea9c ;
               I460bbb250271f3fa5414de2e68474fbc =  I3c484edf6cf740303824b22ad09ecdf1 ;
               I1e29e4b5d18509694df3a0e7b7cd2a7d =  I015c6af005c8eb5a6ccdf97fd0073bbd ;
               Ie25c961fe6b06030e848c7b9eb751909 =  Ic9143d7200fec6ef38e6cde1fc13d859 ;
               I16c56d8b22dd23fbb09ebf4f36107cc9 =  Ie7d8d3754dc7cc7ac9fc8ebcbd3bf82a ;
               I1e10a4b5844d25334b74e1088e2d3deb =  I2e1e3933f8ec5db47edbec59fd1772b5 ;
               Ic524b9ac09a3499b67313edee303c53f =  I5c9eba93bf9c01e161dd3bd508980acb ;
               Ie332a236ba72fed22c9d7670390dc3d1 =  I0be6fa3f4ae264a84a3b241edd706034 ;
               Ia04ae82f80fd35c0eb30fd17ec9f74a2 =  I501a61dbbe9a6edfbf51d18b14d96f10 ;
               I009b2657f941367412da0645c61a6161 =  I9a432f4a190d752c5e723107243daa1d ;
               If84fc94571af2905f59753301bfb7fec =  I97a78caa8c75ef80934e8d013fee43a4 ;
               I782050339f5fcecb44819e7cb6dac5d6 =  Iaf87541d81d0e3cefb78aecf3ae9c92f ;
               I5ce602af9806ed123e70480c643be643 =  I19a49d3680e5786fad7060cbc4be4a16 ;
               Id2450e8bc8cad7c46f1d47372a344f12 =  I25054529bc0fe35bd08f6294a2d51f5e ;
               Id074a700da35c1548c27b5d1c7e9eea0 =  I12d2ea504991199ca905ca91925f2d26 ;
               I689e819fcdc296cb4b537538012615f6 =  I5f3af0ef6d4722a508201707b6994fed ;
               Ic2824f1963f1158e7ad33e9c81bc7d08 =  I626fef2cd9d071cb8c797471055cf245 ;
               Id0ae33a482904b109068ad943d76d758 =  Iacdb27c060a48b7ade76d256e858b314 ;
              I7b7386e46768f03c912485c3c80065dc = 
          (!flogtanh_sel[0]) ? 
                       I3dfcd0d247d56f8167bcbc6aea6e3504: 
                       I477e8f9e2ac8c5d142856ec6787e28ac;
               Ib0e71935bab4a9ebf00d9b2d170b571a =  I2865e7f35c36e2cd4a4e3435aa8c7c14 ;
               I4613dca4c7c67e9dffb22110f62d93a1 =  I7d5b2a7bca99f2164a7ba2cfe46b20e1 ;
               Ifc0a83912f31329972ce02109fe40df0 =  I6296deff598d27ebc1a06cb1316a3eb4 ;
               I021270a1b11bc14783313a27684e1a08 =  I6a993db6733d3efe90511bbe7f4d5654 ;
               I0f8f6a239a05dba04dd3b845c9e8ac9b =  I0f8f8ce5dfbc020b547758c239f923c4 ;
               I99d616bf2017cd8e4f019fa9356a4c9f =  I361c911024ff757958306a38c4bf4465 ;
               I48c538d54789fc85a7349065dc33b20d =  I56a419f6f3b841e7e5dbbbcc0e6af190 ;
               Idf3ebc5f6ef593255d94f70583e028ba =  I807e19c30c0328199d5ab2d64593d509 ;
               I5ec053664237ddc305a831b20239a5b3 =  I2ba381005b1ffbcf163c40f2dd92d2f9 ;
               I2150bffc35644044c52346accf50c6a6 =  Ib0db88e9d645459a03e908dbbf6b5803 ;
               I9a16fe81b2e09494fb280b564b2d8447 =  Iec7ceaf0d09a3629dbe42f8926383e83 ;
               I3a78158e0bcd94e117696bd698f00e43 =  Iece0c68af7dff6bbe73e9e2d468585c2 ;
               Ia674fb4751c28067672ed365648d4046 =  I3d2bc0bd4abfa1286242b841ef4f04ba ;
               I7c2f789de92dcd3106cd534d547ff653 =  Ib9161bcd780dcb77507b4851bb21193d ;
               I42484fc96375ed4f28054b45a7a573a4 =  Ie3ac6cf6fedf997b6839abbcee584fce ;
               Ife0e6d58f356f10d7f769f225de5a7cc =  I8506a14aacf97d360aa4c10a91ef184f ;
               Id958719d49aab2d0b082a6d24fe4c3ed =  Iaf3e9f18da33e20e42838b4467d9741c ;
               I6f030649ec413f3a8b1b2818f11fdeb9 =  I8ff4739a83ed374704f039515b99162f ;
               I1b4cbdf5cfa3d8c53d2000918dab9d92 =  I9653890e840ec994e81844c9a34b10ba ;
               Id48425985a33f1512c0dd32361ceb85e =  Iad493aff89cf569ffcc57b8f204c11ad ;
               I37d45d42016be2e2bc96ae6fd4287f97 =  I98207474d16dc958a7e695a56a81b614 ;
               I6715c7f4ac584103721a33ead7ed395b =  I2911a1c5c49beebcd2fe684678ab89ca ;
               Ia8e9d2fd6a51de4383c16a35737a1831 =  I10d423113bbfd394aca2695798b2d4ad ;
               I3efa217d3d93a9a2f15bdcd906a2a230 =  I1e24b9c9e023b6f0b00cdeaa071366a2 ;
               I016707bf26cc19976929a8b14f535455 =  I3d0c2d0d76d54c59e1d282a37e0aeae8 ;
               I698072a5328a85b0b22ec7bc94b8372e =  I929ddfd7ec9bf7b7c2dd2378395a403a ;
               I70a428ae2a62212ed93be37b860e8231 =  I88d063cb6f169e9f1ae067641fc0d802 ;
               I5193a317b4c9d2bf1992ca5cf9936681 =  I4b139847ca9cce5281ceb1d63a453d05 ;
               I9cb0c1a404a77903890379f0f658c70a =  I7648b4562836acb77aebba8b19dc62e8 ;
               I861bb6fa26ecdc43776d01811abe7bc3 =  I159acdea94fb6185fccd6310e9d1b071 ;
               I92ad6f4d3a62fbd3e86cda7457115093 =  Ifa65fb0d14e454b62f138630d2f9f370 ;
               I17f6c0345023a3824d5e40506e4c1919 =  Ic888c593409b429e20523b414861da69 ;
               Ic309d272e0e79647de87c07aae1e798c =  I3c6576aed9ae9c1a1e86afdc00082fc0 ;
               I24a4c216e917b9b9ad744c7bfa4a7d24 =  Ic6e2dd06abadb6b0613d8be1d3e91da7 ;
              I7112d906a2a8245dd62b7ef26d7e54ee = 
          (!flogtanh_sel[0]) ? 
                       Ieb48cc2ae37e2d9dd9144b587cce78da: 
                       I0c2ea6ea58ccc53502b8765d9ab08a56;
