 reg  ['h3ff:0] [$clog2('h7000+1)-1:0] I810764ca41a2b12d686e115c79b0578f ;
