 reg  ['h3fff:0] [$clog2('h7000+1)-1:0] Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748 ;
