 reg  ['h3f:0] [$clog2('h7000+1)-1:0] I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef ;
