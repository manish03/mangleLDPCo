              I702f756fc12e54b5d0cba9e129e16e40 = 
          (!fgallag_sel[7]) ? 
                       Iac8fa9870b8eea066f71cf779822ae8c: 
                       I21bf34a5a15ad45c1589e27caefe01b3;
              I8ed18c5f09ca2d107ccf511f4efee704 = 
          (!fgallag_sel[7]) ? 
                       I741862871bd1eede0465be591cb86701: 
                       I89a7e0136bed29f84bb4a16c895927e7;
