`include "flogtanh/GF2_LDPC_flogtanh.sv.1"
`include "flogtanh/GF2_LDPC_flogtanh.sv.2"
