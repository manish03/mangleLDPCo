 reg  ['h1:0] [$clog2('h7000+1)-1:0] Id639acb3a3eafcec248bdf33943866f07fefacf8e1d90896c6a07bb83a1177a8 ;
