 reg  ['hff:0] [$clog2('h7000+1)-1:0] I1a62004aa5608ddf7a551106f9a8a7ac ;
