 reg  ['hfff:0] [$clog2('h7000+1)-1:0] I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9 ;
