//`include "GF2_LDPC_flogtanh_0x00011_assign_inc.sv"
//always_comb begin
              Ic7e91188980d728ad34dbe693d9a6e04['h00000] = 
          (!flogtanh_sel['h00011]) ? 
                       Ib43d6a3ec9a1741fe7beed3535eddb34['h00000] : //%
                       Ib43d6a3ec9a1741fe7beed3535eddb34['h00001] ;
//end
//always_comb begin // 
               Ic7e91188980d728ad34dbe693d9a6e04['h00001] =  Ib43d6a3ec9a1741fe7beed3535eddb34['h00002] ;
//end
