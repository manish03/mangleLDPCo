              Ic95a3f9bce1f573855ca615170882870 = 
          (!fgallag_sel[5]) ? 
                       I45d771e861cb0c71b24703a4630c0cf2: 
                       I5da352fc142fd74387413bbd1fba6775;
              I7b13a2539c028f1b1704554ec14280f5 = 
          (!fgallag_sel[5]) ? 
                       I404ff307c40124efe47cd1aa98a26ed2: 
                       I437d32d746b0a046d3b0620972b129a1;
              I9b426da62c1159dd95754d51e3d8b4e8 = 
          (!fgallag_sel[5]) ? 
                       I4b608f7adccf4eefe0909c711022bc17: 
                       Ief186188e0a216ead6c35d9a77ec4b76;
              I77a77a7a6a437c395358b6f0beafd9f2 = 
          (!fgallag_sel[5]) ? 
                       I09e7fa2c8569782c6c9a3e507c5bec16: 
                       I784d791eaf69fdc5ea6c1033592ab5e8;
              I1efd99d9686a0c7e1187d852a3572023 = 
          (!fgallag_sel[5]) ? 
                       I1a54ecd582987b3bbbdc797c8abc7f30: 
                       I1977cd7fe67cd9d9b7f2aeabbdbe4b0e;
              Ia0c03de62b7bfb76e6fea17bd0e8d003 = 
          (!fgallag_sel[5]) ? 
                       Ia8b47732674c465cea9957ee0eea7f22: 
                       I7cdb7e144a06928d0a616bda0b1fb4c0;
