//`include "GF2_LDPC_flogtanh_0x0000e_assign_inc.sv"
//always_comb begin
              Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00000] = 
          (!flogtanh_sel['h0000e]) ? 
                       Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00000] : //%
                       Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00001] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00001] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00002] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00002] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00004] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00003] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00006] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00004] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00008] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00005] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000a] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00006] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000c] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00007] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000e] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00008] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00010] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h00009] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00012] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000a] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00014] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000b] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00016] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000c] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00018] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000d] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001a] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000e] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001c] ;
//end
//always_comb begin // 
               Ica808b9c1910a49740bb889b7521538bc786bf51f6b2c7c3ad1af9712127147b['h0000f] =  Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001e] ;
//end
