 reg  ['h0:0] [$clog2('h7000+1)-1:0] Ia9be81772a42d1908d7f14f7ec313644 ;
