 reg  ['h7ff:0] [$clog2('h7000+1)-1:0] Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756 ;
