reg [fgallag_WDTH -1:0] Iad95cb311111b88124c0d2a123589b68, I45d771e861cb0c71b24703a4630c0cf2;
reg [fgallag_WDTH -1:0] I8efbaa789c07fd87b2bd52379ef30fd6, I5da352fc142fd74387413bbd1fba6775;
reg [fgallag_WDTH -1:0] I75d6885c5406c2c71dc966efa9c6826d, I404ff307c40124efe47cd1aa98a26ed2;
reg [fgallag_WDTH -1:0] I3f698aa4ba3738ea0af307eff19d7322, I437d32d746b0a046d3b0620972b129a1;
reg [fgallag_WDTH -1:0] I3dcfc9ea0f47bae945b7b823693115ad, I4b608f7adccf4eefe0909c711022bc17;
reg [fgallag_WDTH -1:0] Id1a3fd12101241027e2f457a826ed09d, Ief186188e0a216ead6c35d9a77ec4b76;
reg [fgallag_WDTH -1:0] I7bfcc4e396adf33cfc50d06be12d9007, I09e7fa2c8569782c6c9a3e507c5bec16;
reg [fgallag_WDTH -1:0] I5ce36b9e0a8e3e118e1f1b9eae183b7b, I784d791eaf69fdc5ea6c1033592ab5e8;
reg [fgallag_WDTH -1:0] I98f08554298bf8e87fc54a4f8c668314, I1a54ecd582987b3bbbdc797c8abc7f30;
reg [fgallag_WDTH -1:0] Ic05153bb88b7db4e173fd73841f88bf2, I1977cd7fe67cd9d9b7f2aeabbdbe4b0e;
reg [fgallag_WDTH -1:0] I75df32ec8d8f7096f5f7ef1d17cfb8e7, Ia8b47732674c465cea9957ee0eea7f22;
reg [fgallag_WDTH -1:0] Ia3c542d3f12470683609d561d9cd0e35, I7cdb7e144a06928d0a616bda0b1fb4c0;
reg If677b4bb108ef735b4ad076cbbfd3094 ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I45d771e861cb0c71b24703a4630c0cf2 <= 'h0;
 I5da352fc142fd74387413bbd1fba6775 <= 'h0;
 I404ff307c40124efe47cd1aa98a26ed2 <= 'h0;
 I437d32d746b0a046d3b0620972b129a1 <= 'h0;
 I4b608f7adccf4eefe0909c711022bc17 <= 'h0;
 Ief186188e0a216ead6c35d9a77ec4b76 <= 'h0;
 I09e7fa2c8569782c6c9a3e507c5bec16 <= 'h0;
 I784d791eaf69fdc5ea6c1033592ab5e8 <= 'h0;
 I1a54ecd582987b3bbbdc797c8abc7f30 <= 'h0;
 I1977cd7fe67cd9d9b7f2aeabbdbe4b0e <= 'h0;
 Ia8b47732674c465cea9957ee0eea7f22 <= 'h0;
 I7cdb7e144a06928d0a616bda0b1fb4c0 <= 'h0;
 If677b4bb108ef735b4ad076cbbfd3094 <= 'h0;
end
else
begin
 I45d771e861cb0c71b24703a4630c0cf2 <=  Iad95cb311111b88124c0d2a123589b68;
 I5da352fc142fd74387413bbd1fba6775 <=  I8efbaa789c07fd87b2bd52379ef30fd6;
 I404ff307c40124efe47cd1aa98a26ed2 <=  I75d6885c5406c2c71dc966efa9c6826d;
 I437d32d746b0a046d3b0620972b129a1 <=  I3f698aa4ba3738ea0af307eff19d7322;
 I4b608f7adccf4eefe0909c711022bc17 <=  I3dcfc9ea0f47bae945b7b823693115ad;
 Ief186188e0a216ead6c35d9a77ec4b76 <=  Id1a3fd12101241027e2f457a826ed09d;
 I09e7fa2c8569782c6c9a3e507c5bec16 <=  I7bfcc4e396adf33cfc50d06be12d9007;
 I784d791eaf69fdc5ea6c1033592ab5e8 <=  I5ce36b9e0a8e3e118e1f1b9eae183b7b;
 I1a54ecd582987b3bbbdc797c8abc7f30 <=  I98f08554298bf8e87fc54a4f8c668314;
 I1977cd7fe67cd9d9b7f2aeabbdbe4b0e <=  Ic05153bb88b7db4e173fd73841f88bf2;
 Ia8b47732674c465cea9957ee0eea7f22 <=  I75df32ec8d8f7096f5f7ef1d17cfb8e7;
 I7cdb7e144a06928d0a616bda0b1fb4c0 <=  Ia3c542d3f12470683609d561d9cd0e35;
 If677b4bb108ef735b4ad076cbbfd3094 <=  I64ddd9e95d971d161174a6dd0c3d2fbe;
end
