`include "GF2_LDPC_fgallag_inc.sv"
`include "GF2_LDPC_fgallag_0x00000_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00001_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00002_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00003_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00004_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00005_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00006_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00007_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00008_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00009_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x0000a_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x0000b_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x0000c_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x0000d_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x0000e_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x0000f_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00010_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00011_assign_inc.sv"
`include "GF2_LDPC_fgallag_0x00012_assign_inc.sv"
