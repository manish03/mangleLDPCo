`include "flogtanh/GF2_LDPC_flogtanh_0x00000_assign.sv.1"
`include "flogtanh/GF2_LDPC_flogtanh_0x00000_assign.sv.2"
