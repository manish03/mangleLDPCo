//`include "GF2_LDPC_flogtanh_0x00005_assign_inc.sv"
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00000] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00000] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00001] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00001] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00002] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00003] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00002] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00004] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00005] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00003] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00006] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00007] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00004] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00008] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00009] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00005] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00006] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00007] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0000f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00008] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00010] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00011] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00009] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00012] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00013] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00014] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00015] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00016] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00017] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00018] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00019] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0000f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0001f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00010] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00020] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00021] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00011] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00022] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00023] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00012] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00024] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00025] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00013] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00026] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00027] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00014] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00028] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00029] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00015] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00016] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00017] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0002f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00018] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00030] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00031] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00019] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00032] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00033] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00034] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00035] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00036] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00037] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00038] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00039] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0001f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0003f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00020] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00040] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00041] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00021] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00042] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00043] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00022] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00044] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00045] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00023] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00046] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00047] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00024] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00048] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00049] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00025] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00026] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00027] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0004f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00028] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00050] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00051] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00029] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00052] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00053] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00054] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00055] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00056] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00057] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00058] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00059] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0002f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0005f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00030] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00060] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00061] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00031] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00062] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00063] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00032] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00064] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00065] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00033] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00066] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00067] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00034] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00068] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00069] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00035] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00036] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00037] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0006f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00038] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00070] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00071] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00039] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00072] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00073] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00074] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00075] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00076] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00077] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00078] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00079] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0003f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0007f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00040] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00080] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00081] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00041] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00082] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00083] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00042] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00084] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00085] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00043] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00086] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00087] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00044] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00088] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00089] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00045] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00046] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00047] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0008f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00048] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00090] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00091] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00049] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00092] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00093] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00094] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00095] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00096] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00097] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00098] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00099] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0004f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0009f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00050] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a0] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a1] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00051] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a2] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a3] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00052] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a4] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a5] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00053] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a6] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a7] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00054] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a8] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000a9] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00055] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000aa] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ab] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00056] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ac] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ad] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00057] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ae] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000af] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00058] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b0] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b1] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00059] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b2] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b3] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b4] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b5] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b6] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b7] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b8] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000b9] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ba] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000bb] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000bc] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000bd] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0005f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000be] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000bf] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00060] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c0] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c1] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00061] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c2] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c3] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00062] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c4] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c5] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00063] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c6] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c7] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00064] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c8] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000c9] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00065] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ca] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000cb] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00066] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000cc] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000cd] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00067] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ce] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000cf] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00068] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d0] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d1] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00069] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d2] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d3] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d4] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d5] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d6] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d7] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d8] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000d9] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000da] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000db] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000dc] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000dd] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0006f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000de] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000df] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00070] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e0] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e1] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00071] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e2] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e3] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00072] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e4] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e5] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00073] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e6] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e7] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00074] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e8] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000e9] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00075] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ea] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000eb] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00076] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ec] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ed] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00077] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ee] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ef] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00078] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f0] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f1] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00079] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f2] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f3] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f4] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f5] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f6] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f7] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f8] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000f9] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fa] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fb] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fc] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fd] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0007f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000fe] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h000ff] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00080] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00100] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00101] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00081] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00102] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00103] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00082] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00104] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00105] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00083] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00106] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00107] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00084] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00108] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00109] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00085] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00086] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00087] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0010f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00088] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00110] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00111] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00089] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00112] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00113] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00114] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00115] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00116] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00117] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00118] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00119] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0008f] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0011f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00090] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00120] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00121] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00091] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00122] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00123] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00092] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00124] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00125] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00093] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00126] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00127] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00094] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00128] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00129] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00095] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00096] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012d] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00097] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012e] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0012f] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00098] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00130] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00131] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00099] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00132] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00133] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009a] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00134] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00135] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009b] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00136] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00137] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009c] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00138] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00139] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009d] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009e] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013d] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0009f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0013e] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a0] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00140] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00141] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a1] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00142] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00143] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a2] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00144] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00145] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a3] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00146] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00147] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00148] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a5] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014b] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a6] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014d] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0014e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00150] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000a9] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00152] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00153] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00154] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ab] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00156] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00157] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ac] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00158] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00159] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015a] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ae] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015d] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0015e] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b0] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00160] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00161] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00162] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b2] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00164] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00165] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00166] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b4] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00168] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00169] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016a] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b6] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016d] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0016e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00170] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000b9] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00172] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00173] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00174] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00176] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000bc] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00178] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00179] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017a] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000be] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017d] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0017e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00180] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00182] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c2] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00184] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00185] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00186] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00188] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c5] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018a] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018b] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0018e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00190] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000c9] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00192] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00193] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00194] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00196] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00198] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019a] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ce] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019c] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019d] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0019e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a4] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d3] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a6] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a7] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b2] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000da] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b4] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b5] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c2] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e2] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c4] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c5] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d6] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ec] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d8] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001d9] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001f8] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fd] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fa] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fb] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h000ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h001fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00100] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00200] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00101] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00202] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00102] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00204] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00103] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00206] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00104] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00208] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00105] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00106] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00107] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0020e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00108] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00210] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00109] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00212] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00214] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00216] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00218] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0010f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0021e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00110] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00220] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00111] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00222] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00112] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00224] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00113] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00226] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00114] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00228] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00115] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00116] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00117] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0022e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00118] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00230] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00119] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00232] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00234] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00236] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00238] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0011f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0023e] ;
//end
//always_comb begin
              I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00120] = 
          (!flogtanh_sel['h00005]) ? 
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00240] : //%
                       Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00241] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00121] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00242] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00122] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00244] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00123] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00246] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00124] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00248] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00125] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00126] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00127] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0024e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00128] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00250] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00129] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00252] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00254] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00256] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00258] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0012f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0025e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00130] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00260] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00131] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00262] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00132] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00264] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00133] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00266] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00134] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00268] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00135] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00136] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00137] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0026e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00138] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00270] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00139] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00272] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00274] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00276] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00278] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0013f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0027e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00140] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00280] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00141] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00282] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00142] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00284] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00143] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00286] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00144] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00288] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00145] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00146] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00147] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0028e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00148] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00290] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00149] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00292] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00294] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00296] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00298] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0014f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0029e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00150] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00151] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00152] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00153] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00154] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00155] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00156] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00157] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00158] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00159] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0015f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00160] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00161] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00162] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00163] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00164] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00165] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00166] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00167] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00168] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00169] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0016f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00170] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00171] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00172] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00173] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00174] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00175] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00176] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00177] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00178] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00179] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0017f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h002fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00180] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00300] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00181] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00302] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00182] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00304] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00183] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00306] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00184] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00308] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00185] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00186] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00187] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0030e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00188] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00310] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00189] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00312] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00314] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00316] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00318] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0018f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0031e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00190] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00320] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00191] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00322] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00192] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00324] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00193] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00326] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00194] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00328] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00195] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00196] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00197] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0032e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00198] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00330] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00199] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00332] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00334] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00336] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00338] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0019f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0033e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00340] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00342] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00344] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00346] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00348] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0034e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00350] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00352] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00354] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00356] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00358] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0035e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00360] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00362] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00364] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00366] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00368] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0036e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00370] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00372] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00374] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00376] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00378] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0037e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00380] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00382] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00384] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00386] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00388] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0038e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00390] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00392] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00394] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00396] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00398] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0039e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h001ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h003fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00200] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00400] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00201] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00402] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00202] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00404] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00203] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00406] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00204] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00408] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00205] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00206] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00207] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0040e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00208] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00410] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00209] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00412] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00414] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00416] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00418] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0020f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0041e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00210] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00420] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00211] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00422] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00212] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00424] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00213] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00426] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00214] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00428] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00215] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00216] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00217] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0042e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00218] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00430] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00219] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00432] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00434] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00436] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00438] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0021f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0043e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00220] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00440] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00221] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00442] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00222] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00444] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00223] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00446] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00224] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00448] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00225] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00226] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00227] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0044e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00228] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00450] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00229] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00452] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00454] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00456] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00458] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0022f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0045e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00230] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00460] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00231] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00462] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00232] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00464] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00233] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00466] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00234] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00468] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00235] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00236] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00237] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0046e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00238] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00470] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00239] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00472] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00474] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00476] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00478] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0023f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0047e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00240] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00480] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00241] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00482] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00242] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00484] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00243] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00486] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00244] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00488] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00245] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00246] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00247] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0048e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00248] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00490] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00249] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00492] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00494] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00496] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00498] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0024f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0049e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00250] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00251] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00252] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00253] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00254] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00255] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00256] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00257] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00258] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00259] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0025f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00260] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00261] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00262] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00263] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00264] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00265] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00266] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00267] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00268] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00269] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0026f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00270] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00271] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00272] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00273] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00274] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00275] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00276] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00277] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00278] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00279] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0027f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h004fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00280] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00500] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00281] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00502] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00282] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00504] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00283] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00506] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00284] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00508] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00285] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00286] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00287] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0050e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00288] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00510] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00289] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00512] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00514] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00516] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00518] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0028f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0051e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00290] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00520] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00291] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00522] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00292] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00524] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00293] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00526] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00294] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00528] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00295] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00296] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00297] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0052e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00298] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00530] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00299] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00532] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00534] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00536] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00538] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0029f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0053e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00540] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00542] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00544] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00546] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00548] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0054e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00550] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00552] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00554] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00556] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00558] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0055e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00560] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00562] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00564] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00566] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00568] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0056e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00570] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00572] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00574] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00576] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00578] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0057e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00580] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00582] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00584] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00586] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00588] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0058e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00590] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00592] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00594] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00596] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00598] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0059e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h002ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h005fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00300] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00600] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00301] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00602] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00302] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00604] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00303] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00606] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00304] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00608] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00305] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00306] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00307] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0060e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00308] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00610] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00309] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00612] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00614] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00616] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00618] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0030f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0061e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00310] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00620] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00311] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00622] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00312] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00624] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00313] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00626] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00314] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00628] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00315] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00316] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00317] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0062e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00318] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00630] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00319] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00632] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00634] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00636] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00638] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0031f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0063e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00320] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00640] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00321] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00642] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00322] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00644] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00323] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00646] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00324] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00648] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00325] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00326] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00327] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0064e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00328] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00650] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00329] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00652] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00654] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00656] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00658] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0032f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0065e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00330] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00660] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00331] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00662] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00332] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00664] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00333] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00666] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00334] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00668] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00335] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00336] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00337] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0066e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00338] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00670] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00339] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00672] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00674] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00676] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00678] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0033f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0067e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00340] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00680] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00341] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00682] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00342] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00684] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00343] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00686] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00344] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00688] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00345] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00346] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00347] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0068e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00348] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00690] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00349] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00692] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00694] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00696] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00698] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0034f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0069e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00350] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00351] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00352] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00353] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00354] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00355] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00356] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00357] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00358] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00359] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0035f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00360] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00361] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00362] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00363] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00364] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00365] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00366] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00367] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00368] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00369] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0036f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00370] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00371] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00372] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00373] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00374] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00375] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00376] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00377] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00378] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00379] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0037f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h006fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00380] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00700] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00381] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00702] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00382] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00704] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00383] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00706] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00384] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00708] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00385] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00386] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00387] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0070e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00388] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00710] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00389] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00712] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00714] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00716] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00718] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0038f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0071e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00390] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00720] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00391] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00722] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00392] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00724] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00393] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00726] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00394] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00728] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00395] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00396] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00397] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0072e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00398] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00730] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00399] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00732] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00734] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00736] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00738] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0039f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0073e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00740] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00742] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00744] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00746] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00748] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0074e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00750] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00752] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00754] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00756] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00758] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0075e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00760] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00762] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00764] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00766] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00768] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0076e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00770] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00772] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00774] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00776] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00778] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0077e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00780] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00782] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00784] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00786] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00788] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0078e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00790] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00792] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00794] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00796] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00798] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0079e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h003ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h007fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00400] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00800] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00401] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00802] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00402] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00804] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00403] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00806] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00404] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00808] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00405] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00406] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00407] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0080e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00408] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00810] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00409] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00812] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00814] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00816] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00818] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0040f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0081e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00410] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00820] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00411] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00822] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00412] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00824] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00413] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00826] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00414] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00828] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00415] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00416] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00417] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0082e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00418] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00830] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00419] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00832] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00834] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00836] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00838] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0041f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0083e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00420] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00840] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00421] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00842] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00422] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00844] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00423] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00846] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00424] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00848] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00425] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00426] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00427] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0084e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00428] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00850] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00429] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00852] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00854] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00856] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00858] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0042f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0085e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00430] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00860] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00431] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00862] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00432] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00864] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00433] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00866] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00434] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00868] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00435] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00436] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00437] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0086e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00438] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00870] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00439] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00872] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00874] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00876] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00878] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0043f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0087e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00440] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00880] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00441] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00882] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00442] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00884] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00443] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00886] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00444] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00888] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00445] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00446] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00447] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0088e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00448] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00890] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00449] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00892] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00894] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00896] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00898] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0044f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0089e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00450] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00451] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00452] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00453] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00454] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00455] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00456] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00457] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00458] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00459] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0045f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00460] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00461] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00462] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00463] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00464] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00465] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00466] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00467] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00468] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00469] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0046f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00470] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00471] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00472] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00473] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00474] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00475] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00476] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00477] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00478] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00479] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0047f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h008fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00480] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00900] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00481] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00902] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00482] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00904] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00483] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00906] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00484] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00908] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00485] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00486] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00487] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0090e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00488] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00910] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00489] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00912] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00914] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00916] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00918] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0048f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0091e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00490] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00920] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00491] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00922] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00492] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00924] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00493] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00926] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00494] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00928] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00495] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00496] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00497] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0092e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00498] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00930] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00499] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00932] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00934] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00936] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00938] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0049f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0093e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00940] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00942] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00944] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00946] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00948] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0094e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00950] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00952] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00954] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00956] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00958] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0095e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00960] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00962] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00964] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00966] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00968] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0096e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00970] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00972] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00974] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00976] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00978] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0097e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00980] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00982] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00984] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00986] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00988] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0098e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00990] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00992] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00994] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00996] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00998] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0099e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h004ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h009fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00500] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00501] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00502] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00503] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00504] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00505] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00506] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00507] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00508] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00509] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0050f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00510] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00511] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00512] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00513] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00514] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00515] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00516] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00517] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00518] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00519] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0051f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00520] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00521] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00522] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00523] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00524] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00525] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00526] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00527] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00528] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00529] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0052f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00530] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00531] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00532] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00533] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00534] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00535] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00536] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00537] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00538] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00539] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0053f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00540] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00541] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00542] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00543] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00544] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00545] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00546] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00547] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00548] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00549] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0054f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00a9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00550] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00551] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00552] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00553] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00554] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aa8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00555] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aaa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00556] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00557] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00558] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00559] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ab8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00abc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0055f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00abe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00560] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00561] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00562] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00563] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00564] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ac8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00565] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00566] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00acc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00567] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ace] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00568] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00569] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ad8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ada] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00adc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0056f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ade] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00570] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00571] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00572] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00573] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00574] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ae8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00575] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00576] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00577] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00aee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00578] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00579] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00af8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00afa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00afc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0057f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00afe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00580] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00581] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00582] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00583] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00584] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00585] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00586] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00587] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00588] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00589] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0058f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00590] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00591] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00592] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00593] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00594] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00595] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00596] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00597] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00598] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00599] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0059f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00b9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ba8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00baa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00be8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bf8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h005ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00bfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00600] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00601] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00602] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00603] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00604] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00605] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00606] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00607] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00608] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00609] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0060f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00610] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00611] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00612] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00613] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00614] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00615] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00616] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00617] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00618] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00619] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0061f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00620] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00621] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00622] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00623] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00624] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00625] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00626] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00627] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00628] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00629] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0062f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00630] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00631] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00632] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00633] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00634] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00635] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00636] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00637] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00638] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00639] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0063f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00640] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00641] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00642] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00643] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00644] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00645] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00646] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00647] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00648] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00649] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0064f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00c9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00650] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00651] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00652] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00653] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00654] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ca8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00655] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00caa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00656] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00657] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00658] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00659] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0065f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00660] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00661] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00662] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00663] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00664] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00665] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00666] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ccc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00667] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00668] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00669] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0066f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00670] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00671] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00672] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00673] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00674] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ce8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00675] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00676] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00677] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00678] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00679] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cf8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0067f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00cfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00680] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00681] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00682] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00683] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00684] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00685] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00686] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00687] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00688] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00689] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0068f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00690] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00691] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00692] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00693] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00694] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00695] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00696] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00697] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00698] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00699] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0069f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00d9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00da8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00daa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00db8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ddc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00de8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00df8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h006ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00dfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00700] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00701] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00702] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00703] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00704] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00705] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00706] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00707] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00708] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00709] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0070f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00710] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00711] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00712] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00713] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00714] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00715] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00716] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00717] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00718] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00719] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0071f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00720] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00721] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00722] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00723] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00724] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00725] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00726] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00727] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00728] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00729] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0072f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00730] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00731] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00732] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00733] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00734] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00735] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00736] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00737] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00738] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00739] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0073f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00740] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00741] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00742] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00743] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00744] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00745] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00746] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00747] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00748] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00749] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0074f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00e9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00750] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00751] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00752] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00753] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00754] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ea8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00755] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eaa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00756] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00757] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00758] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00759] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ebc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0075f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ebe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00760] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00761] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00762] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00763] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00764] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ec8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00765] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00766] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ecc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00767] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ece] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00768] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00769] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ed8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00edc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0076f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ede] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00770] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00771] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00772] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00773] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00774] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ee8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00775] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00776] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00777] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00eee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00778] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00779] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ef8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00efa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00efc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0077f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00efe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00780] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00781] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00782] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00783] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00784] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00785] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00786] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00787] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00788] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00789] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0078f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00790] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00791] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00792] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00793] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00794] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00795] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00796] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00797] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00798] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00799] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0079f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00f9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fa8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00faa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fe8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00fee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ff8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ffa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ffc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h007ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h00ffe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00800] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01000] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00801] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01002] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00802] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01004] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00803] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01006] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00804] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01008] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00805] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00806] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00807] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0100e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00808] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01010] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00809] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01012] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01014] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01016] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01018] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0080f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0101e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00810] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01020] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00811] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01022] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00812] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01024] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00813] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01026] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00814] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01028] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00815] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00816] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00817] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0102e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00818] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01030] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00819] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01032] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01034] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01036] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01038] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0081f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0103e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00820] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01040] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00821] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01042] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00822] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01044] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00823] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01046] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00824] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01048] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00825] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00826] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00827] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0104e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00828] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01050] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00829] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01052] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01054] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01056] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01058] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0082f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0105e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00830] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01060] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00831] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01062] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00832] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01064] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00833] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01066] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00834] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01068] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00835] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00836] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00837] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0106e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00838] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01070] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00839] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01072] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01074] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01076] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01078] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0083f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0107e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00840] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01080] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00841] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01082] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00842] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01084] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00843] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01086] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00844] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01088] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00845] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00846] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00847] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0108e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00848] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01090] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00849] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01092] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01094] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01096] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01098] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0084f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0109e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00850] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00851] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00852] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00853] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00854] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00855] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00856] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00857] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00858] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00859] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0085f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00860] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00861] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00862] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00863] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00864] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00865] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00866] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00867] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00868] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00869] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0086f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00870] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00871] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00872] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00873] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00874] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00875] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00876] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00877] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00878] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00879] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0087f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h010fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00880] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01100] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00881] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01102] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00882] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01104] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00883] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01106] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00884] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01108] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00885] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00886] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00887] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0110e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00888] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01110] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00889] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01112] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01114] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01116] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01118] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0088f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0111e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00890] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01120] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00891] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01122] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00892] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01124] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00893] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01126] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00894] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01128] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00895] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00896] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00897] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0112e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00898] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01130] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00899] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01132] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01134] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01136] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01138] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0089f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0113e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01140] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01142] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01144] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01146] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01148] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0114e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01150] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01152] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01154] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01156] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01158] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0115e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01160] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01162] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01164] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01166] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01168] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0116e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01170] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01172] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01174] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01176] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01178] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0117e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01180] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01182] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01184] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01186] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01188] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0118e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01190] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01192] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01194] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01196] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01198] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0119e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h008ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h011fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00900] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01200] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00901] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01202] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00902] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01204] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00903] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01206] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00904] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01208] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00905] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00906] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00907] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0120e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00908] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01210] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00909] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01212] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01214] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01216] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01218] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0090f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0121e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00910] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01220] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00911] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01222] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00912] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01224] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00913] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01226] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00914] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01228] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00915] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00916] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00917] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0122e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00918] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01230] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00919] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01232] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01234] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01236] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01238] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0091f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0123e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00920] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01240] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00921] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01242] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00922] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01244] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00923] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01246] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00924] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01248] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00925] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00926] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00927] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0124e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00928] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01250] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00929] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01252] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01254] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01256] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01258] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0092f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0125e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00930] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01260] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00931] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01262] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00932] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01264] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00933] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01266] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00934] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01268] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00935] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00936] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00937] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0126e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00938] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01270] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00939] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01272] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01274] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01276] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01278] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0093f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0127e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00940] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01280] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00941] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01282] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00942] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01284] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00943] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01286] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00944] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01288] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00945] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00946] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00947] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0128e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00948] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01290] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00949] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01292] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01294] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01296] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01298] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0094f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0129e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00950] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00951] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00952] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00953] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00954] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00955] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00956] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00957] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00958] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00959] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0095f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00960] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00961] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00962] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00963] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00964] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00965] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00966] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00967] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00968] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00969] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0096f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00970] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00971] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00972] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00973] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00974] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00975] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00976] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00977] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00978] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00979] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0097f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h012fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00980] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01300] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00981] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01302] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00982] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01304] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00983] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01306] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00984] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01308] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00985] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00986] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00987] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0130e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00988] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01310] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00989] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01312] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01314] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01316] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01318] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0098f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0131e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00990] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01320] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00991] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01322] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00992] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01324] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00993] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01326] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00994] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01328] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00995] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00996] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00997] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0132e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00998] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01330] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00999] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01332] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01334] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01336] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01338] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0099f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0133e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01340] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01342] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01344] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01346] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01348] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0134e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01350] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01352] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01354] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01356] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01358] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0135e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01360] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01362] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01364] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01366] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01368] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0136e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01370] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01372] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01374] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01376] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01378] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0137e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01380] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01382] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01384] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01386] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01388] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0138e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01390] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01392] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01394] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01396] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01398] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0139e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h009ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h013fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01400] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01402] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01404] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01406] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01408] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0140e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01410] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01412] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01414] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01416] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01418] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0141e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01420] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01422] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01424] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01426] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01428] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0142e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01430] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01432] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01434] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01436] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01438] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0143e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01440] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01442] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01444] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01446] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01448] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0144e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01450] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01452] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01454] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01456] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01458] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0145e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01460] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01462] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01464] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01466] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01468] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0146e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01470] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01472] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01474] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01476] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01478] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0147e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01480] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01482] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01484] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01486] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01488] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0148e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01490] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01492] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01494] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01496] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01498] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0149e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h014fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01500] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01502] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01504] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01506] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01508] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0150e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01510] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01512] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01514] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01516] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01518] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0151e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01520] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01522] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01524] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01526] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01528] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0152e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01530] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01532] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01534] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01536] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01538] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00a9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0153e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01540] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01542] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01544] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01546] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01548] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0154e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01550] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aa9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01552] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aaa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01554] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01556] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01558] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aaf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0155e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01560] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01562] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01564] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01566] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01568] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0156e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01570] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ab9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01572] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01574] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00abb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01576] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00abc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01578] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00abd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00abe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00abf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0157e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01580] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01582] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01584] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01586] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01588] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0158e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01590] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ac9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01592] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01594] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00acb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01596] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00acc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01598] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00acd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ace] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00acf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0159e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ad9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ada] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00adb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00adc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00add] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ade] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00adf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ae9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aeb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00af9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00afa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00afb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00afc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00afd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00afe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00aff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h015fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01600] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01602] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01604] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01606] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01608] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0160e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01610] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01612] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01614] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01616] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01618] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0161e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01620] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01622] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01624] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01626] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01628] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0162e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01630] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01632] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01634] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01636] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01638] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0163e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01640] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01642] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01644] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01646] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01648] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0164e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01650] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01652] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01654] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01656] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01658] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0165e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01660] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01662] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01664] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01666] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01668] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0166e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01670] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01672] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01674] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01676] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01678] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0167e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01680] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01682] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01684] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01686] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01688] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0168e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01690] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01692] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01694] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01696] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01698] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0169e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h016fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01700] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01702] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01704] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01706] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01708] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0170e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01710] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01712] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01714] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01716] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01718] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0171e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01720] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01722] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01724] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01726] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01728] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0172e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01730] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01732] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01734] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01736] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01738] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00b9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0173e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01740] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01742] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01744] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01746] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01748] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0174e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01750] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ba9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01752] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00baa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01754] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01756] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01758] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00baf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0175e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01760] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01762] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01764] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01766] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01768] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0176e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01770] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bb9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01772] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01774] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bbb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01776] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bbc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01778] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bbd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bbe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bbf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0177e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01780] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01782] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01784] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01786] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01788] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0178e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01790] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bc9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01792] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01794] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bcb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01796] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bcc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01798] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bcd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bcf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0179e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bd9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bdb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bdc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bdd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bde] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bdf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00be9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00beb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bf9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bfa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bfb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bfc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bfd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bfe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00bff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h017fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01800] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01802] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01804] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01806] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01808] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0180e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01810] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01812] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01814] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01816] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01818] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0181e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01820] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01822] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01824] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01826] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01828] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0182e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01830] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01832] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01834] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01836] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01838] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0183e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01840] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01842] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01844] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01846] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01848] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0184e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01850] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01852] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01854] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01856] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01858] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0185e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01860] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01862] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01864] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01866] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01868] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0186e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01870] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01872] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01874] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01876] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01878] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0187e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01880] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01882] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01884] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01886] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01888] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0188e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01890] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01892] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01894] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01896] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01898] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0189e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h018fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01900] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01902] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01904] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01906] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01908] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0190e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01910] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01912] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01914] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01916] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01918] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0191e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01920] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01922] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01924] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01926] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01928] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0192e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01930] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01932] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01934] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01936] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01938] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00c9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0193e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01940] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01942] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01944] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01946] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01948] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0194e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01950] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ca9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01952] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00caa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01954] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01956] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01958] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00caf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0195e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01960] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01962] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01964] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01966] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01968] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0196e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01970] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cb9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01972] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01974] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cbb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01976] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cbc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01978] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cbd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cbe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cbf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0197e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01980] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01982] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01984] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01986] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01988] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0198e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01990] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cc9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01992] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01994] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ccb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01996] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ccc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01998] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ccd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ccf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0199e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cd9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cdb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cdc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cdd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cde] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cdf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ce9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ceb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ced] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cf9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cfa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cfb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cfc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cfd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cfe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00cff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h019fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01a9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aa8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aaa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ab8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01abc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01abe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ac8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01acc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ace] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ad8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ada] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01adc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ade] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ae8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01aee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01af8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01afa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01afc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01afe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00d9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00da9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00daa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00daf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00db9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dbb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dbc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dbd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dbe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dbf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dc9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dcb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dcc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dcd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dcf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01b9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ba8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01baa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dd9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ddb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ddc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ddd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dde] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ddf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00de9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00deb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ded] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00def] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01be8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00df9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dfa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dfb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dfc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bf8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dfd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dfe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00dff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01bfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01c9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ca8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01caa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ccc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ce8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cf8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01cfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00e9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ea9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eaa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ead] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eaf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eb9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ebb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ebc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ebd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ebe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ebf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ec9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ecb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ecc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ecd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ece] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ecf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01d9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01da8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01daa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ed9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00edb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00edc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01db8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00edd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ede] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00edf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ee9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eeb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ddc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01de8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ef9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00efa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00efb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00efc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01df8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00efd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00efe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00eff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01dfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01e9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ea8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eaa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ebc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ebe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ec8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ecc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ece] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ed8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01edc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ede] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ee8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01eee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ef8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01efa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01efc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01efe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00f9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fa9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00faa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00faf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fb9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fbb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fbc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fbd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fbe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fbf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fc9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fcb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fcc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fcd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fcf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01f9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fa8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01faa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fd9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fdb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fdc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fdd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fde] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fdf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fe9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00feb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fe8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01fee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ff9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ffa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ffb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ffc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ff8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ffd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ffa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00ffe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ffc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h00fff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h01ffe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01000] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02000] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01001] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02002] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01002] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02004] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01003] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02006] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01004] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02008] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01005] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01006] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01007] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0200e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01008] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02010] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01009] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02012] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02014] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02016] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02018] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0100f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0201e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01010] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02020] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01011] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02022] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01012] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02024] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01013] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02026] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01014] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02028] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01015] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01016] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01017] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0202e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01018] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02030] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01019] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02032] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02034] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02036] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02038] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0101f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0203e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01020] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02040] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01021] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02042] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01022] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02044] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01023] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02046] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01024] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02048] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01025] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01026] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01027] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0204e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01028] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02050] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01029] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02052] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02054] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02056] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02058] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0102f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0205e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01030] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02060] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01031] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02062] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01032] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02064] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01033] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02066] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01034] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02068] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01035] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01036] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01037] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0206e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01038] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02070] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01039] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02072] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02074] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02076] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02078] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0103f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0207e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01040] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02080] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01041] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02082] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01042] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02084] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01043] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02086] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01044] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02088] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01045] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01046] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01047] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0208e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01048] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02090] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01049] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02092] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02094] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02096] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02098] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0104f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0209e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01050] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01051] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01052] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01053] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01054] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01055] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01056] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01057] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01058] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01059] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0105f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01060] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01061] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01062] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01063] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01064] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01065] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01066] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01067] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01068] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01069] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0106f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01070] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01071] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01072] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01073] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01074] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01075] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01076] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01077] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01078] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01079] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0107f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h020fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01080] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02100] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01081] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02102] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01082] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02104] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01083] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02106] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01084] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02108] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01085] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01086] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01087] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0210e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01088] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02110] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01089] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02112] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02114] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02116] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02118] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0108f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0211e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01090] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02120] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01091] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02122] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01092] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02124] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01093] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02126] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01094] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02128] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01095] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01096] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01097] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0212e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01098] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02130] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01099] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02132] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02134] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02136] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02138] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0109f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0213e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02140] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02142] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02144] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02146] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02148] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0214e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02150] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02152] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02154] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02156] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02158] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0215e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02160] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02162] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02164] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02166] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02168] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0216e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02170] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02172] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02174] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02176] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02178] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0217e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02180] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02182] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02184] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02186] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02188] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0218e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02190] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02192] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02194] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02196] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02198] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0219e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h010ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h021fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01100] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02200] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01101] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02202] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01102] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02204] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01103] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02206] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01104] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02208] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01105] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01106] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01107] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0220e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01108] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02210] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01109] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02212] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02214] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02216] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02218] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0110f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0221e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01110] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02220] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01111] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02222] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01112] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02224] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01113] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02226] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01114] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02228] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01115] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01116] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01117] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0222e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01118] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02230] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01119] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02232] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02234] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02236] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02238] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0111f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0223e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01120] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02240] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01121] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02242] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01122] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02244] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01123] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02246] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01124] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02248] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01125] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01126] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01127] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0224e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01128] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02250] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01129] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02252] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02254] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02256] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02258] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0112f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0225e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01130] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02260] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01131] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02262] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01132] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02264] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01133] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02266] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01134] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02268] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01135] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01136] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01137] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0226e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01138] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02270] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01139] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02272] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02274] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02276] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02278] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0113f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0227e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01140] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02280] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01141] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02282] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01142] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02284] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01143] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02286] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01144] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02288] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01145] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01146] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01147] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0228e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01148] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02290] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01149] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02292] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02294] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02296] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02298] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0114f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0229e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01150] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01151] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01152] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01153] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01154] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01155] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01156] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01157] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01158] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01159] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0115f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01160] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01161] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01162] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01163] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01164] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01165] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01166] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01167] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01168] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01169] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0116f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01170] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01171] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01172] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01173] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01174] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01175] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01176] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01177] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01178] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01179] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0117f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h022fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01180] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02300] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01181] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02302] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01182] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02304] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01183] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02306] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01184] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02308] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01185] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01186] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01187] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0230e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01188] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02310] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01189] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02312] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02314] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02316] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02318] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0118f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0231e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01190] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02320] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01191] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02322] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01192] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02324] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01193] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02326] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01194] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02328] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01195] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01196] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01197] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0232e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01198] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02330] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01199] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02332] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02334] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02336] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02338] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0119f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0233e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02340] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02342] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02344] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02346] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02348] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0234e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02350] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02352] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02354] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02356] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02358] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0235e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02360] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02362] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02364] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02366] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02368] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0236e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02370] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02372] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02374] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02376] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02378] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0237e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02380] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02382] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02384] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02386] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02388] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0238e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02390] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02392] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02394] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02396] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02398] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0239e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h011ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h023fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01200] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02400] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01201] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02402] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01202] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02404] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01203] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02406] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01204] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02408] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01205] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01206] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01207] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0240e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01208] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02410] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01209] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02412] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02414] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02416] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02418] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0120f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0241e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01210] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02420] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01211] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02422] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01212] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02424] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01213] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02426] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01214] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02428] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01215] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01216] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01217] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0242e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01218] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02430] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01219] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02432] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02434] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02436] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02438] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0121f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0243e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01220] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02440] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01221] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02442] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01222] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02444] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01223] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02446] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01224] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02448] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01225] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01226] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01227] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0244e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01228] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02450] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01229] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02452] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02454] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02456] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02458] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0122f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0245e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01230] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02460] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01231] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02462] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01232] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02464] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01233] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02466] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01234] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02468] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01235] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01236] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01237] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0246e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01238] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02470] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01239] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02472] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02474] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02476] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02478] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0123f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0247e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01240] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02480] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01241] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02482] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01242] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02484] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01243] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02486] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01244] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02488] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01245] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01246] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01247] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0248e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01248] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02490] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01249] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02492] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02494] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02496] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02498] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0124f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0249e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01250] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01251] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01252] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01253] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01254] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01255] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01256] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01257] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01258] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01259] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0125f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01260] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01261] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01262] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01263] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01264] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01265] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01266] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01267] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01268] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01269] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0126f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01270] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01271] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01272] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01273] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01274] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01275] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01276] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01277] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01278] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01279] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0127f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h024fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01280] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02500] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01281] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02502] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01282] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02504] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01283] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02506] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01284] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02508] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01285] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01286] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01287] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0250e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01288] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02510] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01289] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02512] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02514] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02516] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02518] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0128f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0251e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01290] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02520] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01291] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02522] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01292] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02524] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01293] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02526] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01294] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02528] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01295] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01296] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01297] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0252e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01298] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02530] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01299] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02532] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02534] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02536] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02538] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0129f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0253e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02540] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02542] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02544] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02546] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02548] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0254e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02550] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02552] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02554] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02556] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02558] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0255e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02560] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02562] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02564] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02566] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02568] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0256e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02570] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02572] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02574] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02576] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02578] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0257e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02580] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02582] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02584] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02586] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02588] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0258e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02590] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02592] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02594] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02596] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02598] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0259e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h012ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h025fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01300] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02600] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01301] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02602] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01302] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02604] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01303] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02606] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01304] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02608] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01305] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01306] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01307] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0260e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01308] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02610] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01309] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02612] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02614] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02616] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02618] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0130f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0261e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01310] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02620] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01311] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02622] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01312] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02624] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01313] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02626] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01314] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02628] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01315] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01316] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01317] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0262e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01318] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02630] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01319] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02632] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02634] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02636] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02638] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0131f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0263e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01320] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02640] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01321] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02642] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01322] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02644] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01323] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02646] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01324] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02648] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01325] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01326] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01327] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0264e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01328] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02650] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01329] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02652] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02654] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02656] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02658] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0132f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0265e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01330] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02660] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01331] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02662] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01332] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02664] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01333] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02666] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01334] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02668] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01335] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01336] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01337] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0266e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01338] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02670] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01339] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02672] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02674] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02676] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02678] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0133f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0267e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01340] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02680] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01341] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02682] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01342] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02684] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01343] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02686] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01344] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02688] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01345] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01346] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01347] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0268e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01348] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02690] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01349] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02692] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02694] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02696] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02698] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0134f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0269e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01350] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01351] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01352] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01353] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01354] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01355] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01356] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01357] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01358] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01359] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0135f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01360] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01361] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01362] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01363] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01364] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01365] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01366] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01367] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01368] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01369] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0136f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01370] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01371] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01372] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01373] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01374] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01375] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01376] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01377] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01378] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01379] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0137f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h026fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01380] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02700] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01381] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02702] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01382] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02704] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01383] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02706] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01384] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02708] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01385] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01386] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01387] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0270e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01388] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02710] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01389] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02712] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02714] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02716] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02718] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0138f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0271e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01390] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02720] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01391] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02722] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01392] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02724] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01393] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02726] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01394] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02728] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01395] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01396] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01397] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0272e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01398] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02730] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01399] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02732] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02734] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02736] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02738] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0139f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0273e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02740] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02742] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02744] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02746] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02748] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0274e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02750] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02752] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02754] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02756] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02758] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0275e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02760] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02762] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02764] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02766] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02768] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0276e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02770] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02772] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02774] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02776] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02778] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0277e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02780] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02782] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02784] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02786] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02788] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0278e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02790] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02792] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02794] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02796] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02798] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0279e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h013ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h027fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01400] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02800] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01401] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02802] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01402] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02804] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01403] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02806] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01404] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02808] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01405] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01406] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01407] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0280e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01408] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02810] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01409] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02812] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02814] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02816] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02818] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0140f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0281e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01410] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02820] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01411] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02822] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01412] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02824] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01413] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02826] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01414] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02828] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01415] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01416] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01417] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0282e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01418] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02830] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01419] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02832] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02834] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02836] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02838] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0141f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0283e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01420] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02840] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01421] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02842] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01422] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02844] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01423] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02846] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01424] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02848] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01425] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01426] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01427] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0284e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01428] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02850] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01429] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02852] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02854] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02856] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02858] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0142f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0285e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01430] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02860] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01431] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02862] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01432] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02864] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01433] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02866] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01434] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02868] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01435] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01436] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01437] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0286e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01438] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02870] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01439] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02872] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02874] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02876] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02878] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0143f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0287e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01440] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02880] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01441] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02882] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01442] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02884] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01443] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02886] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01444] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02888] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01445] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01446] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01447] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0288e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01448] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02890] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01449] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02892] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02894] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02896] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02898] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0144f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0289e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01450] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01451] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01452] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01453] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01454] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01455] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01456] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01457] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01458] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01459] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0145f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01460] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01461] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01462] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01463] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01464] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01465] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01466] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01467] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01468] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01469] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0146f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01470] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01471] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01472] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01473] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01474] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01475] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01476] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01477] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01478] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01479] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0147f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h028fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01480] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02900] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01481] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02902] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01482] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02904] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01483] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02906] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01484] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02908] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01485] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01486] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01487] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0290e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01488] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02910] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01489] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02912] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02914] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02916] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02918] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0148f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0291e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01490] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02920] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01491] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02922] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01492] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02924] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01493] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02926] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01494] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02928] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01495] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01496] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01497] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0292e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01498] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02930] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01499] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02932] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02934] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02936] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02938] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0149f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0293e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02940] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02942] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02944] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02946] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02948] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0294e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02950] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02952] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02954] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02956] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02958] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0295e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02960] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02962] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02964] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02966] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02968] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0296e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02970] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02972] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02974] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02976] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02978] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0297e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02980] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02982] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02984] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02986] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02988] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0298e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02990] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02992] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02994] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02996] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02998] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0299e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h014ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h029fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01500] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01501] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01502] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01503] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01504] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01505] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01506] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01507] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01508] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01509] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0150f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01510] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01511] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01512] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01513] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01514] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01515] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01516] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01517] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01518] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01519] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0151f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01520] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01521] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01522] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01523] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01524] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01525] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01526] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01527] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01528] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01529] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0152f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01530] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01531] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01532] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01533] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01534] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01535] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01536] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01537] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01538] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01539] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0153f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01540] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01541] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01542] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01543] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01544] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01545] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01546] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01547] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01548] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01549] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0154f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02a9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01550] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01551] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01552] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01553] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01554] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aa8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01555] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aaa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01556] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01557] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01558] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01559] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ab8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02abc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0155f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02abe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01560] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01561] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01562] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01563] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01564] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ac8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01565] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01566] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02acc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01567] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ace] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01568] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01569] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ad8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ada] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02adc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0156f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ade] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01570] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01571] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01572] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01573] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01574] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ae8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01575] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01576] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01577] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02aee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01578] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01579] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02af8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02afa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02afc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0157f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02afe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01580] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01581] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01582] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01583] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01584] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01585] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01586] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01587] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01588] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01589] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0158f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01590] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01591] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01592] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01593] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01594] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01595] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01596] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01597] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01598] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01599] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0159f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02b9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ba8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02baa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02be8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bf8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h015ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02bfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01600] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01601] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01602] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01603] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01604] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01605] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01606] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01607] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01608] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01609] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0160f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01610] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01611] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01612] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01613] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01614] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01615] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01616] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01617] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01618] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01619] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0161f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01620] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01621] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01622] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01623] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01624] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01625] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01626] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01627] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01628] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01629] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0162f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01630] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01631] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01632] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01633] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01634] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01635] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01636] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01637] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01638] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01639] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0163f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01640] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01641] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01642] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01643] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01644] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01645] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01646] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01647] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01648] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01649] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0164f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02c9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01650] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01651] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01652] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01653] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01654] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ca8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01655] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02caa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01656] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01657] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01658] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01659] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0165f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01660] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01661] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01662] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01663] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01664] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01665] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01666] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ccc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01667] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01668] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01669] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0166f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01670] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01671] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01672] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01673] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01674] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ce8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01675] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01676] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01677] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01678] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01679] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cf8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0167f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02cfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01680] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01681] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01682] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01683] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01684] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01685] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01686] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01687] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01688] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01689] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0168f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01690] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01691] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01692] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01693] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01694] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01695] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01696] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01697] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01698] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01699] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0169f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02d9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02da8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02daa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02db8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ddc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02de8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02df8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h016ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02dfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01700] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01701] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01702] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01703] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01704] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01705] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01706] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01707] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01708] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01709] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0170f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01710] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01711] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01712] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01713] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01714] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01715] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01716] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01717] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01718] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01719] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0171f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01720] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01721] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01722] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01723] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01724] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01725] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01726] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01727] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01728] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01729] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0172f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01730] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01731] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01732] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01733] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01734] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01735] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01736] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01737] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01738] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01739] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0173f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01740] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01741] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01742] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01743] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01744] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01745] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01746] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01747] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01748] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01749] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0174f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02e9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01750] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01751] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01752] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01753] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01754] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ea8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01755] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eaa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01756] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01757] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01758] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01759] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ebc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0175f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ebe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01760] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01761] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01762] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01763] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01764] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ec8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01765] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01766] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ecc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01767] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ece] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01768] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01769] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ed8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02edc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0176f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ede] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01770] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01771] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01772] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01773] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01774] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ee8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01775] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01776] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01777] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02eee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01778] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01779] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ef8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02efa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02efc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0177f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02efe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01780] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01781] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01782] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01783] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01784] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01785] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01786] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01787] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01788] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01789] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0178f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01790] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01791] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01792] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01793] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01794] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01795] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01796] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01797] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01798] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01799] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0179f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02f9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fa8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02faa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fe8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02fee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ff8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ffa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ffc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h017ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h02ffe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01800] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03000] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01801] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03002] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01802] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03004] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01803] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03006] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01804] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03008] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01805] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01806] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01807] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0300e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01808] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03010] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01809] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03012] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03014] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03016] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03018] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0180f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0301e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01810] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03020] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01811] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03022] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01812] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03024] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01813] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03026] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01814] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03028] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01815] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01816] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01817] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0302e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01818] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03030] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01819] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03032] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03034] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03036] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03038] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0181f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0303e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01820] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03040] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01821] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03042] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01822] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03044] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01823] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03046] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01824] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03048] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01825] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01826] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01827] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0304e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01828] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03050] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01829] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03052] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03054] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03056] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03058] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0182f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0305e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01830] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03060] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01831] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03062] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01832] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03064] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01833] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03066] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01834] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03068] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01835] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01836] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01837] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0306e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01838] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03070] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01839] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03072] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03074] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03076] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03078] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0183f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0307e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01840] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03080] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01841] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03082] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01842] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03084] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01843] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03086] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01844] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03088] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01845] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01846] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01847] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0308e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01848] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03090] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01849] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03092] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03094] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03096] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03098] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0184f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0309e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01850] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01851] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01852] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01853] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01854] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01855] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01856] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01857] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01858] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01859] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0185f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01860] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01861] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01862] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01863] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01864] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01865] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01866] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01867] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01868] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01869] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0186f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01870] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01871] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01872] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01873] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01874] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01875] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01876] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01877] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01878] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01879] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0187f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h030fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01880] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03100] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01881] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03102] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01882] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03104] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01883] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03106] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01884] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03108] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01885] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01886] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01887] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0310e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01888] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03110] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01889] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03112] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03114] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03116] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03118] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0188f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0311e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01890] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03120] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01891] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03122] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01892] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03124] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01893] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03126] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01894] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03128] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01895] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01896] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01897] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0312e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01898] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03130] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01899] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03132] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03134] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03136] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03138] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0189f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0313e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03140] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03142] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03144] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03146] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03148] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0314e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03150] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03152] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03154] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03156] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03158] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0315e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03160] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03162] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03164] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03166] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03168] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0316e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03170] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03172] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03174] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03176] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03178] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0317e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03180] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03182] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03184] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03186] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03188] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0318e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03190] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03192] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03194] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03196] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03198] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0319e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h018ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h031fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01900] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03200] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01901] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03202] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01902] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03204] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01903] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03206] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01904] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03208] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01905] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01906] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01907] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0320e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01908] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03210] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01909] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03212] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03214] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03216] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03218] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0190f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0321e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01910] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03220] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01911] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03222] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01912] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03224] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01913] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03226] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01914] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03228] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01915] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01916] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01917] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0322e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01918] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03230] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01919] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03232] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03234] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03236] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03238] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0191f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0323e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01920] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03240] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01921] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03242] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01922] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03244] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01923] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03246] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01924] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03248] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01925] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01926] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01927] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0324e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01928] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03250] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01929] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03252] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03254] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03256] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03258] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0192f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0325e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01930] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03260] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01931] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03262] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01932] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03264] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01933] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03266] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01934] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03268] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01935] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01936] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01937] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0326e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01938] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03270] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01939] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03272] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03274] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03276] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03278] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0193f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0327e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01940] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03280] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01941] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03282] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01942] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03284] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01943] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03286] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01944] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03288] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01945] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01946] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01947] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0328e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01948] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03290] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01949] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03292] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03294] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03296] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03298] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0194f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0329e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01950] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01951] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01952] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01953] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01954] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01955] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01956] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01957] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01958] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01959] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0195f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01960] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01961] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01962] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01963] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01964] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01965] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01966] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01967] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01968] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01969] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0196f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01970] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01971] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01972] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01973] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01974] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01975] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01976] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01977] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01978] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01979] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0197f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h032fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01980] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03300] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01981] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03302] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01982] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03304] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01983] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03306] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01984] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03308] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01985] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01986] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01987] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0330e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01988] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03310] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01989] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03312] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03314] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03316] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03318] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0198f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0331e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01990] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03320] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01991] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03322] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01992] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03324] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01993] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03326] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01994] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03328] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01995] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01996] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01997] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0332e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01998] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03330] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01999] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03332] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03334] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03336] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03338] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h0199f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0333e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03340] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03342] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03344] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03346] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03348] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0334e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03350] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019a9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03352] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019aa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03354] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03356] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03358] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019af] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0335e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03360] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03362] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03364] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03366] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03368] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0336e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03370] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019b9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03372] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03374] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019bb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03376] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019bc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03378] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019bd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019be] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019bf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0337e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03380] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03382] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03384] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03386] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03388] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0338e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03390] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019c9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03392] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03394] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019cb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03396] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019cc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03398] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019cd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019cf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0339e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019d9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019da] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019db] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019dc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019dd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019de] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019df] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019e9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019eb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019f9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019fa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019fb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019fc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019fd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019fe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h019ff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h033fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03400] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03402] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03404] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03406] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03408] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0340e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03410] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03412] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03414] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03416] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03418] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0341e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03420] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03422] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03424] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03426] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03428] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0342e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03430] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03432] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03434] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03436] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03438] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0343e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03440] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03442] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03444] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03446] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03448] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0344e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03450] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03452] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03454] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03456] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03458] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0345e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03460] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03462] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03464] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03466] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03468] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0346e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03470] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03472] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03474] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03476] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03478] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0347e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03480] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03482] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03484] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03486] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03488] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0348e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03490] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03492] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03494] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03496] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03498] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0349e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h034fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03500] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03502] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03504] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03506] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03508] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0350e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03510] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03512] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03514] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03516] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03518] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0351e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03520] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03522] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03524] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03526] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03528] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0352e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03530] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03532] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03534] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03536] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03538] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01a9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0353e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03540] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03542] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03544] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03546] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03548] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0354e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03550] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aa9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03552] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aaa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03554] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03556] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03558] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aaf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0355e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03560] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03562] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03564] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03566] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03568] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0356e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03570] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ab9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03572] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03574] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01abb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03576] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01abc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03578] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01abd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01abe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01abf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0357e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03580] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03582] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03584] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03586] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03588] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0358e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03590] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ac9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03592] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03594] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01acb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03596] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01acc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03598] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01acd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ace] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01acf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0359e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ad9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ada] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01adb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01adc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01add] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ade] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01adf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ae9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aeb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01af9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01afa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01afb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01afc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01afd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01afe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01aff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h035fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03600] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03602] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03604] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03606] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03608] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0360e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03610] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03612] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03614] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03616] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03618] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0361e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03620] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03622] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03624] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03626] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03628] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0362e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03630] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03632] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03634] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03636] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03638] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0363e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03640] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03642] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03644] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03646] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03648] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0364e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03650] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03652] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03654] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03656] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03658] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0365e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03660] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03662] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03664] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03666] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03668] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0366e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03670] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03672] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03674] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03676] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03678] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0367e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03680] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03682] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03684] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03686] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03688] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0368e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03690] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03692] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03694] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03696] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03698] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0369e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h036fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03700] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03702] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03704] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03706] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03708] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0370e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03710] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03712] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03714] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03716] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03718] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0371e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03720] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03722] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03724] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03726] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03728] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0372e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03730] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03732] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03734] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03736] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03738] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01b9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0373e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03740] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03742] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03744] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03746] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03748] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0374e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03750] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ba9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03752] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01baa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03754] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03756] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03758] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01baf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0375e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03760] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03762] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03764] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03766] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03768] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0376e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03770] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bb9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03772] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03774] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bbb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03776] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bbc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03778] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bbd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bbe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bbf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0377e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03780] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03782] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03784] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03786] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03788] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0378e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03790] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bc9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03792] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03794] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bcb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03796] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bcc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03798] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bcd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bcf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0379e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bd9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bdb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bdc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bdd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bde] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bdf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01be9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01beb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bf9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bfa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bfb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bfc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bfd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bfe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01bff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h037fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03800] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03802] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03804] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03806] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03808] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0380e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03810] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03812] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03814] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03816] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03818] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0381e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03820] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03822] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03824] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03826] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03828] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0382e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03830] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03832] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03834] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03836] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03838] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0383e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03840] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03842] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03844] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03846] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03848] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0384e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03850] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03852] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03854] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03856] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03858] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0385e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03860] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03862] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03864] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03866] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03868] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0386e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03870] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03872] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03874] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03876] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03878] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0387e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03880] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03882] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03884] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03886] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03888] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0388e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03890] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03892] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03894] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03896] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03898] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0389e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h038fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03900] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03902] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03904] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03906] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03908] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0390e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03910] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03912] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03914] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03916] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03918] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0391e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03920] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03922] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03924] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03926] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03928] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0392e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03930] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03932] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03934] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03936] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03938] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01c9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0393e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03940] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03942] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03944] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03946] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03948] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0394e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03950] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ca9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03952] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01caa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03954] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03956] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03958] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01caf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0395e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03960] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03962] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03964] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03966] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03968] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0396e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03970] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cb9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03972] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03974] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cbb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03976] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cbc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03978] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cbd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cbe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cbf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0397e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03980] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03982] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03984] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03986] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03988] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0398e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03990] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cc9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03992] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03994] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ccb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03996] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ccc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03998] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ccd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ccf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h0399e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039a8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039aa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cd9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cdb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cdc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039b8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cdd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cde] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039bc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cdf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039be] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039c8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039cc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ce9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ceb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039d8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ced] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039da] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039dc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039de] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039e8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039ee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cf9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cfa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cfb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cfc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039f8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cfd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039fa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cfe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039fc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01cff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h039fe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03a9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aa8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aaa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ab8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03abc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03abe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ac8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03acc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ace] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ad8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ada] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03adc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ade] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ae8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03aee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03af8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03afa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03afc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03afe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01d9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01da9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01daa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01daf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01db9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dbb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dbc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dbd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dbe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dbf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dc9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dcb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dcc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dcd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dcf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03b9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ba8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03baa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dd9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ddb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ddc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ddd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dde] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ddf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01de9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01deb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ded] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01def] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03be8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01df9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dfa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dfb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dfc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bf8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dfd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dfe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01dff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03bfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03c9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ca8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03caa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ccc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ce8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cf8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03cfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01e9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ea9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eaa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ead] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eaf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eb9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ebb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ebc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ebd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ebe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ebf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ec9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ecb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ecc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ecd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ece] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ecf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03d9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03da8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03daa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ed9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01edb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01edc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03db8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01edd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ede] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01edf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ee9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eeb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ddc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03de8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ef9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01efa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01efb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01efc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03df8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01efd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dfa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01efe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dfc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01eff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03dfe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f00] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f01] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f02] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f03] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f04] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f05] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f06] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f07] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f08] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f09] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f0f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f10] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f11] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f12] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f13] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f14] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f15] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f16] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f17] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f18] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f19] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f1f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f20] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f21] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f22] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f23] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f24] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f25] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f26] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f27] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f28] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f29] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f2f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f30] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f31] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f32] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f33] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f34] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f35] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f36] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f37] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f38] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f39] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f3f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f40] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f41] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f42] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f43] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f44] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f45] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f46] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f47] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f48] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f49] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f4f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03e9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f50] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f51] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f52] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f53] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f54] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ea8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f55] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eaa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f56] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f57] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f58] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f59] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ebc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f5f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ebe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f60] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f61] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f62] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f63] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f64] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ec8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f65] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f66] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ecc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f67] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ece] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f68] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f69] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ed8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03edc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f6f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ede] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f70] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f71] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f72] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f73] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f74] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ee8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f75] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f76] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f77] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03eee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f78] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f79] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ef8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03efa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03efc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f7f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03efe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f80] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f00] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f81] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f02] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f82] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f04] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f83] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f06] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f84] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f08] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f85] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f86] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f87] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f0e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f88] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f10] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f89] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f12] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f14] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f16] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f18] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f8f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f1e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f90] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f20] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f91] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f22] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f92] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f24] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f93] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f26] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f94] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f28] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f95] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f96] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f97] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f2e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f98] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f30] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f99] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f32] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9a] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f34] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9b] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f36] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9c] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f38] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9d] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9e] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01f9f] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f3e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f40] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f42] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f44] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f46] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f48] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f4e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f50] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fa9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f52] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01faa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f54] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fab] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f56] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fac] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f58] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fad] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fae] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01faf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f5e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f60] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f62] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f64] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f66] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f68] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f6e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f70] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fb9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f72] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fba] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f74] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fbb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f76] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fbc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f78] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fbd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fbe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fbf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f7e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f80] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f82] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f84] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f86] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f88] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f8e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f90] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fc9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f92] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fca] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f94] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fcb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f96] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fcc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f98] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fcd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9a] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fce] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9c] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fcf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03f9e] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fa8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03faa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fac] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fae] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fd9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fda] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fdb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fdc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fb8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fdd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fba] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fde] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fbc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fdf] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fbe] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fc8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fca] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fcc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fce] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fe9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fea] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01feb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fec] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fd8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fed] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fda] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fee] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fdc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fef] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fde] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff0] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff1] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff2] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff3] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff4] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fe8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff5] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fea] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff6] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fec] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff7] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03fee] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff8] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff0] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ff9] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff2] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ffa] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff4] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ffb] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff6] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ffc] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ff8] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ffd] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ffa] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01ffe] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ffc] ;
//end
//always_comb begin // 
               I1b5811486f7a6670fb1b4d36b84beb7b32860428e990713b5714655ff65df1f2['h01fff] =  Ieafd9525846c58bc50d97b888c56259ef9df96a08d8897927069698b763f4748['h03ffe] ;
//end
