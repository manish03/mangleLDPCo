 reg  ['hfff:0] [$clog2('h7000+1)-1:0] I1b23c494e0c04cc5a8a3ff99b6cdf26d ;
