         I0c1c52a843a5de4bb5e0eb6897ea37c4 =   'h00380 ;
         Ice4c8b10e41f361db2bd4a7b8470b05e =   'h0013a ;
         I612d62c35e606e6e91220910fd8448f1 =   'h0010b ;
         I4f664d460f924a71ebd3cc05f0916521 =   'h000f1 ;
         I0e38bd43118f53204e169f324066b75c =   'h000de ;
         I46878ad6c93d318bf7a959c78090bf66 =   'h000d0 ;
         Ie2c597c226457d94ec76f1513d95aab2 =   'h000c4 ;
         I2c72e48d1e2274c662c18b729af96161 =   'h000ba ;
         Id416e2e4f204401c79d97ae6ae1414ae =   'h000b2 ;
         I8fa96c5580fd6050e2a8c5fcb77c9927 =   'h000aa ;
         Ia9569f758e6bc743aae3a2bb51d941ee =   'h000a3 ;
         I00ae3aaf6b44b2f7fd9bbceafb9c4e22 =   'h0009d ;
         Ibfea7f98ec3bbe5588eb75cbcef739d7 =   'h00098 ;
         Id9eff948ed9da8502308740b4ae17dbf =   'h00093 ;
         If9d08c27c57ed8293171486ad65ed95c =   'h0008e ;
         Iace1409bfc12437ef093b91d50c8175a =   'h0008a ;
         I506d9cf5c368c130a8517f994e7f7a43 =   'h00085 ;
         I0f3fb929c6ee46d33daeba7024107aff =   'h00082 ;
         Id3ac7026a6f63b1dc8588f9bdfd50068 =   'h0007e ;
         I680caae24965f4516cbd8642d4d43b3b =   'h0007b ;
         I7b240e087870bef3e01b2de04cdbae13 =   'h00077 ;
         Ic2b7c4749006adaa1dfa0ca1c5d7a371 =   'h00074 ;
         I2abc1d3ddcecbdbdc971abb93be58744 =   'h00071 ;
         I9fcc49fa3eb8ad62633822ff3ac5973a =   'h0006f ;
         I6b938059b8a71491bf1718326233b688 =   'h0006c ;
         I5d98a20b0eef6a335b29f017cd3120df =   'h00069 ;
         I69d5314c6ba43f6d015acf00c8a2a7be =   'h00067 ;
         I64ce8a8f7f046222c963820f37362021 =   'h00065 ;
         I4e1c98665268d59e19c3068ff9efe9a8 =   'h00062 ;
         I1399a46a42c2cc384efc8ca681b1b249 =   'h00060 ;
         I3e0d577c49e0fcba84112e3afab2edbe =   'h0005e ;
         Ic266aa3f20103455635f801a0fe1056a =   'h0005c ;
         I285c0d0dbcb505b98bbf005805067396 =   'h0005a ;
         Icba253e44f98c391c02e864856715f49 =   'h00058 ;
         Iaa4b6b01007d9836ae0092101c4065db =   'h00056 ;
         Ia2f4d61e666ea4e0d8085325cdaa7344 =   'h00055 ;
         I84ed644f3578e53744802bab05d17011 =   'h00053 ;
         I5fbdad2d56ab8f5435a712b512190645 =   'h00051 ;
         I670a7cf3b4948b0d31c871ba641af4c1 =   'h00050 ;
         I227702af9307eb6600ed78a648bb71e9 =   'h0004e ;
         If0c4078bb97b3a246a91be4180ee7af9 =   'h0004c ;
         I913f1af34aaf3d51d3c60489979a81d5 =   'h0004b ;
         I22e712371781d71cbb80680359ccd708 =   'h0004a ;
         I5e9450b27761da0b895a4f6ace1ad171 =   'h00048 ;
         I0b1bc20ea62f64bae807d8ac1166139f =   'h00047 ;
         Idddfbcad405258a5434d8b94eb26654c =   'h00045 ;
         I8beef0ea5356b2f46d7d5f16db49ebef =   'h00044 ;
         I499586880161ca66628afed78e7e495d =   'h00043 ;
         Ie909ad4a9ba2fde8fd6451e7eda2088d =   'h00042 ;
         Iee75fb439b2200aba94b03fd69cd7adc =   'h00040 ;
         Id8a8555f4bf9003a0ac0dcafaa67e68d =   'h0003f ;
         I10065fe206e6700159260af61afa61c2 =   'h0003e ;
         Ia41593b7790fde4ae4dd986dd583286f =   'h0003d ;
         I44490a711aece8f1a24c080cd0f37607 =   'h0003c ;
         Ic35377a5686c5a6edace93b58129cbdd =   'h0003b ;
         Iccd1e1793be28ddad794782e2700a4d0 =   'h0003a ;
         Id112833f079dcf6e092d48cd13120d47 =   'h00039 ;
         Ia550c5040df02dc8a8735562e71ddf6f =   'h00038 ;
         Ibcaed8bfefd254ded778d760cd533b81 =   'h00037 ;
         I19c7906957daf8e2a04b013e95db9c6e =   'h00036 ;
         I4bbddbcd811dc6936fd20d18559e3aac =   'h00035 ;
         Idaf09a27ce68e8877da2d4c48be4c8ca =   'h00034 ;
         I82ad270d36061ef06232de9b92742dfd =   'h00033 ;
         Ieb5d1ef84057ceba02d9db624be39285 =   'h00032 ;
         I7ebd34e6a95c3589b44cc0941f54bfa9 =   'h00031 ;
         I46432f8bb8f39efef70554ea0e8573de =   'h00031 ;
         I1fb7b6a528ec8d5871cb15a490bbfda2 =   'h00030 ;
         I25d429f4a9f397a0d0ca515241b3c1b5 =   'h0002f ;
         I3ca008900582aea13c5cf09b6c3af78e =   'h0002e ;
         Id9a5e1c4a044b3006d620dd52e2e8ddc =   'h0002d ;
         I63f34eddeedc5ded8721b40546c758c3 =   'h0002d ;
         I8ec5f00523507f51358081e52a5bc55c =   'h0002c ;
         Ib77465ae19c99c6e2c39e2ab6438730d =   'h0002b ;
         I025a54040366d4505896c1179d580dc1 =   'h0002a ;
         I0ac7e4f7f0e68450455e4a3d3ed57c56 =   'h0002a ;
         If6f5c61447dbeeaef688c670c9802649 =   'h00029 ;
         I968168f5cd481033283f24425f7862b9 =   'h00028 ;
         Ie364b2799febe180ea9c2361279bcdc3 =   'h00028 ;
         I76cc2a7d1f750a49780fe7e7f1651d5e =   'h00027 ;
         I2e3ac4cb975151fcb26d716ef80a24f9 =   'h00026 ;
         I6da8878ff3f8680907597ba4ab49e7e4 =   'h00026 ;
         I28db3b4aa4f26a48ef6a28956536d15a =   'h00025 ;
         I7b95e7f8f8f6d01ad095fdfbe36e7f6d =   'h00025 ;
         Ieb56b02269e16c20b5f626afc1b97c98 =   'h00024 ;
         I486565b0e63446c0b122a62bac6644da =   'h00023 ;
         Ibd4082b5df0c5bca554397e77fbf589e =   'h00023 ;
         I6361b4f6c6266288a5f53dfbf0e514cc =   'h00022 ;
         I0590fa4c4cb5194e038b57fd416210b9 =   'h00022 ;
         If8409ca3930cc882752b4efe399aa107 =   'h00021 ;
         I509f64436f6d698c58fa255372adf7e7 =   'h00021 ;
         Ib6319f6f8e74409bd60d624b07fc75d2 =   'h00020 ;
         I344f88b13d6f536724dd33ed2d9fa07a =   'h00020 ;
         Ia9c1251bf7d48ef32d67ee176ca55e07 =   'h0001f ;
         I8a885ced1613614d0bc3e1d2ce31cd34 =   'h0001e ;
         I084e8923b177a76c4fbed301ae5f905f =   'h0001e ;
         I58d2c7aa1ec77bc041b6b1e2e4ad8277 =   'h0001e ;
         I9be477a653c8d0bd98ea404fa8876dd5 =   'h0001d ;
         Ifefb2b21271a5578ec1e1d9ddae2047c =   'h0001d ;
         I708bb50785dd2710e712438dcfec5eb1 =   'h0001c ;
         I12e20bdca30dd5a4695333353faaafe1 =   'h0001c ;
         I37da1f9f97e273359be9e4912f8a8ee7 =   'h0001b ;
         I0df8e26f5e3a60744a02e8b50cff23a5 =   'h0001b ;
         I0f005326cad2001188a9fc4b919bd19a =   'h0001a ;
         I1b7f0cb10a2a1c63083aa2e5d5fe84d8 =   'h0001a ;
         I43240748b90a2f1b2738d7773256f36c =   'h0001a ;
         I9d301fb4da56021d4bf0df8dd2719eb4 =   'h00019 ;
         I50188fbeeabb5bbc1549229769cc58d3 =   'h00019 ;
         I85af941bfb4adc588579de64e51887bb =   'h00018 ;
         I6baa38fdfb9b81d807b09ca3b7cd5d32 =   'h00018 ;
         Ica83cfc4696601a6936e577389a395cc =   'h00018 ;
         I9ae9897faacb46733dcec0b985a590ce =   'h00017 ;
         Ibcf6f538d26631634b6ceafdd3ee991f =   'h00017 ;
         Ia2d7c7007306e7b2ca65518fcc005588 =   'h00016 ;
         I5db8abcf5c9f55ffbe360502c0acf592 =   'h00016 ;
         Iebf161a4f32971bd911356670349e894 =   'h00016 ;
         Iba78cb5ab1da071088bf8f924095d1dd =   'h00015 ;
         Ib8bc0d119e76d93a801d9749ff205d30 =   'h00015 ;
         I7d760437e7830701c90db6653febff5a =   'h00015 ;
         Ie7d3e4264ef52d194bcd054dc421e97e =   'h00014 ;
         I2271582af0c776dadff851456aa6e4a7 =   'h00014 ;
         I851e3c75bf75803e1d745053721aa9ad =   'h00014 ;
         Ifa32facd628d97fa55482c63464bbeed =   'h00013 ;
         I37a83fa1dac26d4614760db718790dfb =   'h00013 ;
         Icdfa771d45c36fef80efda13b0481130 =   'h00013 ;
         Ic72a44c59c204b5d5b77523429df133b =   'h00013 ;
         I1395b926b6d89fdfe41444e3a94d0d10 =   'h00012 ;
         I8393828bf7f4ce64ef97785fcd0d65fb =   'h00012 ;
         I2f6dc9f6f5d1316b9426bbe277b82427 =   'h00012 ;
         I60098787140a26167a69e135e08c6e8b =   'h00011 ;
         Ice5b808b49ac5331f4fd6f36e74f0897 =   'h00011 ;
         I3480a29289d8eca6cbf762b798ec68fc =   'h00011 ;
         Ie8718369d950a31dd1e9b307ce68984c =   'h00011 ;
         I954ad53f646754aa0c8db5073aff65fe =   'h00010 ;
         I8f9194a8b73a5008a74dfe09429e455b =   'h00010 ;
         I9b0851ae1b88864bd086003066137b86 =   'h00010 ;
         Ia8d552e62e3c642796936c2c4188f8a4 =   'h00010 ;
         Idaffd115023b38f3f7e7cafe8e2cedb8 =   'h0000f ;
         Id6ff758a9c646a75ea986fe323b91966 =   'h0000f ;
         Iabbe6a5d643c1d8c3f7e2c8ddb41f8f2 =   'h0000f ;
         Id4b54da5ca05664d454c620a63622da2 =   'h0000f ;
         I0e4e792c6af3f2575e3e36eed213e7bb =   'h0000e ;
         I2c7afb36c88b388e24d0edf20acf3bf5 =   'h0000e ;
         Ibb053ae1486e202396d69ec80ceb37b5 =   'h0000e ;
         I88a88c8c4b3a9af4f49565aac9e5f248 =   'h0000e ;
         I359e996afe4b35d29d9180b990a27fcd =   'h0000e ;
         I899a8e3a18bc3f9e4f3a5af73fa61dcb =   'h0000d ;
         Ic124969a8cfb359b1ccc12c38b92f031 =   'h0000d ;
         Ibd06fe0881c395a5e679d87fb9ffdef4 =   'h0000d ;
         I8d0c94e6e41f653eeefb5b911e56e229 =   'h0000d ;
         I06d6e9bf2bf5fe1d0d06a7a7bf9aef4a =   'h0000d ;
         I3df5795d906a0f00bf42bf6e3ea2da66 =   'h0000c ;
         Idf0aba59612a66e3e74e0a90e1f24024 =   'h0000c ;
         I4ebe1cce938e487efd6289f437e5dc5a =   'h0000c ;
         Ia2818dffb7609ae601acc9bad920308c =   'h0000c ;
         I26a3e6a339b41ad00866844786681513 =   'h0000c ;
         I76b2e256804d1913c453dc19742869fb =   'h0000b ;
         I2ff4e3eb141f0d9f284bab6b5c9eb9bc =   'h0000b ;
         Ife7243ad867ecc4e311906fc4ede4451 =   'h0000b ;
         If65d250d229376f2091caa5d0eed8b8c =   'h0000b ;
         Iab0e973383f884115980f16a6261ebfb =   'h0000b ;
         I2c4e82e4c7fe3917596e9dfe8f01f865 =   'h0000b ;
         Ie17470e1d818de84c8e5e0269c5a18c3 =   'h0000a ;
         I25a3a01cc23b7303e828c5a76d108335 =   'h0000a ;
         I393c613e2dc208cf7724920ccf7da4a2 =   'h0000a ;
         I6dcc14bced84384b08b054ad1ed5d6ba =   'h0000a ;
         I93713849034deecf3189479b9012f123 =   'h0000a ;
         Ia20663615bcd8de7a403e368c23aa942 =   'h0000a ;
         I2623b7a7673b4061c0cfdd92e0119112 =   'h00009 ;
         I37517b2fa41b7fa2d25a45058b8369d1 =   'h00009 ;
         I613289d33f6a2742ef380880a6e4fe0b =   'h00009 ;
         I79d675be55634575c1ca36153e9b3637 =   'h00009 ;
         I5a21a18c1e1992154869c922fa691c74 =   'h00009 ;
         If8be80c27161a6257e0f1d41359727e0 =   'h00009 ;
         I7991f753713b02ebd49178ca1ca2f1cc =   'h00009 ;
         I040f9f3dc40e2bcc958191055ca6b6d2 =   'h00008 ;
         I70a8f1f9966c63b414a3bb68e5e3972c =   'h00008 ;
         Id8f36cdae93ca8a388aff8fb4806f4a3 =   'h00008 ;
         I906be6a8bc43d22dd04b47c2bba5c2f9 =   'h00008 ;
         Id4df0a1c44ea75f32970739cb4c5a2cc =   'h00008 ;
         I971cb87b4023114252557346c9a07d0e =   'h00008 ;
         I6e1912c5b6a09ff090f2d49d51002030 =   'h00008 ;
         Ia276ca65e85b9ccd4a9553b970b418a9 =   'h00008 ;
         Ia0b083b9bf3175a9961f79464d1b6bde =   'h00007 ;
         I6aea13b6ec3703c9c919731b7c43e44f =   'h00007 ;
         Ieb8b3cb38d28c4357bbd35d485f66dfe =   'h00007 ;
         I25fcdd6fea9bc9d728e5b6dc28cabee4 =   'h00007 ;
         I0ef97b8205f4a544cc31d1ab9fd62d90 =   'h00007 ;
         I157f4891b58262db67a57781e6789205 =   'h00007 ;
         I0306b43f29eb07e97472616ba7516f54 =   'h00007 ;
         Id8c72b2670ca8001c69b60551519f4b8 =   'h00007 ;
         If32e24d0be817c10df587ed0aac48af2 =   'h00007 ;
         I6c17cb40f5ab67595f89afc0aa3e570d =   'h00006 ;
         I2789fbaed627ab6bea83080a0634f73d =   'h00006 ;
         Id4415bf69046a95359a7f23a0ec3d5a3 =   'h00006 ;
         I25862ee3c8452b8f0d3187132477b77f =   'h00006 ;
         I5e8114931cbd9da66eec0a9e96b647b3 =   'h00006 ;
         I01a946c09a7ce0b62c7ba805e301de52 =   'h00006 ;
         Ice805f2d2607178baf73b8c8bdd1b725 =   'h00006 ;
         I77767e8e8a46c270774c64d18eebca4c =   'h00006 ;
         Iac7d03545a18a22c01e97d9f8ca93e40 =   'h00006 ;
         I1a60f16daa4667129838097d94c932b2 =   'h00006 ;
         I8f08550281859dc884c13197e046ef10 =   'h00006 ;
         I23978d82bd6e911f5366f97765be24aa =   'h00005 ;
         Ib26450dc355c3ca34ba704abe7350e2d =   'h00005 ;
         I29c302625d14d028e34ae65f37961e3a =   'h00005 ;
         Iede527989cec0a93d78423b7df14d707 =   'h00005 ;
         Ic0b1d8a6c00df4a35e285accfd1d149b =   'h00005 ;
         Ic82e6892a22a0fd064bdfbe31cc171f3 =   'h00005 ;
         Icd96d324832586b90e3d89709934fc9a =   'h00005 ;
         I07aea291890873ea17e211143a7a8291 =   'h00005 ;
         I424af84f8e7d7f4c85fe9e4632d0a5b1 =   'h00005 ;
         Ied903684ae1a9f6b1d39d3714b6db7d1 =   'h00005 ;
         I07e0123a7a61773a58a82d037140d1bc =   'h00005 ;
         Ideeabf83d0b70f18efb7a46d88efc352 =   'h00005 ;
         I148d4ff69853a123a3c5a306e978d9a2 =   'h00005 ;
         If578b689c5609b11df900bf92d0a388a =   'h00004 ;
         Ibc5a4c442eab539e5bb136a83112191f =   'h00004 ;
         Ia19a1d1736d5feb515750e680b83db4d =   'h00004 ;
         I98f9daa53631a03ce5f4d21fa499a734 =   'h00004 ;
         I3a1a9a79b0dd6856b5d6ef8eda18c564 =   'h00004 ;
         I9268175b692637227825c86f87dad083 =   'h00004 ;
         I1571e04768855319692febc19c86f630 =   'h00004 ;
         I382b613b4744799d708ecb0c361c7293 =   'h00004 ;
         I736ed9a09ea1b83b13fc3b53ded0c560 =   'h00004 ;
         I0e2430406a0c161380cfd60e7bbfa542 =   'h00004 ;
         Icfce7d26af22431c30d34d5738109a18 =   'h00004 ;
         I070f6f095b8a43ed92048d9fcd6625b2 =   'h00004 ;
         I7b5d1412081b2bad3b5dd0cffe78238f =   'h00004 ;
         I04e76b2c5bf274bc2d8b9862c3690980 =   'h00004 ;
         I7fdb420f639b22294c896a20c8036f02 =   'h00004 ;
         I7a40ef6e10e3406e1d8c57ae53c6c3a1 =   'h00004 ;
         I2e3fbfe6dd237424289f6f4d00ad486e =   'h00003 ;
         I2cef2ca61302b60079b80fd9f252c56c =   'h00003 ;
         Ib44222bf07803a788687a877f1491ef1 =   'h00003 ;
         Id5fbe2f0dbe2a2d864202212c5db88cc =   'h00003 ;
         I6f4cc724a3e77e3b282e08a162448b75 =   'h00003 ;
         I573fcd75e769729647bc1c5fc8e54852 =   'h00003 ;
         I806e05d43c46bf4f67ccf2f1afa2911e =   'h00003 ;
         Ia2f45ae7f344cf3de7a61fcc35ae4651 =   'h00003 ;
         I3debb601b68a3cd58ecdaa7d78e66c7f =   'h00003 ;
         I9bc3698d4111848c8ff7f5082b4e6f3f =   'h00003 ;
         I4f5449753716964b3600bbcbd44902f0 =   'h00003 ;
         I39de7cf13d732f3d5c89eaa718407a97 =   'h00003 ;
         I1936f1a842424a3fdc777207a05433c7 =   'h00003 ;
         I2b5d24b895e1386c5acec6ec51af70ee =   'h00003 ;
         I9cdec4376c54fd0d5892b20f7f3944e5 =   'h00003 ;
         Ic3dc6389680526e4e9f3db1a31c4e954 =   'h00003 ;
         I6de265c429ab7ef182f2ed2b52f413b3 =   'h00003 ;
         I17dd943cac50d93f041a310edf916616 =   'h00003 ;
         I2a2db61ae5f793391b0388d1139c1003 =   'h00003 ;
         I3a4a24d886c2c06e283081c1b0079aff =   'h00003 ;
         I1ae5bf5c035790ca6279076719f7d218 =   'h00003 ;
         Ic98fdc1a35fc3c698dd9c5bfe2fdd1ac =   'h00002 ;
         I0b771b927e8acb823e30239c89aafe9f =   'h00002 ;
         Ic3caaaecbbca186ebf9cc35e554ff62e =   'h00002 ;
         I33fc4ecd929152c59d62af65ecb38414 =   'h00002 ;
         I09a3008676f21e58545563dff1cc9328 =   'h00002 ;
         I566a0851428acd33e432b33fe3c42b4c =   'h00002 ;
         I96884d5c0babd2437ec14429856c0414 =   'h00002 ;
         I6a3539539860b98d7a310f63314a2932 =   'h00002 ;
         Ice31c844af4b8c3b966b778cca601527 =   'h00002 ;
         I8eec3d66ef763226b960a24192aafe27 =   'h00002 ;
         I093a0ecd0a1aaea8a97d08d54cd37fec =   'h00002 ;
         I3b2708fccba619958a392242efbbeea7 =   'h00002 ;
         I543deb703bb9eb808f4381f543e408de =   'h00002 ;
         I0e0c7e753509c664971fd12be9183537 =   'h00002 ;
         I68577e7dec24946ec0745c5d4255795f =   'h00002 ;
         If53e38b5b6031a7e927a65f90acf5120 =   'h00002 ;
         I372a38a8675f65c5257b645fb5d809af =   'h00002 ;
         I0d37309bb37b707e10a4e12425157fe3 =   'h00002 ;
         I5935a4ee604a8c6259d88bd4b679babf =   'h00002 ;
         If4ed201fbbaa5ce9bfd05d65d79458d0 =   'h00002 ;
         I9b11c7aa2d35ee4589dec055ab0df2ca =   'h00002 ;
         I45a6d3691aef6c693ae6ee25c25a4b24 =   'h00002 ;
         Ia15364dea1e0f0243204b4bc4c9b8bb9 =   'h00002 ;
         I2f31acde416c079c48ce54697eac5e60 =   'h00002 ;
         Idab577631403b170aa07d02c7d455315 =   'h00002 ;
         I36b79e4befc1673140076d2f9cbc9d82 =   'h00002 ;
         I9f263275a24efe9297aa995282c48360 =   'h00002 ;
         I7915e8a9a775ea1bc1bf7fe71648303d =   'h00002 ;
         I4a7ac8c9709967341ededa935aa65581 =   'h00002 ;
         Ibd7437a655d4985728ce070004e3b419 =   'h00002 ;
         I8a834fd9d1425a79f7ff0713777fcdcc =   'h00002 ;
         Ia60cc135f03b89516e61d52335e69674 =   'h00002 ;
         Ia1b1f012b02265afed03cb146e88f2a0 =   'h00002 ;
         I6095ee8675c10be082abccd7cef7ceeb =   'h00001 ;
         I2be07fc5652209f0e8eda31090dbb162 =   'h00001 ;
         Ic60fc4bb6e7ccb8bee260e5b982bc5a1 =   'h00001 ;
         I217d1876f768c7dd3eed096e2de59dfd =   'h00001 ;
         Ibb297f22ba2e0d4786042f7503ff3f61 =   'h00001 ;
         I8d917a51d32729f4a5a98b5d3a40f947 =   'h00001 ;
         I08213a1a86aa27e3d3ed2d294d972ea7 =   'h00001 ;
         I271dfdeef4359fa9b2ebf80ca950a08e =   'h00001 ;
         Iff44a32b2e9a1a65d820b0839313015e =   'h00001 ;
         I2882587956babd713eb3a53af6afe389 =   'h00001 ;
         I4f1ca888cae3ee3efeefafcfb12e16b3 =   'h00001 ;
         Icff2aa823d2f0e9421f3fbce6d21f510 =   'h00001 ;
         I2cd19bf0afc4563ea24619849ab7d8b7 =   'h00001 ;
         I80cae65874911e05bc77db3e5fe0fcd2 =   'h00001 ;
         I18c43491892bd258dfd07aa0263c5479 =   'h00001 ;
         If322bf2a59be9bf7b33a49a6baf72ed7 =   'h00001 ;
         I2bb21cbf03db27c0b9d814517033b56e =   'h00001 ;
         Ib408b39624c6576c228f32eed26ccf8b =   'h00001 ;
         Ib6dee36145f77a6f1364c218140266b4 =   'h00001 ;
         Iafa25738d96fb115c78d8d295902c263 =   'h00001 ;
         Ie7cb395e7ce65ca399d99a5e62a7efad =   'h00001 ;
         I1bee0c6e3a24ee319d219799ce58f13e =   'h00001 ;
         I7fcbf3d532ed0c810cdc1c5be536d263 =   'h00001 ;
         Ied7f9cbbcacc43332f1219e8bd0a07bb =   'h00001 ;
         I491888fefe23bb0bef60f293668491af =   'h00001 ;
         I1b9368c7a0d236ed73a6783281144bca =   'h00001 ;
         I2adf1f34eb55f6f7e5f37b328b2bcf21 =   'h00001 ;
         Iaa61cf5ca911de351708963438768cee =   'h00001 ;
         Iacba64081faa56ef9190aa65fc89ae7f =   'h00001 ;
         I5d41596aeb3aeb4f07dbc0c995b5f4a3 =   'h00001 ;
         I1c01c903faacd546e44a6fd6564ef3bd =   'h00001 ;
         I3e3195b93f03e3c8c24655259f745374 =   'h00001 ;
         Ie229e972daab0a41969c5cc066e52e61 =   'h00001 ;
         I5a646f85f9e6d52063b0c0e6f479f6f1 =   'h00001 ;
         I01a50cb46ae1b229eda9094867090aae =   'h00001 ;
         I68026b1eb748133551563bea029c3488 =   'h00001 ;
         I726047b0a4d45f8ad1f394301dbfb78d =   'h00001 ;
         I2cddfa0b89e0aececac2dd7d983beb26 =   'h00001 ;
         Ic5e1dd806582ee08eb6d1048d6617b13 =   'h00001 ;
         I9040f68430c75ce7527990dd702b7feb =   'h00001 ;
         I40ebb4eb571f18c2fb810daab0d5770f =   'h00001 ;
         Ia4738ee511867aa46e0e92f3d86c4ccf =   'h00001 ;
         Ic10326eae7434399af6e611e31389963 =   'h00001 ;
         I8fafe7fe582d027b97dbf2cc58763096 =   'h00001 ;
         I8a329168f83731c15dbedb1f1f966d78 =   'h00001 ;
         I603a5f82891f62b59f7890d631d0b6df =   'h00001 ;
         I620517db078658289fcde4200f15ac06 =   'h00001 ;
         I51271c02c6fd9cbda153c9b28aa099e3 =   'h00001 ;
         I8def31183d1a648a6a50245eeb6b57a1 =   'h00001 ;
         I0c3a1185a9fbb05c0dcec0d655068786 =   'h00001 ;
         Icf0284aeb5d603e893733d2139a79ef3 =   'h00001 ;
         I3d0e6fa7f7edbd105fd8f7823722bcf0 =   'h00001 ;
         I55e28dff0ebd1007f4f00c512f1df1b7 =   'h00001 ;
         I2b33fef3c83dab2f2d254cb295264482 =   'h00001 ;
         I1689bfa3340ff4798ef7eb160714ede5 =   'h00001 ;
         I1b5deee5754dcc0762ca2691fd927056 =   'h00001 ;
         I1e63fce77120b91dc6195d2febce4d42 =   'h00001 ;
         I1d3f5624cb6f217fac422833ed8b7195 =   'h00001 ;
         I1fde6652c1fb298d84e88620edc9e91a =   'h00001 ;
         Iffd2d0fd17d604ddadcfc2dd9e46276a =   'h00001 ;
         I8295b6fa92e241d4b689ad0e26f6a2db =   'h00001 ;
         I8573b3db0d36442c2f233d12586d82f5 =   'h00001 ;
         I5319144e65be1e69c9ef767bfecd4ea3 =   'h00001 ;
         Ie7da9e9fdd626504cb2f00a3ec899718 =   'h00001 ;
         I8293d7dc145b31d28c05c02677760e9a =   'h00001 ;
         Ia372f6e388ed5cf8e9810c52d3749136 =   'h00001 ;
         Ibd959e3bf9ef7ee76ec2754a06926d9a =   'h00001 ;
         I8f03815159c11486a4805e7f72c84a38 =   'h00001 ;
         I15e5e06b7dcf6616094faeb798a0fdc8 =   'h00001 ;
         If23f4bc5d45a3e7a22a9e8596b99c575 =   'h00001 ;
         I70afe2bb83173aa96269271270d03f2e =   'h00000 ;
