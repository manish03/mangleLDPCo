reg [flogtanh_WDTH -1:0] I0c1c52a843a5de4bb5e0eb6897ea37c4,  I371284eed470112cb89e1d361a9d40f7;
reg [flogtanh_WDTH -1:0] Ice4c8b10e41f361db2bd4a7b8470b05e,  If0fb2e90431d89d99912918f83036f4c;
reg [flogtanh_WDTH -1:0] I612d62c35e606e6e91220910fd8448f1,  I0ee915f21334d38c75f0207e3b052a69;
reg [flogtanh_WDTH -1:0] I4f664d460f924a71ebd3cc05f0916521,  Icf5a9bd712d310ac17eb2354f884a237;
reg [flogtanh_WDTH -1:0] I0e38bd43118f53204e169f324066b75c,  I3222cf2f98878be3f453560ddb3dc43c;
reg [flogtanh_WDTH -1:0] I46878ad6c93d318bf7a959c78090bf66,  I2dd9e89f2842e748c1574ad0e7f4dba9;
reg [flogtanh_WDTH -1:0] Ie2c597c226457d94ec76f1513d95aab2,  I667adc16c92bec8f413a1a9bbfc41ce5;
reg [flogtanh_WDTH -1:0] I2c72e48d1e2274c662c18b729af96161,  Ie6aa50a44574542826b78fed7d77b76f;
reg [flogtanh_WDTH -1:0] Id416e2e4f204401c79d97ae6ae1414ae,  Ie97072fa52f483bbd89f019c21152cdf;
reg [flogtanh_WDTH -1:0] I8fa96c5580fd6050e2a8c5fcb77c9927,  I47f153e1cecaa77f1e6e6f07c0220557;
reg [flogtanh_WDTH -1:0] Ia9569f758e6bc743aae3a2bb51d941ee,  I1b9dcfaf144b48a64b990e5b020d4a02;
reg [flogtanh_WDTH -1:0] I00ae3aaf6b44b2f7fd9bbceafb9c4e22,  Ie32d4bd927d02e547850331db8028177;
reg [flogtanh_WDTH -1:0] Ibfea7f98ec3bbe5588eb75cbcef739d7,  I0988db7ca497541e372131a0b0e8075e;
reg [flogtanh_WDTH -1:0] Id9eff948ed9da8502308740b4ae17dbf,  Id13b5577b8baa586fedd34d4aab9d9c5;
reg [flogtanh_WDTH -1:0] If9d08c27c57ed8293171486ad65ed95c,  Iedd0e0f6ee682a131d4f14c4762ea0eb;
reg [flogtanh_WDTH -1:0] Iace1409bfc12437ef093b91d50c8175a,  I875d7c55914414298f0fbec0b345c92e;
reg [flogtanh_WDTH -1:0] I506d9cf5c368c130a8517f994e7f7a43,  Ide64c9647c7898867e0d036e9ff95f6e;
reg [flogtanh_WDTH -1:0] I0f3fb929c6ee46d33daeba7024107aff,  Ied6ccabb348ed7e20567011e027c86ad;
reg [flogtanh_WDTH -1:0] Id3ac7026a6f63b1dc8588f9bdfd50068,  Id030b072054c623c7aac5c571d052951;
reg [flogtanh_WDTH -1:0] I680caae24965f4516cbd8642d4d43b3b,  Ice55fb2e506accf518b4aa18298d017e;
reg [flogtanh_WDTH -1:0] I7b240e087870bef3e01b2de04cdbae13,  I07a0167dcdfc76612e1b0da251337a7b;
reg [flogtanh_WDTH -1:0] Ic2b7c4749006adaa1dfa0ca1c5d7a371,  I045e08f48738d395af2b79f25af73732;
reg [flogtanh_WDTH -1:0] I2abc1d3ddcecbdbdc971abb93be58744,  I7df57f27a880fe45f78c108f8faba963;
reg [flogtanh_WDTH -1:0] I9fcc49fa3eb8ad62633822ff3ac5973a,  I60204c1d3a96524bbbdf715f95f08fe4;
reg [flogtanh_WDTH -1:0] I6b938059b8a71491bf1718326233b688,  Id5b9ae91dc900060caffff2520236f66;
reg [flogtanh_WDTH -1:0] I5d98a20b0eef6a335b29f017cd3120df,  I861fe9da6d004ce3998ab54a8c0d62af;
reg [flogtanh_WDTH -1:0] I69d5314c6ba43f6d015acf00c8a2a7be,  I95caae0432aeadc0cbe279f9d6f9062b;
reg [flogtanh_WDTH -1:0] I64ce8a8f7f046222c963820f37362021,  Ic9c3b015d5830bf4834a435eba89caa5;
reg [flogtanh_WDTH -1:0] I4e1c98665268d59e19c3068ff9efe9a8,  I6e18dd1a579e09b80ac113fe85b483b4;
reg [flogtanh_WDTH -1:0] I1399a46a42c2cc384efc8ca681b1b249,  I51c1c8e8df14396c5c77b5013531a84f;
reg [flogtanh_WDTH -1:0] I3e0d577c49e0fcba84112e3afab2edbe,  Ie8f75e8e020d43f6a357b5175047c254;
reg [flogtanh_WDTH -1:0] Ic266aa3f20103455635f801a0fe1056a,  Ie762d8aa151448cbaa0d005a3c01572a;
reg [flogtanh_WDTH -1:0] I285c0d0dbcb505b98bbf005805067396,  I293b32c043e20d6baab178319dd1e2f6;
reg [flogtanh_WDTH -1:0] Icba253e44f98c391c02e864856715f49,  I200aae813b664e02075eeefbc3b4450d;
reg [flogtanh_WDTH -1:0] Iaa4b6b01007d9836ae0092101c4065db,  I006264bde45d8df078ef711c221ff387;
reg [flogtanh_WDTH -1:0] Ia2f4d61e666ea4e0d8085325cdaa7344,  I9200a0071528b14dc52e92082768ca97;
reg [flogtanh_WDTH -1:0] I84ed644f3578e53744802bab05d17011,  I55761decd7043b4dc82737b9d6ef6e7d;
reg [flogtanh_WDTH -1:0] I5fbdad2d56ab8f5435a712b512190645,  I4f51d114002bdfd69a31f95c2fa5234c;
reg [flogtanh_WDTH -1:0] I670a7cf3b4948b0d31c871ba641af4c1,  I796cb71b28957405c10015a2ab7124c6;
reg [flogtanh_WDTH -1:0] I227702af9307eb6600ed78a648bb71e9,  Ic85bacce5db48b4dd3f626749f6effa8;
reg [flogtanh_WDTH -1:0] If0c4078bb97b3a246a91be4180ee7af9,  I2a508066cf0e07bbe8a91f276fbb3078;
reg [flogtanh_WDTH -1:0] I913f1af34aaf3d51d3c60489979a81d5,  I85913ae95fcd63de45030d583846b1d6;
reg [flogtanh_WDTH -1:0] I22e712371781d71cbb80680359ccd708,  I971cff06a60916ea3e136b397d4c620b;
reg [flogtanh_WDTH -1:0] I5e9450b27761da0b895a4f6ace1ad171,  I2c363f7abf62c9026d0b0dfe5a51207a;
reg [flogtanh_WDTH -1:0] I0b1bc20ea62f64bae807d8ac1166139f,  Ia5043b0c8ee086c66e683eb115a75484;
reg [flogtanh_WDTH -1:0] Idddfbcad405258a5434d8b94eb26654c,  I6b7b63ea23c5b4f3c597f121284cd2da;
reg [flogtanh_WDTH -1:0] I8beef0ea5356b2f46d7d5f16db49ebef,  I3cf82abadcee2faa1849d0a9a45b051e;
reg [flogtanh_WDTH -1:0] I499586880161ca66628afed78e7e495d,  I8b42f5455dd8f6323d7a4e28c0eaa1a9;
reg [flogtanh_WDTH -1:0] Ie909ad4a9ba2fde8fd6451e7eda2088d,  I608597017b046d92b77226999df90600;
reg [flogtanh_WDTH -1:0] Iee75fb439b2200aba94b03fd69cd7adc,  Ia39b908f8d6b63777376ca560cd0cc8d;
reg [flogtanh_WDTH -1:0] Id8a8555f4bf9003a0ac0dcafaa67e68d,  I87ad38ab473927df7c0bd69c6b4b4c5e;
reg [flogtanh_WDTH -1:0] I10065fe206e6700159260af61afa61c2,  I8e70752f74ecdbe95a7b33ca264d4589;
reg [flogtanh_WDTH -1:0] Ia41593b7790fde4ae4dd986dd583286f,  I6e768e27a3f1804919e3f83c050e19ba;
reg [flogtanh_WDTH -1:0] I44490a711aece8f1a24c080cd0f37607,  I2285f424ef2b8b2041267c1652155ad0;
reg [flogtanh_WDTH -1:0] Ic35377a5686c5a6edace93b58129cbdd,  Ibc5b97632aab1e763ac51f8d18edc792;
reg [flogtanh_WDTH -1:0] Iccd1e1793be28ddad794782e2700a4d0,  Ic4a0165bd71d9e586fdc66c824e45224;
reg [flogtanh_WDTH -1:0] Id112833f079dcf6e092d48cd13120d47,  I40de7aeac837276e7b3f0c4b29ce5eca;
reg [flogtanh_WDTH -1:0] Ia550c5040df02dc8a8735562e71ddf6f,  I024a746142e5ff074724f92af62f3bd3;
reg [flogtanh_WDTH -1:0] Ibcaed8bfefd254ded778d760cd533b81,  I1e54f934fa92e681472d03199991f0b2;
reg [flogtanh_WDTH -1:0] I19c7906957daf8e2a04b013e95db9c6e,  I8cabd17b81e99a86fc8704aaaae629a3;
reg [flogtanh_WDTH -1:0] I4bbddbcd811dc6936fd20d18559e3aac,  I54c1bf986182c83540d950762048a5e3;
reg [flogtanh_WDTH -1:0] Idaf09a27ce68e8877da2d4c48be4c8ca,  Ia5fbeb5be349b8088a749e25a9e6e416;
reg [flogtanh_WDTH -1:0] I82ad270d36061ef06232de9b92742dfd,  I987b220a4729d14e9fc97b57867436e4;
reg [flogtanh_WDTH -1:0] Ieb5d1ef84057ceba02d9db624be39285,  I7f1d9309d3053256134130574b970425;
reg [flogtanh_WDTH -1:0] I7ebd34e6a95c3589b44cc0941f54bfa9,  I9fd9d5a2a3a34b532bad740b16ce66fb;
reg [flogtanh_WDTH -1:0] I46432f8bb8f39efef70554ea0e8573de,  I66a648a9f6b10b1d580e72b36a1ed9e7;
reg [flogtanh_WDTH -1:0] I1fb7b6a528ec8d5871cb15a490bbfda2,  Ia08c041d1aacfbbd1f8d7980923b9b05;
reg [flogtanh_WDTH -1:0] I25d429f4a9f397a0d0ca515241b3c1b5,  I6805a2f26b1e51f7ac0087e6829b3c5c;
reg [flogtanh_WDTH -1:0] I3ca008900582aea13c5cf09b6c3af78e,  Icc11f9d183454b33624bd411710342a0;
reg [flogtanh_WDTH -1:0] Id9a5e1c4a044b3006d620dd52e2e8ddc,  I18f145bedd3864fcebd983f9533a5877;
reg [flogtanh_WDTH -1:0] I63f34eddeedc5ded8721b40546c758c3,  Ifa25d4c9ccc3efd1af4e711d3c32e9c5;
reg [flogtanh_WDTH -1:0] I8ec5f00523507f51358081e52a5bc55c,  I5bbf8f01c5ddaa02516dde3867ec3d78;
reg [flogtanh_WDTH -1:0] Ib77465ae19c99c6e2c39e2ab6438730d,  I3f8fe2d052a6df20dfaac6f88d4fff8a;
reg [flogtanh_WDTH -1:0] I025a54040366d4505896c1179d580dc1,  I9fbf9bcb6022bb550bc2dbd52f20d05f;
reg [flogtanh_WDTH -1:0] I0ac7e4f7f0e68450455e4a3d3ed57c56,  Iacd71ce5854c85450463a0a45ebc6a2d;
reg [flogtanh_WDTH -1:0] If6f5c61447dbeeaef688c670c9802649,  Id7c1a8f42cc90b7846105cd103b07228;
reg [flogtanh_WDTH -1:0] I968168f5cd481033283f24425f7862b9,  Ic6d94b59cd6f4c7765463694c9fbae3c;
reg [flogtanh_WDTH -1:0] Ie364b2799febe180ea9c2361279bcdc3,  I11a9409c814372a31d771888692ae955;
reg [flogtanh_WDTH -1:0] I76cc2a7d1f750a49780fe7e7f1651d5e,  I760f9ff7bc594c98e71080485cc1a082;
reg [flogtanh_WDTH -1:0] I2e3ac4cb975151fcb26d716ef80a24f9,  Idb9be12ba6807752b0c36f4cc18843cb;
reg [flogtanh_WDTH -1:0] I6da8878ff3f8680907597ba4ab49e7e4,  I192119ad6ad1396dd6fd1fab6e4c4cca;
reg [flogtanh_WDTH -1:0] I28db3b4aa4f26a48ef6a28956536d15a,  Ib4c62a865f79eaa2aa5fbd12860f2e80;
reg [flogtanh_WDTH -1:0] I7b95e7f8f8f6d01ad095fdfbe36e7f6d,  I5fb195f29a4e02620d2cca6e7f2a8fa0;
reg [flogtanh_WDTH -1:0] Ieb56b02269e16c20b5f626afc1b97c98,  I41b4d1d3d5ae22c8fe4f1e0fe20ccac7;
reg [flogtanh_WDTH -1:0] I486565b0e63446c0b122a62bac6644da,  Ib2afa3be272607c236cbd5410a88e8c2;
reg [flogtanh_WDTH -1:0] Ibd4082b5df0c5bca554397e77fbf589e,  I43587e6827dc7dc1ef38d552f6a73ca4;
reg [flogtanh_WDTH -1:0] I6361b4f6c6266288a5f53dfbf0e514cc,  Ic27ed0f98cad254a72ade8253ccc01d2;
reg [flogtanh_WDTH -1:0] I0590fa4c4cb5194e038b57fd416210b9,  I5860a511728dad8112a9246843f0fdab;
reg [flogtanh_WDTH -1:0] If8409ca3930cc882752b4efe399aa107,  I6f83f4d8681a17b7e700a38a78917822;
reg [flogtanh_WDTH -1:0] I509f64436f6d698c58fa255372adf7e7,  Ic902ce884c81efed3160715af43eb19b;
reg [flogtanh_WDTH -1:0] Ib6319f6f8e74409bd60d624b07fc75d2,  I8297012f23a474aa863c56e6ab9f77f4;
reg [flogtanh_WDTH -1:0] I344f88b13d6f536724dd33ed2d9fa07a,  I703fa28fdfb32f8e7fe5062a3332ff6a;
reg [flogtanh_WDTH -1:0] Ia9c1251bf7d48ef32d67ee176ca55e07,  I4d60a4630a93dbf6460fc525f16fb69b;
reg [flogtanh_WDTH -1:0] I8a885ced1613614d0bc3e1d2ce31cd34,  If6a1f518420fbc246e2524469689a5e7;
reg [flogtanh_WDTH -1:0] I084e8923b177a76c4fbed301ae5f905f,  I48c55cdc6c1e3bb5e36a5451cb43c5a9;
reg [flogtanh_WDTH -1:0] I58d2c7aa1ec77bc041b6b1e2e4ad8277,  I147accfb14f15341869779b74c8cadb6;
reg [flogtanh_WDTH -1:0] I9be477a653c8d0bd98ea404fa8876dd5,  I0d302535ee6928ed74d7b456efaf01e6;
reg [flogtanh_WDTH -1:0] Ifefb2b21271a5578ec1e1d9ddae2047c,  I0039a78cbf75de3d875c319e3bc08d22;
reg [flogtanh_WDTH -1:0] I708bb50785dd2710e712438dcfec5eb1,  I7a43154a62ef625844cda08b1dfc9c79;
reg [flogtanh_WDTH -1:0] I12e20bdca30dd5a4695333353faaafe1,  I8e05a477fab7c0c6f70c681626640b93;
reg [flogtanh_WDTH -1:0] I37da1f9f97e273359be9e4912f8a8ee7,  I51393ac63dc5f8c0898ffa6dd59ee183;
reg [flogtanh_WDTH -1:0] I0df8e26f5e3a60744a02e8b50cff23a5,  Ib4f7dd6e43c7a291d753f96b1aac8ce6;
reg [flogtanh_WDTH -1:0] I0f005326cad2001188a9fc4b919bd19a,  Ibf76adf5511e851727200f4fd60bf34b;
reg [flogtanh_WDTH -1:0] I1b7f0cb10a2a1c63083aa2e5d5fe84d8,  Id90de24703e5b15356a8ab3862612957;
reg [flogtanh_WDTH -1:0] I43240748b90a2f1b2738d7773256f36c,  I2b42badcbe3d18d033edbd6d4663fac6;
reg [flogtanh_WDTH -1:0] I9d301fb4da56021d4bf0df8dd2719eb4,  I72450aa2c2f2f501a5465f008e95ba4f;
reg [flogtanh_WDTH -1:0] I50188fbeeabb5bbc1549229769cc58d3,  Ib802f2c9c1265a47e5acfc419034488d;
reg [flogtanh_WDTH -1:0] I85af941bfb4adc588579de64e51887bb,  Idb28449172f54add7ac6fd1287543a5b;
reg [flogtanh_WDTH -1:0] I6baa38fdfb9b81d807b09ca3b7cd5d32,  I6b33174bb2786da0ba9ba988a96aa5bf;
reg [flogtanh_WDTH -1:0] Ica83cfc4696601a6936e577389a395cc,  Ib68892cce1de9f46fb391a7ee8a01afb;
reg [flogtanh_WDTH -1:0] I9ae9897faacb46733dcec0b985a590ce,  Ia0e39ef7db11ff2f95f50e6a912e945e;
reg [flogtanh_WDTH -1:0] Ibcf6f538d26631634b6ceafdd3ee991f,  I1f3153881fc6a7fc767a33253f80e06f;
reg [flogtanh_WDTH -1:0] Ia2d7c7007306e7b2ca65518fcc005588,  I994e4d13d16c12025cb60205b8f7559f;
reg [flogtanh_WDTH -1:0] I5db8abcf5c9f55ffbe360502c0acf592,  I3e4b2dbb8f44350c5cff7430502401b7;
reg [flogtanh_WDTH -1:0] Iebf161a4f32971bd911356670349e894,  Id1e6e9ac8ddad3aedd347aee9f615d9f;
reg [flogtanh_WDTH -1:0] Iba78cb5ab1da071088bf8f924095d1dd,  I5a6da3732e0f265ad95269f5a629c1e8;
reg [flogtanh_WDTH -1:0] Ib8bc0d119e76d93a801d9749ff205d30,  If8773fa380ec5c1199794d4128d443f1;
reg [flogtanh_WDTH -1:0] I7d760437e7830701c90db6653febff5a,  I63283e5286a737d3ba1f99ae29902bb9;
reg [flogtanh_WDTH -1:0] Ie7d3e4264ef52d194bcd054dc421e97e,  Iedcc3a589dba858f1193b1be582db24b;
reg [flogtanh_WDTH -1:0] I2271582af0c776dadff851456aa6e4a7,  I8a87d3adcb2989738d70db84c3b97a3a;
reg [flogtanh_WDTH -1:0] I851e3c75bf75803e1d745053721aa9ad,  I267e058f7db05744d80df6b52be83475;
reg [flogtanh_WDTH -1:0] Ifa32facd628d97fa55482c63464bbeed,  I5e121581d8a5f81fc84da2fa982d8fd6;
reg [flogtanh_WDTH -1:0] I37a83fa1dac26d4614760db718790dfb,  I51f875fbf103d8b8093d73279f127843;
reg [flogtanh_WDTH -1:0] Icdfa771d45c36fef80efda13b0481130,  Ifcbf9c1d4d6f111f06212e58764d29ea;
reg [flogtanh_WDTH -1:0] Ic72a44c59c204b5d5b77523429df133b,  Ie0e816b57f511fc0479210deebbd9fc1;
reg [flogtanh_WDTH -1:0] I1395b926b6d89fdfe41444e3a94d0d10,  Ia7673dc1d477d486371935040ff7dce9;
reg [flogtanh_WDTH -1:0] I8393828bf7f4ce64ef97785fcd0d65fb,  I7df5c4ad52bf35d254a4a14771a28fe7;
reg [flogtanh_WDTH -1:0] I2f6dc9f6f5d1316b9426bbe277b82427,  I9ae2d00bf699c7f12c3f5d78ad2c405c;
reg [flogtanh_WDTH -1:0] I60098787140a26167a69e135e08c6e8b,  Icb740a93e2adc0a9f18ac25d0c5d018c;
reg [flogtanh_WDTH -1:0] Ice5b808b49ac5331f4fd6f36e74f0897,  Ia9691e7c587528f3ca0d85d842225da4;
reg [flogtanh_WDTH -1:0] I3480a29289d8eca6cbf762b798ec68fc,  Iab732884bb2d4b1781e31c7a1c109000;
reg [flogtanh_WDTH -1:0] Ie8718369d950a31dd1e9b307ce68984c,  I67d8e4c822cc57b150a76dbb3478b5b5;
reg [flogtanh_WDTH -1:0] I954ad53f646754aa0c8db5073aff65fe,  I3bb2f03bf7d2f7480187062b45c6fdd9;
reg [flogtanh_WDTH -1:0] I8f9194a8b73a5008a74dfe09429e455b,  I8e57236f80078ae72706aa8102e1bf53;
reg [flogtanh_WDTH -1:0] I9b0851ae1b88864bd086003066137b86,  I1732bcc59b7bad3d08b232d099fdefdc;
reg [flogtanh_WDTH -1:0] Ia8d552e62e3c642796936c2c4188f8a4,  I4b568309171ac557250c2ec600b9d7b0;
reg [flogtanh_WDTH -1:0] Idaffd115023b38f3f7e7cafe8e2cedb8,  I886251a3307e5fe20788c8e947f4ef37;
reg [flogtanh_WDTH -1:0] Id6ff758a9c646a75ea986fe323b91966,  Ic0d064e8436ad001f7e9d97e800e5636;
reg [flogtanh_WDTH -1:0] Iabbe6a5d643c1d8c3f7e2c8ddb41f8f2,  I9f2ba5b0600c5eb81cef40d0822d0aea;
reg [flogtanh_WDTH -1:0] Id4b54da5ca05664d454c620a63622da2,  I2aaf6ff0daa3d3e26b197e6895cabf3c;
reg [flogtanh_WDTH -1:0] I0e4e792c6af3f2575e3e36eed213e7bb,  I2e8c68a51f1f1f4e413897791a6823a0;
reg [flogtanh_WDTH -1:0] I2c7afb36c88b388e24d0edf20acf3bf5,  I1a318a04ba3cf92f4ba0dc132a564040;
reg [flogtanh_WDTH -1:0] Ibb053ae1486e202396d69ec80ceb37b5,  Id32b88b33bfbcf79ff0a10d447f69619;
reg [flogtanh_WDTH -1:0] I88a88c8c4b3a9af4f49565aac9e5f248,  Ia41215dbdcd4b27a8ab41f48d40d644a;
reg [flogtanh_WDTH -1:0] I359e996afe4b35d29d9180b990a27fcd,  I53c239961c5745db892194a0a62b5d57;
reg [flogtanh_WDTH -1:0] I899a8e3a18bc3f9e4f3a5af73fa61dcb,  I0ffed4dfc4e97bb477647e5eab3a18f3;
reg [flogtanh_WDTH -1:0] Ic124969a8cfb359b1ccc12c38b92f031,  I46fcaa5311cc831199bb4a5a3dba797e;
reg [flogtanh_WDTH -1:0] Ibd06fe0881c395a5e679d87fb9ffdef4,  I69b693e03eccfe9a889894988c0c9a53;
reg [flogtanh_WDTH -1:0] I8d0c94e6e41f653eeefb5b911e56e229,  Id0ca109680ce0cb6603139baeebac59f;
reg [flogtanh_WDTH -1:0] I06d6e9bf2bf5fe1d0d06a7a7bf9aef4a,  I7bcf3409fb1f7bf880f945db8f2eb6c2;
reg [flogtanh_WDTH -1:0] I3df5795d906a0f00bf42bf6e3ea2da66,  I873254d95f4a9976acf9210228365521;
reg [flogtanh_WDTH -1:0] Idf0aba59612a66e3e74e0a90e1f24024,  I2a437c10a562e8e7f4cef30bbfde2fd3;
reg [flogtanh_WDTH -1:0] I4ebe1cce938e487efd6289f437e5dc5a,  I50e26d2184d04613f297357308e7c91e;
reg [flogtanh_WDTH -1:0] Ia2818dffb7609ae601acc9bad920308c,  I8b14ff6b303ae081ae414ca7a00da3eb;
reg [flogtanh_WDTH -1:0] I26a3e6a339b41ad00866844786681513,  Ibf3a99967d7cbab53676fed78da28eb8;
reg [flogtanh_WDTH -1:0] I76b2e256804d1913c453dc19742869fb,  Ifb6cf60f578b5a5dd0c27da72408cbce;
reg [flogtanh_WDTH -1:0] I2ff4e3eb141f0d9f284bab6b5c9eb9bc,  I000bdba9ccdb068a02fd37d2991675b6;
reg [flogtanh_WDTH -1:0] Ife7243ad867ecc4e311906fc4ede4451,  I5110f5370812f6d0319c0f42a6638b5b;
reg [flogtanh_WDTH -1:0] If65d250d229376f2091caa5d0eed8b8c,  Ic36cb86884806afb677ac8fb42aead36;
reg [flogtanh_WDTH -1:0] Iab0e973383f884115980f16a6261ebfb,  Ie4dba51278ebf8a9358c2019383fbaf8;
reg [flogtanh_WDTH -1:0] I2c4e82e4c7fe3917596e9dfe8f01f865,  I96373fc8bdf40551ef8206b4ba38cd98;
reg [flogtanh_WDTH -1:0] Ie17470e1d818de84c8e5e0269c5a18c3,  I7b8a50810f6a4c27a23c82330707c4b6;
reg [flogtanh_WDTH -1:0] I25a3a01cc23b7303e828c5a76d108335,  Id84a4cc9f82244c2357edc537824eb30;
reg [flogtanh_WDTH -1:0] I393c613e2dc208cf7724920ccf7da4a2,  I8866b1e80ead799943d3ad273ee0c97e;
reg [flogtanh_WDTH -1:0] I6dcc14bced84384b08b054ad1ed5d6ba,  I33d92c1bdacf71fa60865f1741288cdf;
reg [flogtanh_WDTH -1:0] I93713849034deecf3189479b9012f123,  I834a4a93056d8777cd2d4996ae33122a;
reg [flogtanh_WDTH -1:0] Ia20663615bcd8de7a403e368c23aa942,  I51bc583f480542f3f95241643bb39eee;
reg [flogtanh_WDTH -1:0] I2623b7a7673b4061c0cfdd92e0119112,  I35539407bedb7d43642e952787216ce6;
reg [flogtanh_WDTH -1:0] I37517b2fa41b7fa2d25a45058b8369d1,  Ifa78beaa6ae7a7a32f4886a14e4d1532;
reg [flogtanh_WDTH -1:0] I613289d33f6a2742ef380880a6e4fe0b,  Iae691c305b2fd52617ef92705568a8b8;
reg [flogtanh_WDTH -1:0] I79d675be55634575c1ca36153e9b3637,  Ie87c6bd3452b53ef57df5f420f351434;
reg [flogtanh_WDTH -1:0] I5a21a18c1e1992154869c922fa691c74,  I03106ddaebe00bc59e1611573835f727;
reg [flogtanh_WDTH -1:0] If8be80c27161a6257e0f1d41359727e0,  I8b947b6c3139066fbd5873d5b818183e;
reg [flogtanh_WDTH -1:0] I7991f753713b02ebd49178ca1ca2f1cc,  Ibb1c668cb8ad3eb49b9bff842d118aa7;
reg [flogtanh_WDTH -1:0] I040f9f3dc40e2bcc958191055ca6b6d2,  I4c3bda40c1fe5dbacee1829e0d60bcab;
reg [flogtanh_WDTH -1:0] I70a8f1f9966c63b414a3bb68e5e3972c,  I405504d762cd698722b183721df7243f;
reg [flogtanh_WDTH -1:0] Id8f36cdae93ca8a388aff8fb4806f4a3,  Iae9c6245aa98b5758df6d57f8c33ab31;
reg [flogtanh_WDTH -1:0] I906be6a8bc43d22dd04b47c2bba5c2f9,  I35f897e994d6fb9ae452bee5b423c4e9;
reg [flogtanh_WDTH -1:0] Id4df0a1c44ea75f32970739cb4c5a2cc,  I413a7fe2255064627ed283d35d910de4;
reg [flogtanh_WDTH -1:0] I971cb87b4023114252557346c9a07d0e,  Ic930f61e087bf2477712e8fef9c413d3;
reg [flogtanh_WDTH -1:0] I6e1912c5b6a09ff090f2d49d51002030,  I61ce1d41fa5221c01f7e9571965eb3fe;
reg [flogtanh_WDTH -1:0] Ia276ca65e85b9ccd4a9553b970b418a9,  Ic70b0be144931713bc160b7b4d8038e2;
reg [flogtanh_WDTH -1:0] Ia0b083b9bf3175a9961f79464d1b6bde,  Ic854870518bb942314f6269c6833ff5a;
reg [flogtanh_WDTH -1:0] I6aea13b6ec3703c9c919731b7c43e44f,  Ifdbf3e9abf7bff7ce4c689bb7e1226f4;
reg [flogtanh_WDTH -1:0] Ieb8b3cb38d28c4357bbd35d485f66dfe,  I4576ad4e2708a5635d93b304f1f10677;
reg [flogtanh_WDTH -1:0] I25fcdd6fea9bc9d728e5b6dc28cabee4,  Ibe54160f877c63dfaace0fc2c41ff11e;
reg [flogtanh_WDTH -1:0] I0ef97b8205f4a544cc31d1ab9fd62d90,  I04e75fe6916169cea741152b9fc6600b;
reg [flogtanh_WDTH -1:0] I157f4891b58262db67a57781e6789205,  I60fc524227900d3fcb19263336db4383;
reg [flogtanh_WDTH -1:0] I0306b43f29eb07e97472616ba7516f54,  I11555ad63e8caa81cb02dd9264668a3d;
reg [flogtanh_WDTH -1:0] Id8c72b2670ca8001c69b60551519f4b8,  Ie9feb0382e321c4cc1602c4fab33f939;
reg [flogtanh_WDTH -1:0] If32e24d0be817c10df587ed0aac48af2,  I21a1b05b4e659507fc3ff2077e7d2e8d;
reg [flogtanh_WDTH -1:0] I6c17cb40f5ab67595f89afc0aa3e570d,  I5af0b1d227ed007db9cd98d8a93b89a6;
reg [flogtanh_WDTH -1:0] I2789fbaed627ab6bea83080a0634f73d,  If9bdb9270926fe47e645cea702bf7775;
reg [flogtanh_WDTH -1:0] Id4415bf69046a95359a7f23a0ec3d5a3,  Ie6694b28f83262c5051dd00e336eb8da;
reg [flogtanh_WDTH -1:0] I25862ee3c8452b8f0d3187132477b77f,  I500e2c4d34270abc5a6f51cec578a7b5;
reg [flogtanh_WDTH -1:0] I5e8114931cbd9da66eec0a9e96b647b3,  I4c4c87637fc7973a58e933ffa76e611e;
reg [flogtanh_WDTH -1:0] I01a946c09a7ce0b62c7ba805e301de52,  Id7d81b33ad4bd7ae9df6a69b8e1e3351;
reg [flogtanh_WDTH -1:0] Ice805f2d2607178baf73b8c8bdd1b725,  I9eae9bcc567e9c051d268bd446b238ec;
reg [flogtanh_WDTH -1:0] I77767e8e8a46c270774c64d18eebca4c,  I614d496a5262a7f6ebd9a2d078ad30ac;
reg [flogtanh_WDTH -1:0] Iac7d03545a18a22c01e97d9f8ca93e40,  Ifdde7e51b6c92f13208685e0dc05c95f;
reg [flogtanh_WDTH -1:0] I1a60f16daa4667129838097d94c932b2,  I0ce07744582a47bf9cfcbdb2776a04c3;
reg [flogtanh_WDTH -1:0] I8f08550281859dc884c13197e046ef10,  I4b0ae6a7608a5ba8b1d66f7dac61bd11;
reg [flogtanh_WDTH -1:0] I23978d82bd6e911f5366f97765be24aa,  I6c2a048243ceddc9e31b7a37f74eeac1;
reg [flogtanh_WDTH -1:0] Ib26450dc355c3ca34ba704abe7350e2d,  I461cf1d25b347dd378a48f0dd2f5c5ae;
reg [flogtanh_WDTH -1:0] I29c302625d14d028e34ae65f37961e3a,  If32b0bc17ee8e3a95335b09550f05167;
reg [flogtanh_WDTH -1:0] Iede527989cec0a93d78423b7df14d707,  I2f751a32b067b688a98c0d98a8461265;
reg [flogtanh_WDTH -1:0] Ic0b1d8a6c00df4a35e285accfd1d149b,  Ib8528ee13f669ca3b7d0fddcc4fe697c;
reg [flogtanh_WDTH -1:0] Ic82e6892a22a0fd064bdfbe31cc171f3,  Ic0698d2eab5cdc70666a51ac0962e5f4;
reg [flogtanh_WDTH -1:0] Icd96d324832586b90e3d89709934fc9a,  I2ff4fa27b4aef5cca03eff8bb129a9eb;
reg [flogtanh_WDTH -1:0] I07aea291890873ea17e211143a7a8291,  I7770f02fbe5d3c1c49b9d5a3ffe4cd24;
reg [flogtanh_WDTH -1:0] I424af84f8e7d7f4c85fe9e4632d0a5b1,  Ib731ae113881b22a9abea15970d8c906;
reg [flogtanh_WDTH -1:0] Ied903684ae1a9f6b1d39d3714b6db7d1,  Iaef6a7213e546e24b635fd39c69b22a1;
reg [flogtanh_WDTH -1:0] I07e0123a7a61773a58a82d037140d1bc,  I5f2f0073edbf2de118fb329b9d2f6d2c;
reg [flogtanh_WDTH -1:0] Ideeabf83d0b70f18efb7a46d88efc352,  Idf85836a87828a65b1a189608df72380;
reg [flogtanh_WDTH -1:0] I148d4ff69853a123a3c5a306e978d9a2,  Ib3f304bc897f97659a51764e156f4002;
reg [flogtanh_WDTH -1:0] If578b689c5609b11df900bf92d0a388a,  I02c642372452e4dc5069ceb96098ff71;
reg [flogtanh_WDTH -1:0] Ibc5a4c442eab539e5bb136a83112191f,  Ie6a18db9c01142eb719b8426919a114d;
reg [flogtanh_WDTH -1:0] Ia19a1d1736d5feb515750e680b83db4d,  Ia96c18f8eef3c498f310b2aace71b9cd;
reg [flogtanh_WDTH -1:0] I98f9daa53631a03ce5f4d21fa499a734,  I94c6e4bc6b9ec661a6d76814aafa1e74;
reg [flogtanh_WDTH -1:0] I3a1a9a79b0dd6856b5d6ef8eda18c564,  I3c2369669172ef6a4f0a1b36916e4a34;
reg [flogtanh_WDTH -1:0] I9268175b692637227825c86f87dad083,  If22f0f17b0156ee153508c5e4c9742ff;
reg [flogtanh_WDTH -1:0] I1571e04768855319692febc19c86f630,  Ife58da9674cbcfa416675f629c158399;
reg [flogtanh_WDTH -1:0] I382b613b4744799d708ecb0c361c7293,  Iaefac912d485b61e57075ddb0212fc55;
reg [flogtanh_WDTH -1:0] I736ed9a09ea1b83b13fc3b53ded0c560,  I4b044f5c58a7d4eab6a1d2735e997f44;
reg [flogtanh_WDTH -1:0] I0e2430406a0c161380cfd60e7bbfa542,  I805cf823cf1cc902fe63131647d582c5;
reg [flogtanh_WDTH -1:0] Icfce7d26af22431c30d34d5738109a18,  I468c07efbe31fa2f18ae967a769e5db0;
reg [flogtanh_WDTH -1:0] I070f6f095b8a43ed92048d9fcd6625b2,  I68941b5c1b03152c7425aa0a1e347385;
reg [flogtanh_WDTH -1:0] I7b5d1412081b2bad3b5dd0cffe78238f,  Iee2c7d458d2673fe0cd58bcae0eca7de;
reg [flogtanh_WDTH -1:0] I04e76b2c5bf274bc2d8b9862c3690980,  I49597f093b8baac9c769fce82f7ad0d3;
reg [flogtanh_WDTH -1:0] I7fdb420f639b22294c896a20c8036f02,  I2f80f409a3c59f56aa230c393d6c4297;
reg [flogtanh_WDTH -1:0] I7a40ef6e10e3406e1d8c57ae53c6c3a1,  I87fcfc6fe1957f42e271128cfa0be7e0;
reg [flogtanh_WDTH -1:0] I2e3fbfe6dd237424289f6f4d00ad486e,  I37b6525d09e5cd2be4f64b64d380cf06;
reg [flogtanh_WDTH -1:0] I2cef2ca61302b60079b80fd9f252c56c,  Ib915a0bb2acae5abe82646277a50f211;
reg [flogtanh_WDTH -1:0] Ib44222bf07803a788687a877f1491ef1,  If7d1635e4aceeaeb897a2b9d03caaac6;
reg [flogtanh_WDTH -1:0] Id5fbe2f0dbe2a2d864202212c5db88cc,  Ib8ef3c757de68cd0afc90a6786286248;
reg [flogtanh_WDTH -1:0] I6f4cc724a3e77e3b282e08a162448b75,  I627418190ef1e1115d0346d2db6134ba;
reg [flogtanh_WDTH -1:0] I573fcd75e769729647bc1c5fc8e54852,  Id59e1e3a73e7db64fd4808fed9e3e173;
reg [flogtanh_WDTH -1:0] I806e05d43c46bf4f67ccf2f1afa2911e,  Iad4c43fc6e3ea0cddeb3da00b8faab4f;
reg [flogtanh_WDTH -1:0] Ia2f45ae7f344cf3de7a61fcc35ae4651,  I097da986a541504f1f641404c1749e43;
reg [flogtanh_WDTH -1:0] I3debb601b68a3cd58ecdaa7d78e66c7f,  If307175952944fcf9053a4d0eed964c9;
reg [flogtanh_WDTH -1:0] I9bc3698d4111848c8ff7f5082b4e6f3f,  Ib834d61619c282eb6994727f4b1fe2dd;
reg [flogtanh_WDTH -1:0] I4f5449753716964b3600bbcbd44902f0,  I9c6851db428c373c2fd723c1a374795a;
reg [flogtanh_WDTH -1:0] I39de7cf13d732f3d5c89eaa718407a97,  Ib815852a6d56c5ea21f7a23acb120f3b;
reg [flogtanh_WDTH -1:0] I1936f1a842424a3fdc777207a05433c7,  If80d97d0c5785dd6a0cd9fd3c0a6f870;
reg [flogtanh_WDTH -1:0] I2b5d24b895e1386c5acec6ec51af70ee,  Ifdff70e8ea00c64f13abd0d6da5bc11e;
reg [flogtanh_WDTH -1:0] I9cdec4376c54fd0d5892b20f7f3944e5,  I64fc41bf20b9f82b2bb86fc9f2438e81;
reg [flogtanh_WDTH -1:0] Ic3dc6389680526e4e9f3db1a31c4e954,  I303191eabaa2211774eb1341a7ce1d32;
reg [flogtanh_WDTH -1:0] I6de265c429ab7ef182f2ed2b52f413b3,  Ief8d6b623591a56818c091c5f08e9bcb;
reg [flogtanh_WDTH -1:0] I17dd943cac50d93f041a310edf916616,  I4fa399fc2e70ae442ef421db22b5ea9c;
reg [flogtanh_WDTH -1:0] I2a2db61ae5f793391b0388d1139c1003,  I4580e224188f11052c47c9d7d81178ac;
reg [flogtanh_WDTH -1:0] I3a4a24d886c2c06e283081c1b0079aff,  I3c484edf6cf740303824b22ad09ecdf1;
reg [flogtanh_WDTH -1:0] I1ae5bf5c035790ca6279076719f7d218,  Ic22fe13fadb6b0abb614918dd785552d;
reg [flogtanh_WDTH -1:0] Ic98fdc1a35fc3c698dd9c5bfe2fdd1ac,  I015c6af005c8eb5a6ccdf97fd0073bbd;
reg [flogtanh_WDTH -1:0] I0b771b927e8acb823e30239c89aafe9f,  Iee7fd00e1644e71903c0ca268ba813ec;
reg [flogtanh_WDTH -1:0] Ic3caaaecbbca186ebf9cc35e554ff62e,  Ic9143d7200fec6ef38e6cde1fc13d859;
reg [flogtanh_WDTH -1:0] I33fc4ecd929152c59d62af65ecb38414,  I974755cb3f16a1db503e4d6658d1f4bd;
reg [flogtanh_WDTH -1:0] I09a3008676f21e58545563dff1cc9328,  Ie7d8d3754dc7cc7ac9fc8ebcbd3bf82a;
reg [flogtanh_WDTH -1:0] I566a0851428acd33e432b33fe3c42b4c,  I903284ce681f1526c56a4889306a65ec;
reg [flogtanh_WDTH -1:0] I96884d5c0babd2437ec14429856c0414,  I2e1e3933f8ec5db47edbec59fd1772b5;
reg [flogtanh_WDTH -1:0] I6a3539539860b98d7a310f63314a2932,  Ieccf95256e095c0e79b8ac959cea7655;
reg [flogtanh_WDTH -1:0] Ice31c844af4b8c3b966b778cca601527,  I5c9eba93bf9c01e161dd3bd508980acb;
reg [flogtanh_WDTH -1:0] I8eec3d66ef763226b960a24192aafe27,  I8f66edb2bb1d6c6f228711fc27836a3d;
reg [flogtanh_WDTH -1:0] I093a0ecd0a1aaea8a97d08d54cd37fec,  I0be6fa3f4ae264a84a3b241edd706034;
reg [flogtanh_WDTH -1:0] I3b2708fccba619958a392242efbbeea7,  I7fa9026688537d119b6997572564584d;
reg [flogtanh_WDTH -1:0] I543deb703bb9eb808f4381f543e408de,  I501a61dbbe9a6edfbf51d18b14d96f10;
reg [flogtanh_WDTH -1:0] I0e0c7e753509c664971fd12be9183537,  I4fc839b634aaa2e0b5775984e0dbf6ae;
reg [flogtanh_WDTH -1:0] I68577e7dec24946ec0745c5d4255795f,  I9a432f4a190d752c5e723107243daa1d;
reg [flogtanh_WDTH -1:0] If53e38b5b6031a7e927a65f90acf5120,  I23a1b8a01fbaa3122ef3d1efe362a3ff;
reg [flogtanh_WDTH -1:0] I372a38a8675f65c5257b645fb5d809af,  I97a78caa8c75ef80934e8d013fee43a4;
reg [flogtanh_WDTH -1:0] I0d37309bb37b707e10a4e12425157fe3,  I72d4a7275ddf3d5d41149fbc6e6cce23;
reg [flogtanh_WDTH -1:0] I5935a4ee604a8c6259d88bd4b679babf,  Iaf87541d81d0e3cefb78aecf3ae9c92f;
reg [flogtanh_WDTH -1:0] If4ed201fbbaa5ce9bfd05d65d79458d0,  I55ebb5c7ded985c8911629524e62aa16;
reg [flogtanh_WDTH -1:0] I9b11c7aa2d35ee4589dec055ab0df2ca,  I19a49d3680e5786fad7060cbc4be4a16;
reg [flogtanh_WDTH -1:0] I45a6d3691aef6c693ae6ee25c25a4b24,  I60e4a3789fb3df162298306c815259b2;
reg [flogtanh_WDTH -1:0] Ia15364dea1e0f0243204b4bc4c9b8bb9,  I25054529bc0fe35bd08f6294a2d51f5e;
reg [flogtanh_WDTH -1:0] I2f31acde416c079c48ce54697eac5e60,  I8a471bd6f3fd220a34d9cc870eaeafe4;
reg [flogtanh_WDTH -1:0] Idab577631403b170aa07d02c7d455315,  I12d2ea504991199ca905ca91925f2d26;
reg [flogtanh_WDTH -1:0] I36b79e4befc1673140076d2f9cbc9d82,  If93a23874096c597803aa347c0900cd2;
reg [flogtanh_WDTH -1:0] I9f263275a24efe9297aa995282c48360,  I5f3af0ef6d4722a508201707b6994fed;
reg [flogtanh_WDTH -1:0] I7915e8a9a775ea1bc1bf7fe71648303d,  Ib88cf5d737b09afb18cbce8072be2ea0;
reg [flogtanh_WDTH -1:0] I4a7ac8c9709967341ededa935aa65581,  I626fef2cd9d071cb8c797471055cf245;
reg [flogtanh_WDTH -1:0] Ibd7437a655d4985728ce070004e3b419,  I723088e5c9b31e731220874d2f27f195;
reg [flogtanh_WDTH -1:0] I8a834fd9d1425a79f7ff0713777fcdcc,  Iacdb27c060a48b7ade76d256e858b314;
reg [flogtanh_WDTH -1:0] Ia60cc135f03b89516e61d52335e69674,  I3719da3863fb069e898484ce997c2f40;
reg [flogtanh_WDTH -1:0] Ia1b1f012b02265afed03cb146e88f2a0,  I3dfcd0d247d56f8167bcbc6aea6e3504;
reg [flogtanh_WDTH -1:0] I6095ee8675c10be082abccd7cef7ceeb,  I477e8f9e2ac8c5d142856ec6787e28ac;
reg [flogtanh_WDTH -1:0] I2be07fc5652209f0e8eda31090dbb162,  I2865e7f35c36e2cd4a4e3435aa8c7c14;
reg [flogtanh_WDTH -1:0] Ic60fc4bb6e7ccb8bee260e5b982bc5a1,  I4d83852d202e9f1c49955b59d183cc07;
reg [flogtanh_WDTH -1:0] I217d1876f768c7dd3eed096e2de59dfd,  I7d5b2a7bca99f2164a7ba2cfe46b20e1;
reg [flogtanh_WDTH -1:0] Ibb297f22ba2e0d4786042f7503ff3f61,  I3c7c5071212ff5db857e3f84f6131391;
reg [flogtanh_WDTH -1:0] I8d917a51d32729f4a5a98b5d3a40f947,  I6296deff598d27ebc1a06cb1316a3eb4;
reg [flogtanh_WDTH -1:0] I08213a1a86aa27e3d3ed2d294d972ea7,  Ie6acf5390a3487fca3f8e4b66a640da3;
reg [flogtanh_WDTH -1:0] I271dfdeef4359fa9b2ebf80ca950a08e,  I6a993db6733d3efe90511bbe7f4d5654;
reg [flogtanh_WDTH -1:0] Iff44a32b2e9a1a65d820b0839313015e,  I3ba62f936f0832ff2ebed33f862286ff;
reg [flogtanh_WDTH -1:0] I2882587956babd713eb3a53af6afe389,  I0f8f8ce5dfbc020b547758c239f923c4;
reg [flogtanh_WDTH -1:0] I4f1ca888cae3ee3efeefafcfb12e16b3,  Ife2ceb6bb50cdc7adb4a20e1851d54c5;
reg [flogtanh_WDTH -1:0] Icff2aa823d2f0e9421f3fbce6d21f510,  I361c911024ff757958306a38c4bf4465;
reg [flogtanh_WDTH -1:0] I2cd19bf0afc4563ea24619849ab7d8b7,  I8ca3c12dd3e04f05ca52ebd1ea32cfee;
reg [flogtanh_WDTH -1:0] I80cae65874911e05bc77db3e5fe0fcd2,  I56a419f6f3b841e7e5dbbbcc0e6af190;
reg [flogtanh_WDTH -1:0] I18c43491892bd258dfd07aa0263c5479,  I5ee41fe39af22ebe82e91a1dee0b7221;
reg [flogtanh_WDTH -1:0] If322bf2a59be9bf7b33a49a6baf72ed7,  I807e19c30c0328199d5ab2d64593d509;
reg [flogtanh_WDTH -1:0] I2bb21cbf03db27c0b9d814517033b56e,  Id4a5425f6a2a8a689eb1e5e25131fa0c;
reg [flogtanh_WDTH -1:0] Ib408b39624c6576c228f32eed26ccf8b,  I2ba381005b1ffbcf163c40f2dd92d2f9;
reg [flogtanh_WDTH -1:0] Ib6dee36145f77a6f1364c218140266b4,  I2a48609c13ebc0cc9a8551fdf244a2d8;
reg [flogtanh_WDTH -1:0] Iafa25738d96fb115c78d8d295902c263,  Ib0db88e9d645459a03e908dbbf6b5803;
reg [flogtanh_WDTH -1:0] Ie7cb395e7ce65ca399d99a5e62a7efad,  I9170cf346273d705158f36c2a9e59961;
reg [flogtanh_WDTH -1:0] I1bee0c6e3a24ee319d219799ce58f13e,  Iec7ceaf0d09a3629dbe42f8926383e83;
reg [flogtanh_WDTH -1:0] I7fcbf3d532ed0c810cdc1c5be536d263,  I9d738422a85fb3cd648444a039b96e9d;
reg [flogtanh_WDTH -1:0] Ied7f9cbbcacc43332f1219e8bd0a07bb,  Iece0c68af7dff6bbe73e9e2d468585c2;
reg [flogtanh_WDTH -1:0] I491888fefe23bb0bef60f293668491af,  I66f0d7b1c32cba28b55806d443090f9f;
reg [flogtanh_WDTH -1:0] I1b9368c7a0d236ed73a6783281144bca,  I3d2bc0bd4abfa1286242b841ef4f04ba;
reg [flogtanh_WDTH -1:0] I2adf1f34eb55f6f7e5f37b328b2bcf21,  If83620428cf14f11cbd5eb3584a0e877;
reg [flogtanh_WDTH -1:0] Iaa61cf5ca911de351708963438768cee,  Ib9161bcd780dcb77507b4851bb21193d;
reg [flogtanh_WDTH -1:0] Iacba64081faa56ef9190aa65fc89ae7f,  I584c580e66ed2d89371a7a1a4fd59599;
reg [flogtanh_WDTH -1:0] I5d41596aeb3aeb4f07dbc0c995b5f4a3,  Ie3ac6cf6fedf997b6839abbcee584fce;
reg [flogtanh_WDTH -1:0] I1c01c903faacd546e44a6fd6564ef3bd,  I3a67256306c29f917d28ff55be76d4bc;
reg [flogtanh_WDTH -1:0] I3e3195b93f03e3c8c24655259f745374,  I8506a14aacf97d360aa4c10a91ef184f;
reg [flogtanh_WDTH -1:0] Ie229e972daab0a41969c5cc066e52e61,  I6751092e3a762e4f0ac88e02e8d145df;
reg [flogtanh_WDTH -1:0] I5a646f85f9e6d52063b0c0e6f479f6f1,  Iaf3e9f18da33e20e42838b4467d9741c;
reg [flogtanh_WDTH -1:0] I01a50cb46ae1b229eda9094867090aae,  I83649a386aab66f1c0774263a77831c7;
reg [flogtanh_WDTH -1:0] I68026b1eb748133551563bea029c3488,  I8ff4739a83ed374704f039515b99162f;
reg [flogtanh_WDTH -1:0] I726047b0a4d45f8ad1f394301dbfb78d,  I9851d75a6dcdb74212fd0146a9aa49f7;
reg [flogtanh_WDTH -1:0] I2cddfa0b89e0aececac2dd7d983beb26,  I9653890e840ec994e81844c9a34b10ba;
reg [flogtanh_WDTH -1:0] Ic5e1dd806582ee08eb6d1048d6617b13,  I1322f065e413aef275747decaa48d550;
reg [flogtanh_WDTH -1:0] I9040f68430c75ce7527990dd702b7feb,  Iad493aff89cf569ffcc57b8f204c11ad;
reg [flogtanh_WDTH -1:0] I40ebb4eb571f18c2fb810daab0d5770f,  I99928f669eb8b23feb022a8fb39ef5f6;
reg [flogtanh_WDTH -1:0] Ia4738ee511867aa46e0e92f3d86c4ccf,  I98207474d16dc958a7e695a56a81b614;
reg [flogtanh_WDTH -1:0] Ic10326eae7434399af6e611e31389963,  I422a5ea4034e59d308907e5684f8ad8e;
reg [flogtanh_WDTH -1:0] I8fafe7fe582d027b97dbf2cc58763096,  I2911a1c5c49beebcd2fe684678ab89ca;
reg [flogtanh_WDTH -1:0] I8a329168f83731c15dbedb1f1f966d78,  I0a3206015f8d35fafd10bd4709b95faf;
reg [flogtanh_WDTH -1:0] I603a5f82891f62b59f7890d631d0b6df,  I10d423113bbfd394aca2695798b2d4ad;
reg [flogtanh_WDTH -1:0] I620517db078658289fcde4200f15ac06,  I596999303fc894014a5ae6ba2f09f143;
reg [flogtanh_WDTH -1:0] I51271c02c6fd9cbda153c9b28aa099e3,  I1e24b9c9e023b6f0b00cdeaa071366a2;
reg [flogtanh_WDTH -1:0] I8def31183d1a648a6a50245eeb6b57a1,  I6983ea7dcebc925bd95ee96457a2de66;
reg [flogtanh_WDTH -1:0] I0c3a1185a9fbb05c0dcec0d655068786,  I3d0c2d0d76d54c59e1d282a37e0aeae8;
reg [flogtanh_WDTH -1:0] Icf0284aeb5d603e893733d2139a79ef3,  I6f6c9a635c0ad62e7687a666f98ca4d1;
reg [flogtanh_WDTH -1:0] I3d0e6fa7f7edbd105fd8f7823722bcf0,  I929ddfd7ec9bf7b7c2dd2378395a403a;
reg [flogtanh_WDTH -1:0] I55e28dff0ebd1007f4f00c512f1df1b7,  I6fce04d1f8c9975afa3e6abb203b13db;
reg [flogtanh_WDTH -1:0] I2b33fef3c83dab2f2d254cb295264482,  I88d063cb6f169e9f1ae067641fc0d802;
reg [flogtanh_WDTH -1:0] I1689bfa3340ff4798ef7eb160714ede5,  I2adbad4296c06db0ef231d53e6516986;
reg [flogtanh_WDTH -1:0] I1b5deee5754dcc0762ca2691fd927056,  I4b139847ca9cce5281ceb1d63a453d05;
reg [flogtanh_WDTH -1:0] I1e63fce77120b91dc6195d2febce4d42,  If9c81e3f27ee171ff282cc7fe18947ed;
reg [flogtanh_WDTH -1:0] I1d3f5624cb6f217fac422833ed8b7195,  I7648b4562836acb77aebba8b19dc62e8;
reg [flogtanh_WDTH -1:0] I1fde6652c1fb298d84e88620edc9e91a,  I9f2892cd4e16b8719b5ffcb4b051ac0f;
reg [flogtanh_WDTH -1:0] Iffd2d0fd17d604ddadcfc2dd9e46276a,  I159acdea94fb6185fccd6310e9d1b071;
reg [flogtanh_WDTH -1:0] I8295b6fa92e241d4b689ad0e26f6a2db,  I7a19ff6c711f9ed53df05a4999041a70;
reg [flogtanh_WDTH -1:0] I8573b3db0d36442c2f233d12586d82f5,  Ifa65fb0d14e454b62f138630d2f9f370;
reg [flogtanh_WDTH -1:0] I5319144e65be1e69c9ef767bfecd4ea3,  I0f24875d6dcbc0c7c83602f50ee3a8f5;
reg [flogtanh_WDTH -1:0] Ie7da9e9fdd626504cb2f00a3ec899718,  Ic888c593409b429e20523b414861da69;
reg [flogtanh_WDTH -1:0] I8293d7dc145b31d28c05c02677760e9a,  Ic10e70c69f2401950c31aeaaa1600ed5;
reg [flogtanh_WDTH -1:0] Ia372f6e388ed5cf8e9810c52d3749136,  I3c6576aed9ae9c1a1e86afdc00082fc0;
reg [flogtanh_WDTH -1:0] Ibd959e3bf9ef7ee76ec2754a06926d9a,  If710661738ba49d8040a1aaa6c4a0dfe;
reg [flogtanh_WDTH -1:0] I8f03815159c11486a4805e7f72c84a38,  Ic6e2dd06abadb6b0613d8be1d3e91da7;
reg [flogtanh_WDTH -1:0] I15e5e06b7dcf6616094faeb798a0fdc8,  I6e72837b363b91f0a1301ccc2c3a9e32;
reg [flogtanh_WDTH -1:0] If23f4bc5d45a3e7a22a9e8596b99c575,  Ieb48cc2ae37e2d9dd9144b587cce78da;
reg [flogtanh_WDTH -1:0] I70afe2bb83173aa96269271270d03f2e,  I0c2ea6ea58ccc53502b8765d9ab08a56;
wire start_d_flogtanh0x00000;
reg I2590acd159fd90fe367126ce432e39e8;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I371284eed470112cb89e1d361a9d40f7 <= 'h0;
 If0fb2e90431d89d99912918f83036f4c <= 'h0;
 I0ee915f21334d38c75f0207e3b052a69 <= 'h0;
 Icf5a9bd712d310ac17eb2354f884a237 <= 'h0;
 I3222cf2f98878be3f453560ddb3dc43c <= 'h0;
 I2dd9e89f2842e748c1574ad0e7f4dba9 <= 'h0;
 I667adc16c92bec8f413a1a9bbfc41ce5 <= 'h0;
 Ie6aa50a44574542826b78fed7d77b76f <= 'h0;
 Ie97072fa52f483bbd89f019c21152cdf <= 'h0;
 I47f153e1cecaa77f1e6e6f07c0220557 <= 'h0;
 I1b9dcfaf144b48a64b990e5b020d4a02 <= 'h0;
 Ie32d4bd927d02e547850331db8028177 <= 'h0;
 I0988db7ca497541e372131a0b0e8075e <= 'h0;
 Id13b5577b8baa586fedd34d4aab9d9c5 <= 'h0;
 Iedd0e0f6ee682a131d4f14c4762ea0eb <= 'h0;
 I875d7c55914414298f0fbec0b345c92e <= 'h0;
 Ide64c9647c7898867e0d036e9ff95f6e <= 'h0;
 Ied6ccabb348ed7e20567011e027c86ad <= 'h0;
 Id030b072054c623c7aac5c571d052951 <= 'h0;
 Ice55fb2e506accf518b4aa18298d017e <= 'h0;
 I07a0167dcdfc76612e1b0da251337a7b <= 'h0;
 I045e08f48738d395af2b79f25af73732 <= 'h0;
 I7df57f27a880fe45f78c108f8faba963 <= 'h0;
 I60204c1d3a96524bbbdf715f95f08fe4 <= 'h0;
 Id5b9ae91dc900060caffff2520236f66 <= 'h0;
 I861fe9da6d004ce3998ab54a8c0d62af <= 'h0;
 I95caae0432aeadc0cbe279f9d6f9062b <= 'h0;
 Ic9c3b015d5830bf4834a435eba89caa5 <= 'h0;
 I6e18dd1a579e09b80ac113fe85b483b4 <= 'h0;
 I51c1c8e8df14396c5c77b5013531a84f <= 'h0;
 Ie8f75e8e020d43f6a357b5175047c254 <= 'h0;
 Ie762d8aa151448cbaa0d005a3c01572a <= 'h0;
 I293b32c043e20d6baab178319dd1e2f6 <= 'h0;
 I200aae813b664e02075eeefbc3b4450d <= 'h0;
 I006264bde45d8df078ef711c221ff387 <= 'h0;
 I9200a0071528b14dc52e92082768ca97 <= 'h0;
 I55761decd7043b4dc82737b9d6ef6e7d <= 'h0;
 I4f51d114002bdfd69a31f95c2fa5234c <= 'h0;
 I796cb71b28957405c10015a2ab7124c6 <= 'h0;
 Ic85bacce5db48b4dd3f626749f6effa8 <= 'h0;
 I2a508066cf0e07bbe8a91f276fbb3078 <= 'h0;
 I85913ae95fcd63de45030d583846b1d6 <= 'h0;
 I971cff06a60916ea3e136b397d4c620b <= 'h0;
 I2c363f7abf62c9026d0b0dfe5a51207a <= 'h0;
 Ia5043b0c8ee086c66e683eb115a75484 <= 'h0;
 I6b7b63ea23c5b4f3c597f121284cd2da <= 'h0;
 I3cf82abadcee2faa1849d0a9a45b051e <= 'h0;
 I8b42f5455dd8f6323d7a4e28c0eaa1a9 <= 'h0;
 I608597017b046d92b77226999df90600 <= 'h0;
 Ia39b908f8d6b63777376ca560cd0cc8d <= 'h0;
 I87ad38ab473927df7c0bd69c6b4b4c5e <= 'h0;
 I8e70752f74ecdbe95a7b33ca264d4589 <= 'h0;
 I6e768e27a3f1804919e3f83c050e19ba <= 'h0;
 I2285f424ef2b8b2041267c1652155ad0 <= 'h0;
 Ibc5b97632aab1e763ac51f8d18edc792 <= 'h0;
 Ic4a0165bd71d9e586fdc66c824e45224 <= 'h0;
 I40de7aeac837276e7b3f0c4b29ce5eca <= 'h0;
 I024a746142e5ff074724f92af62f3bd3 <= 'h0;
 I1e54f934fa92e681472d03199991f0b2 <= 'h0;
 I8cabd17b81e99a86fc8704aaaae629a3 <= 'h0;
 I54c1bf986182c83540d950762048a5e3 <= 'h0;
 Ia5fbeb5be349b8088a749e25a9e6e416 <= 'h0;
 I987b220a4729d14e9fc97b57867436e4 <= 'h0;
 I7f1d9309d3053256134130574b970425 <= 'h0;
 I9fd9d5a2a3a34b532bad740b16ce66fb <= 'h0;
 I66a648a9f6b10b1d580e72b36a1ed9e7 <= 'h0;
 Ia08c041d1aacfbbd1f8d7980923b9b05 <= 'h0;
 I6805a2f26b1e51f7ac0087e6829b3c5c <= 'h0;
 Icc11f9d183454b33624bd411710342a0 <= 'h0;
 I18f145bedd3864fcebd983f9533a5877 <= 'h0;
 Ifa25d4c9ccc3efd1af4e711d3c32e9c5 <= 'h0;
 I5bbf8f01c5ddaa02516dde3867ec3d78 <= 'h0;
 I3f8fe2d052a6df20dfaac6f88d4fff8a <= 'h0;
 I9fbf9bcb6022bb550bc2dbd52f20d05f <= 'h0;
 Iacd71ce5854c85450463a0a45ebc6a2d <= 'h0;
 Id7c1a8f42cc90b7846105cd103b07228 <= 'h0;
 Ic6d94b59cd6f4c7765463694c9fbae3c <= 'h0;
 I11a9409c814372a31d771888692ae955 <= 'h0;
 I760f9ff7bc594c98e71080485cc1a082 <= 'h0;
 Idb9be12ba6807752b0c36f4cc18843cb <= 'h0;
 I192119ad6ad1396dd6fd1fab6e4c4cca <= 'h0;
 Ib4c62a865f79eaa2aa5fbd12860f2e80 <= 'h0;
 I5fb195f29a4e02620d2cca6e7f2a8fa0 <= 'h0;
 I41b4d1d3d5ae22c8fe4f1e0fe20ccac7 <= 'h0;
 Ib2afa3be272607c236cbd5410a88e8c2 <= 'h0;
 I43587e6827dc7dc1ef38d552f6a73ca4 <= 'h0;
 Ic27ed0f98cad254a72ade8253ccc01d2 <= 'h0;
 I5860a511728dad8112a9246843f0fdab <= 'h0;
 I6f83f4d8681a17b7e700a38a78917822 <= 'h0;
 Ic902ce884c81efed3160715af43eb19b <= 'h0;
 I8297012f23a474aa863c56e6ab9f77f4 <= 'h0;
 I703fa28fdfb32f8e7fe5062a3332ff6a <= 'h0;
 I4d60a4630a93dbf6460fc525f16fb69b <= 'h0;
 If6a1f518420fbc246e2524469689a5e7 <= 'h0;
 I48c55cdc6c1e3bb5e36a5451cb43c5a9 <= 'h0;
 I147accfb14f15341869779b74c8cadb6 <= 'h0;
 I0d302535ee6928ed74d7b456efaf01e6 <= 'h0;
 I0039a78cbf75de3d875c319e3bc08d22 <= 'h0;
 I7a43154a62ef625844cda08b1dfc9c79 <= 'h0;
 I8e05a477fab7c0c6f70c681626640b93 <= 'h0;
 I51393ac63dc5f8c0898ffa6dd59ee183 <= 'h0;
 Ib4f7dd6e43c7a291d753f96b1aac8ce6 <= 'h0;
 Ibf76adf5511e851727200f4fd60bf34b <= 'h0;
 Id90de24703e5b15356a8ab3862612957 <= 'h0;
 I2b42badcbe3d18d033edbd6d4663fac6 <= 'h0;
 I72450aa2c2f2f501a5465f008e95ba4f <= 'h0;
 Ib802f2c9c1265a47e5acfc419034488d <= 'h0;
 Idb28449172f54add7ac6fd1287543a5b <= 'h0;
 I6b33174bb2786da0ba9ba988a96aa5bf <= 'h0;
 Ib68892cce1de9f46fb391a7ee8a01afb <= 'h0;
 Ia0e39ef7db11ff2f95f50e6a912e945e <= 'h0;
 I1f3153881fc6a7fc767a33253f80e06f <= 'h0;
 I994e4d13d16c12025cb60205b8f7559f <= 'h0;
 I3e4b2dbb8f44350c5cff7430502401b7 <= 'h0;
 Id1e6e9ac8ddad3aedd347aee9f615d9f <= 'h0;
 I5a6da3732e0f265ad95269f5a629c1e8 <= 'h0;
 If8773fa380ec5c1199794d4128d443f1 <= 'h0;
 I63283e5286a737d3ba1f99ae29902bb9 <= 'h0;
 Iedcc3a589dba858f1193b1be582db24b <= 'h0;
 I8a87d3adcb2989738d70db84c3b97a3a <= 'h0;
 I267e058f7db05744d80df6b52be83475 <= 'h0;
 I5e121581d8a5f81fc84da2fa982d8fd6 <= 'h0;
 I51f875fbf103d8b8093d73279f127843 <= 'h0;
 Ifcbf9c1d4d6f111f06212e58764d29ea <= 'h0;
 Ie0e816b57f511fc0479210deebbd9fc1 <= 'h0;
 Ia7673dc1d477d486371935040ff7dce9 <= 'h0;
 I7df5c4ad52bf35d254a4a14771a28fe7 <= 'h0;
 I9ae2d00bf699c7f12c3f5d78ad2c405c <= 'h0;
 Icb740a93e2adc0a9f18ac25d0c5d018c <= 'h0;
 Ia9691e7c587528f3ca0d85d842225da4 <= 'h0;
 Iab732884bb2d4b1781e31c7a1c109000 <= 'h0;
 I67d8e4c822cc57b150a76dbb3478b5b5 <= 'h0;
 I3bb2f03bf7d2f7480187062b45c6fdd9 <= 'h0;
 I8e57236f80078ae72706aa8102e1bf53 <= 'h0;
 I1732bcc59b7bad3d08b232d099fdefdc <= 'h0;
 I4b568309171ac557250c2ec600b9d7b0 <= 'h0;
 I886251a3307e5fe20788c8e947f4ef37 <= 'h0;
 Ic0d064e8436ad001f7e9d97e800e5636 <= 'h0;
 I9f2ba5b0600c5eb81cef40d0822d0aea <= 'h0;
 I2aaf6ff0daa3d3e26b197e6895cabf3c <= 'h0;
 I2e8c68a51f1f1f4e413897791a6823a0 <= 'h0;
 I1a318a04ba3cf92f4ba0dc132a564040 <= 'h0;
 Id32b88b33bfbcf79ff0a10d447f69619 <= 'h0;
 Ia41215dbdcd4b27a8ab41f48d40d644a <= 'h0;
 I53c239961c5745db892194a0a62b5d57 <= 'h0;
 I0ffed4dfc4e97bb477647e5eab3a18f3 <= 'h0;
 I46fcaa5311cc831199bb4a5a3dba797e <= 'h0;
 I69b693e03eccfe9a889894988c0c9a53 <= 'h0;
 Id0ca109680ce0cb6603139baeebac59f <= 'h0;
 I7bcf3409fb1f7bf880f945db8f2eb6c2 <= 'h0;
 I873254d95f4a9976acf9210228365521 <= 'h0;
 I2a437c10a562e8e7f4cef30bbfde2fd3 <= 'h0;
 I50e26d2184d04613f297357308e7c91e <= 'h0;
 I8b14ff6b303ae081ae414ca7a00da3eb <= 'h0;
 Ibf3a99967d7cbab53676fed78da28eb8 <= 'h0;
 Ifb6cf60f578b5a5dd0c27da72408cbce <= 'h0;
 I000bdba9ccdb068a02fd37d2991675b6 <= 'h0;
 I5110f5370812f6d0319c0f42a6638b5b <= 'h0;
 Ic36cb86884806afb677ac8fb42aead36 <= 'h0;
 Ie4dba51278ebf8a9358c2019383fbaf8 <= 'h0;
 I96373fc8bdf40551ef8206b4ba38cd98 <= 'h0;
 I7b8a50810f6a4c27a23c82330707c4b6 <= 'h0;
 Id84a4cc9f82244c2357edc537824eb30 <= 'h0;
 I8866b1e80ead799943d3ad273ee0c97e <= 'h0;
 I33d92c1bdacf71fa60865f1741288cdf <= 'h0;
 I834a4a93056d8777cd2d4996ae33122a <= 'h0;
 I51bc583f480542f3f95241643bb39eee <= 'h0;
 I35539407bedb7d43642e952787216ce6 <= 'h0;
 Ifa78beaa6ae7a7a32f4886a14e4d1532 <= 'h0;
 Iae691c305b2fd52617ef92705568a8b8 <= 'h0;
 Ie87c6bd3452b53ef57df5f420f351434 <= 'h0;
 I03106ddaebe00bc59e1611573835f727 <= 'h0;
 I8b947b6c3139066fbd5873d5b818183e <= 'h0;
 Ibb1c668cb8ad3eb49b9bff842d118aa7 <= 'h0;
 I4c3bda40c1fe5dbacee1829e0d60bcab <= 'h0;
 I405504d762cd698722b183721df7243f <= 'h0;
 Iae9c6245aa98b5758df6d57f8c33ab31 <= 'h0;
 I35f897e994d6fb9ae452bee5b423c4e9 <= 'h0;
 I413a7fe2255064627ed283d35d910de4 <= 'h0;
 Ic930f61e087bf2477712e8fef9c413d3 <= 'h0;
 I61ce1d41fa5221c01f7e9571965eb3fe <= 'h0;
 Ic70b0be144931713bc160b7b4d8038e2 <= 'h0;
 Ic854870518bb942314f6269c6833ff5a <= 'h0;
 Ifdbf3e9abf7bff7ce4c689bb7e1226f4 <= 'h0;
 I4576ad4e2708a5635d93b304f1f10677 <= 'h0;
 Ibe54160f877c63dfaace0fc2c41ff11e <= 'h0;
 I04e75fe6916169cea741152b9fc6600b <= 'h0;
 I60fc524227900d3fcb19263336db4383 <= 'h0;
 I11555ad63e8caa81cb02dd9264668a3d <= 'h0;
 Ie9feb0382e321c4cc1602c4fab33f939 <= 'h0;
 I21a1b05b4e659507fc3ff2077e7d2e8d <= 'h0;
 I5af0b1d227ed007db9cd98d8a93b89a6 <= 'h0;
 If9bdb9270926fe47e645cea702bf7775 <= 'h0;
 Ie6694b28f83262c5051dd00e336eb8da <= 'h0;
 I500e2c4d34270abc5a6f51cec578a7b5 <= 'h0;
 I4c4c87637fc7973a58e933ffa76e611e <= 'h0;
 Id7d81b33ad4bd7ae9df6a69b8e1e3351 <= 'h0;
 I9eae9bcc567e9c051d268bd446b238ec <= 'h0;
 I614d496a5262a7f6ebd9a2d078ad30ac <= 'h0;
 Ifdde7e51b6c92f13208685e0dc05c95f <= 'h0;
 I0ce07744582a47bf9cfcbdb2776a04c3 <= 'h0;
 I4b0ae6a7608a5ba8b1d66f7dac61bd11 <= 'h0;
 I6c2a048243ceddc9e31b7a37f74eeac1 <= 'h0;
 I461cf1d25b347dd378a48f0dd2f5c5ae <= 'h0;
 If32b0bc17ee8e3a95335b09550f05167 <= 'h0;
 I2f751a32b067b688a98c0d98a8461265 <= 'h0;
 Ib8528ee13f669ca3b7d0fddcc4fe697c <= 'h0;
 Ic0698d2eab5cdc70666a51ac0962e5f4 <= 'h0;
 I2ff4fa27b4aef5cca03eff8bb129a9eb <= 'h0;
 I7770f02fbe5d3c1c49b9d5a3ffe4cd24 <= 'h0;
 Ib731ae113881b22a9abea15970d8c906 <= 'h0;
 Iaef6a7213e546e24b635fd39c69b22a1 <= 'h0;
 I5f2f0073edbf2de118fb329b9d2f6d2c <= 'h0;
 Idf85836a87828a65b1a189608df72380 <= 'h0;
 Ib3f304bc897f97659a51764e156f4002 <= 'h0;
 I02c642372452e4dc5069ceb96098ff71 <= 'h0;
 Ie6a18db9c01142eb719b8426919a114d <= 'h0;
 Ia96c18f8eef3c498f310b2aace71b9cd <= 'h0;
 I94c6e4bc6b9ec661a6d76814aafa1e74 <= 'h0;
 I3c2369669172ef6a4f0a1b36916e4a34 <= 'h0;
 If22f0f17b0156ee153508c5e4c9742ff <= 'h0;
 Ife58da9674cbcfa416675f629c158399 <= 'h0;
 Iaefac912d485b61e57075ddb0212fc55 <= 'h0;
 I4b044f5c58a7d4eab6a1d2735e997f44 <= 'h0;
 I805cf823cf1cc902fe63131647d582c5 <= 'h0;
 I468c07efbe31fa2f18ae967a769e5db0 <= 'h0;
 I68941b5c1b03152c7425aa0a1e347385 <= 'h0;
 Iee2c7d458d2673fe0cd58bcae0eca7de <= 'h0;
 I49597f093b8baac9c769fce82f7ad0d3 <= 'h0;
 I2f80f409a3c59f56aa230c393d6c4297 <= 'h0;
 I87fcfc6fe1957f42e271128cfa0be7e0 <= 'h0;
 I37b6525d09e5cd2be4f64b64d380cf06 <= 'h0;
 Ib915a0bb2acae5abe82646277a50f211 <= 'h0;
 If7d1635e4aceeaeb897a2b9d03caaac6 <= 'h0;
 Ib8ef3c757de68cd0afc90a6786286248 <= 'h0;
 I627418190ef1e1115d0346d2db6134ba <= 'h0;
 Id59e1e3a73e7db64fd4808fed9e3e173 <= 'h0;
 Iad4c43fc6e3ea0cddeb3da00b8faab4f <= 'h0;
 I097da986a541504f1f641404c1749e43 <= 'h0;
 If307175952944fcf9053a4d0eed964c9 <= 'h0;
 Ib834d61619c282eb6994727f4b1fe2dd <= 'h0;
 I9c6851db428c373c2fd723c1a374795a <= 'h0;
 Ib815852a6d56c5ea21f7a23acb120f3b <= 'h0;
 If80d97d0c5785dd6a0cd9fd3c0a6f870 <= 'h0;
 Ifdff70e8ea00c64f13abd0d6da5bc11e <= 'h0;
 I64fc41bf20b9f82b2bb86fc9f2438e81 <= 'h0;
 I303191eabaa2211774eb1341a7ce1d32 <= 'h0;
 Ief8d6b623591a56818c091c5f08e9bcb <= 'h0;
 I4fa399fc2e70ae442ef421db22b5ea9c <= 'h0;
 I4580e224188f11052c47c9d7d81178ac <= 'h0;
 I3c484edf6cf740303824b22ad09ecdf1 <= 'h0;
 Ic22fe13fadb6b0abb614918dd785552d <= 'h0;
 I015c6af005c8eb5a6ccdf97fd0073bbd <= 'h0;
 Iee7fd00e1644e71903c0ca268ba813ec <= 'h0;
 Ic9143d7200fec6ef38e6cde1fc13d859 <= 'h0;
 I974755cb3f16a1db503e4d6658d1f4bd <= 'h0;
 Ie7d8d3754dc7cc7ac9fc8ebcbd3bf82a <= 'h0;
 I903284ce681f1526c56a4889306a65ec <= 'h0;
 I2e1e3933f8ec5db47edbec59fd1772b5 <= 'h0;
 Ieccf95256e095c0e79b8ac959cea7655 <= 'h0;
 I5c9eba93bf9c01e161dd3bd508980acb <= 'h0;
 I8f66edb2bb1d6c6f228711fc27836a3d <= 'h0;
 I0be6fa3f4ae264a84a3b241edd706034 <= 'h0;
 I7fa9026688537d119b6997572564584d <= 'h0;
 I501a61dbbe9a6edfbf51d18b14d96f10 <= 'h0;
 I4fc839b634aaa2e0b5775984e0dbf6ae <= 'h0;
 I9a432f4a190d752c5e723107243daa1d <= 'h0;
 I23a1b8a01fbaa3122ef3d1efe362a3ff <= 'h0;
 I97a78caa8c75ef80934e8d013fee43a4 <= 'h0;
 I72d4a7275ddf3d5d41149fbc6e6cce23 <= 'h0;
 Iaf87541d81d0e3cefb78aecf3ae9c92f <= 'h0;
 I55ebb5c7ded985c8911629524e62aa16 <= 'h0;
 I19a49d3680e5786fad7060cbc4be4a16 <= 'h0;
 I60e4a3789fb3df162298306c815259b2 <= 'h0;
 I25054529bc0fe35bd08f6294a2d51f5e <= 'h0;
 I8a471bd6f3fd220a34d9cc870eaeafe4 <= 'h0;
 I12d2ea504991199ca905ca91925f2d26 <= 'h0;
 If93a23874096c597803aa347c0900cd2 <= 'h0;
 I5f3af0ef6d4722a508201707b6994fed <= 'h0;
 Ib88cf5d737b09afb18cbce8072be2ea0 <= 'h0;
 I626fef2cd9d071cb8c797471055cf245 <= 'h0;
 I723088e5c9b31e731220874d2f27f195 <= 'h0;
 Iacdb27c060a48b7ade76d256e858b314 <= 'h0;
 I3719da3863fb069e898484ce997c2f40 <= 'h0;
 I3dfcd0d247d56f8167bcbc6aea6e3504 <= 'h0;
 I477e8f9e2ac8c5d142856ec6787e28ac <= 'h0;
 I2865e7f35c36e2cd4a4e3435aa8c7c14 <= 'h0;
 I4d83852d202e9f1c49955b59d183cc07 <= 'h0;
 I7d5b2a7bca99f2164a7ba2cfe46b20e1 <= 'h0;
 I3c7c5071212ff5db857e3f84f6131391 <= 'h0;
 I6296deff598d27ebc1a06cb1316a3eb4 <= 'h0;
 Ie6acf5390a3487fca3f8e4b66a640da3 <= 'h0;
 I6a993db6733d3efe90511bbe7f4d5654 <= 'h0;
 I3ba62f936f0832ff2ebed33f862286ff <= 'h0;
 I0f8f8ce5dfbc020b547758c239f923c4 <= 'h0;
 Ife2ceb6bb50cdc7adb4a20e1851d54c5 <= 'h0;
 I361c911024ff757958306a38c4bf4465 <= 'h0;
 I8ca3c12dd3e04f05ca52ebd1ea32cfee <= 'h0;
 I56a419f6f3b841e7e5dbbbcc0e6af190 <= 'h0;
 I5ee41fe39af22ebe82e91a1dee0b7221 <= 'h0;
 I807e19c30c0328199d5ab2d64593d509 <= 'h0;
 Id4a5425f6a2a8a689eb1e5e25131fa0c <= 'h0;
 I2ba381005b1ffbcf163c40f2dd92d2f9 <= 'h0;
 I2a48609c13ebc0cc9a8551fdf244a2d8 <= 'h0;
 Ib0db88e9d645459a03e908dbbf6b5803 <= 'h0;
 I9170cf346273d705158f36c2a9e59961 <= 'h0;
 Iec7ceaf0d09a3629dbe42f8926383e83 <= 'h0;
 I9d738422a85fb3cd648444a039b96e9d <= 'h0;
 Iece0c68af7dff6bbe73e9e2d468585c2 <= 'h0;
 I66f0d7b1c32cba28b55806d443090f9f <= 'h0;
 I3d2bc0bd4abfa1286242b841ef4f04ba <= 'h0;
 If83620428cf14f11cbd5eb3584a0e877 <= 'h0;
 Ib9161bcd780dcb77507b4851bb21193d <= 'h0;
 I584c580e66ed2d89371a7a1a4fd59599 <= 'h0;
 Ie3ac6cf6fedf997b6839abbcee584fce <= 'h0;
 I3a67256306c29f917d28ff55be76d4bc <= 'h0;
 I8506a14aacf97d360aa4c10a91ef184f <= 'h0;
 I6751092e3a762e4f0ac88e02e8d145df <= 'h0;
 Iaf3e9f18da33e20e42838b4467d9741c <= 'h0;
 I83649a386aab66f1c0774263a77831c7 <= 'h0;
 I8ff4739a83ed374704f039515b99162f <= 'h0;
 I9851d75a6dcdb74212fd0146a9aa49f7 <= 'h0;
 I9653890e840ec994e81844c9a34b10ba <= 'h0;
 I1322f065e413aef275747decaa48d550 <= 'h0;
 Iad493aff89cf569ffcc57b8f204c11ad <= 'h0;
 I99928f669eb8b23feb022a8fb39ef5f6 <= 'h0;
 I98207474d16dc958a7e695a56a81b614 <= 'h0;
 I422a5ea4034e59d308907e5684f8ad8e <= 'h0;
 I2911a1c5c49beebcd2fe684678ab89ca <= 'h0;
 I0a3206015f8d35fafd10bd4709b95faf <= 'h0;
 I10d423113bbfd394aca2695798b2d4ad <= 'h0;
 I596999303fc894014a5ae6ba2f09f143 <= 'h0;
 I1e24b9c9e023b6f0b00cdeaa071366a2 <= 'h0;
 I6983ea7dcebc925bd95ee96457a2de66 <= 'h0;
 I3d0c2d0d76d54c59e1d282a37e0aeae8 <= 'h0;
 I6f6c9a635c0ad62e7687a666f98ca4d1 <= 'h0;
 I929ddfd7ec9bf7b7c2dd2378395a403a <= 'h0;
 I6fce04d1f8c9975afa3e6abb203b13db <= 'h0;
 I88d063cb6f169e9f1ae067641fc0d802 <= 'h0;
 I2adbad4296c06db0ef231d53e6516986 <= 'h0;
 I4b139847ca9cce5281ceb1d63a453d05 <= 'h0;
 If9c81e3f27ee171ff282cc7fe18947ed <= 'h0;
 I7648b4562836acb77aebba8b19dc62e8 <= 'h0;
 I9f2892cd4e16b8719b5ffcb4b051ac0f <= 'h0;
 I159acdea94fb6185fccd6310e9d1b071 <= 'h0;
 I7a19ff6c711f9ed53df05a4999041a70 <= 'h0;
 Ifa65fb0d14e454b62f138630d2f9f370 <= 'h0;
 I0f24875d6dcbc0c7c83602f50ee3a8f5 <= 'h0;
 Ic888c593409b429e20523b414861da69 <= 'h0;
 Ic10e70c69f2401950c31aeaaa1600ed5 <= 'h0;
 I3c6576aed9ae9c1a1e86afdc00082fc0 <= 'h0;
 If710661738ba49d8040a1aaa6c4a0dfe <= 'h0;
 Ic6e2dd06abadb6b0613d8be1d3e91da7 <= 'h0;
 I6e72837b363b91f0a1301ccc2c3a9e32 <= 'h0;
 Ieb48cc2ae37e2d9dd9144b587cce78da <= 'h0;
 I0c2ea6ea58ccc53502b8765d9ab08a56 <= 'h0;
 I2590acd159fd90fe367126ce432e39e8 <= 'h0;
end
else
begin
 I371284eed470112cb89e1d361a9d40f7 <= I0c1c52a843a5de4bb5e0eb6897ea37c4;
 If0fb2e90431d89d99912918f83036f4c <= Ice4c8b10e41f361db2bd4a7b8470b05e;
 I0ee915f21334d38c75f0207e3b052a69 <= I612d62c35e606e6e91220910fd8448f1;
 Icf5a9bd712d310ac17eb2354f884a237 <= I4f664d460f924a71ebd3cc05f0916521;
 I3222cf2f98878be3f453560ddb3dc43c <= I0e38bd43118f53204e169f324066b75c;
 I2dd9e89f2842e748c1574ad0e7f4dba9 <= I46878ad6c93d318bf7a959c78090bf66;
 I667adc16c92bec8f413a1a9bbfc41ce5 <= Ie2c597c226457d94ec76f1513d95aab2;
 Ie6aa50a44574542826b78fed7d77b76f <= I2c72e48d1e2274c662c18b729af96161;
 Ie97072fa52f483bbd89f019c21152cdf <= Id416e2e4f204401c79d97ae6ae1414ae;
 I47f153e1cecaa77f1e6e6f07c0220557 <= I8fa96c5580fd6050e2a8c5fcb77c9927;
 I1b9dcfaf144b48a64b990e5b020d4a02 <= Ia9569f758e6bc743aae3a2bb51d941ee;
 Ie32d4bd927d02e547850331db8028177 <= I00ae3aaf6b44b2f7fd9bbceafb9c4e22;
 I0988db7ca497541e372131a0b0e8075e <= Ibfea7f98ec3bbe5588eb75cbcef739d7;
 Id13b5577b8baa586fedd34d4aab9d9c5 <= Id9eff948ed9da8502308740b4ae17dbf;
 Iedd0e0f6ee682a131d4f14c4762ea0eb <= If9d08c27c57ed8293171486ad65ed95c;
 I875d7c55914414298f0fbec0b345c92e <= Iace1409bfc12437ef093b91d50c8175a;
 Ide64c9647c7898867e0d036e9ff95f6e <= I506d9cf5c368c130a8517f994e7f7a43;
 Ied6ccabb348ed7e20567011e027c86ad <= I0f3fb929c6ee46d33daeba7024107aff;
 Id030b072054c623c7aac5c571d052951 <= Id3ac7026a6f63b1dc8588f9bdfd50068;
 Ice55fb2e506accf518b4aa18298d017e <= I680caae24965f4516cbd8642d4d43b3b;
 I07a0167dcdfc76612e1b0da251337a7b <= I7b240e087870bef3e01b2de04cdbae13;
 I045e08f48738d395af2b79f25af73732 <= Ic2b7c4749006adaa1dfa0ca1c5d7a371;
 I7df57f27a880fe45f78c108f8faba963 <= I2abc1d3ddcecbdbdc971abb93be58744;
 I60204c1d3a96524bbbdf715f95f08fe4 <= I9fcc49fa3eb8ad62633822ff3ac5973a;
 Id5b9ae91dc900060caffff2520236f66 <= I6b938059b8a71491bf1718326233b688;
 I861fe9da6d004ce3998ab54a8c0d62af <= I5d98a20b0eef6a335b29f017cd3120df;
 I95caae0432aeadc0cbe279f9d6f9062b <= I69d5314c6ba43f6d015acf00c8a2a7be;
 Ic9c3b015d5830bf4834a435eba89caa5 <= I64ce8a8f7f046222c963820f37362021;
 I6e18dd1a579e09b80ac113fe85b483b4 <= I4e1c98665268d59e19c3068ff9efe9a8;
 I51c1c8e8df14396c5c77b5013531a84f <= I1399a46a42c2cc384efc8ca681b1b249;
 Ie8f75e8e020d43f6a357b5175047c254 <= I3e0d577c49e0fcba84112e3afab2edbe;
 Ie762d8aa151448cbaa0d005a3c01572a <= Ic266aa3f20103455635f801a0fe1056a;
 I293b32c043e20d6baab178319dd1e2f6 <= I285c0d0dbcb505b98bbf005805067396;
 I200aae813b664e02075eeefbc3b4450d <= Icba253e44f98c391c02e864856715f49;
 I006264bde45d8df078ef711c221ff387 <= Iaa4b6b01007d9836ae0092101c4065db;
 I9200a0071528b14dc52e92082768ca97 <= Ia2f4d61e666ea4e0d8085325cdaa7344;
 I55761decd7043b4dc82737b9d6ef6e7d <= I84ed644f3578e53744802bab05d17011;
 I4f51d114002bdfd69a31f95c2fa5234c <= I5fbdad2d56ab8f5435a712b512190645;
 I796cb71b28957405c10015a2ab7124c6 <= I670a7cf3b4948b0d31c871ba641af4c1;
 Ic85bacce5db48b4dd3f626749f6effa8 <= I227702af9307eb6600ed78a648bb71e9;
 I2a508066cf0e07bbe8a91f276fbb3078 <= If0c4078bb97b3a246a91be4180ee7af9;
 I85913ae95fcd63de45030d583846b1d6 <= I913f1af34aaf3d51d3c60489979a81d5;
 I971cff06a60916ea3e136b397d4c620b <= I22e712371781d71cbb80680359ccd708;
 I2c363f7abf62c9026d0b0dfe5a51207a <= I5e9450b27761da0b895a4f6ace1ad171;
 Ia5043b0c8ee086c66e683eb115a75484 <= I0b1bc20ea62f64bae807d8ac1166139f;
 I6b7b63ea23c5b4f3c597f121284cd2da <= Idddfbcad405258a5434d8b94eb26654c;
 I3cf82abadcee2faa1849d0a9a45b051e <= I8beef0ea5356b2f46d7d5f16db49ebef;
 I8b42f5455dd8f6323d7a4e28c0eaa1a9 <= I499586880161ca66628afed78e7e495d;
 I608597017b046d92b77226999df90600 <= Ie909ad4a9ba2fde8fd6451e7eda2088d;
 Ia39b908f8d6b63777376ca560cd0cc8d <= Iee75fb439b2200aba94b03fd69cd7adc;
 I87ad38ab473927df7c0bd69c6b4b4c5e <= Id8a8555f4bf9003a0ac0dcafaa67e68d;
 I8e70752f74ecdbe95a7b33ca264d4589 <= I10065fe206e6700159260af61afa61c2;
 I6e768e27a3f1804919e3f83c050e19ba <= Ia41593b7790fde4ae4dd986dd583286f;
 I2285f424ef2b8b2041267c1652155ad0 <= I44490a711aece8f1a24c080cd0f37607;
 Ibc5b97632aab1e763ac51f8d18edc792 <= Ic35377a5686c5a6edace93b58129cbdd;
 Ic4a0165bd71d9e586fdc66c824e45224 <= Iccd1e1793be28ddad794782e2700a4d0;
 I40de7aeac837276e7b3f0c4b29ce5eca <= Id112833f079dcf6e092d48cd13120d47;
 I024a746142e5ff074724f92af62f3bd3 <= Ia550c5040df02dc8a8735562e71ddf6f;
 I1e54f934fa92e681472d03199991f0b2 <= Ibcaed8bfefd254ded778d760cd533b81;
 I8cabd17b81e99a86fc8704aaaae629a3 <= I19c7906957daf8e2a04b013e95db9c6e;
 I54c1bf986182c83540d950762048a5e3 <= I4bbddbcd811dc6936fd20d18559e3aac;
 Ia5fbeb5be349b8088a749e25a9e6e416 <= Idaf09a27ce68e8877da2d4c48be4c8ca;
 I987b220a4729d14e9fc97b57867436e4 <= I82ad270d36061ef06232de9b92742dfd;
 I7f1d9309d3053256134130574b970425 <= Ieb5d1ef84057ceba02d9db624be39285;
 I9fd9d5a2a3a34b532bad740b16ce66fb <= I7ebd34e6a95c3589b44cc0941f54bfa9;
 I66a648a9f6b10b1d580e72b36a1ed9e7 <= I46432f8bb8f39efef70554ea0e8573de;
 Ia08c041d1aacfbbd1f8d7980923b9b05 <= I1fb7b6a528ec8d5871cb15a490bbfda2;
 I6805a2f26b1e51f7ac0087e6829b3c5c <= I25d429f4a9f397a0d0ca515241b3c1b5;
 Icc11f9d183454b33624bd411710342a0 <= I3ca008900582aea13c5cf09b6c3af78e;
 I18f145bedd3864fcebd983f9533a5877 <= Id9a5e1c4a044b3006d620dd52e2e8ddc;
 Ifa25d4c9ccc3efd1af4e711d3c32e9c5 <= I63f34eddeedc5ded8721b40546c758c3;
 I5bbf8f01c5ddaa02516dde3867ec3d78 <= I8ec5f00523507f51358081e52a5bc55c;
 I3f8fe2d052a6df20dfaac6f88d4fff8a <= Ib77465ae19c99c6e2c39e2ab6438730d;
 I9fbf9bcb6022bb550bc2dbd52f20d05f <= I025a54040366d4505896c1179d580dc1;
 Iacd71ce5854c85450463a0a45ebc6a2d <= I0ac7e4f7f0e68450455e4a3d3ed57c56;
 Id7c1a8f42cc90b7846105cd103b07228 <= If6f5c61447dbeeaef688c670c9802649;
 Ic6d94b59cd6f4c7765463694c9fbae3c <= I968168f5cd481033283f24425f7862b9;
 I11a9409c814372a31d771888692ae955 <= Ie364b2799febe180ea9c2361279bcdc3;
 I760f9ff7bc594c98e71080485cc1a082 <= I76cc2a7d1f750a49780fe7e7f1651d5e;
 Idb9be12ba6807752b0c36f4cc18843cb <= I2e3ac4cb975151fcb26d716ef80a24f9;
 I192119ad6ad1396dd6fd1fab6e4c4cca <= I6da8878ff3f8680907597ba4ab49e7e4;
 Ib4c62a865f79eaa2aa5fbd12860f2e80 <= I28db3b4aa4f26a48ef6a28956536d15a;
 I5fb195f29a4e02620d2cca6e7f2a8fa0 <= I7b95e7f8f8f6d01ad095fdfbe36e7f6d;
 I41b4d1d3d5ae22c8fe4f1e0fe20ccac7 <= Ieb56b02269e16c20b5f626afc1b97c98;
 Ib2afa3be272607c236cbd5410a88e8c2 <= I486565b0e63446c0b122a62bac6644da;
 I43587e6827dc7dc1ef38d552f6a73ca4 <= Ibd4082b5df0c5bca554397e77fbf589e;
 Ic27ed0f98cad254a72ade8253ccc01d2 <= I6361b4f6c6266288a5f53dfbf0e514cc;
 I5860a511728dad8112a9246843f0fdab <= I0590fa4c4cb5194e038b57fd416210b9;
 I6f83f4d8681a17b7e700a38a78917822 <= If8409ca3930cc882752b4efe399aa107;
 Ic902ce884c81efed3160715af43eb19b <= I509f64436f6d698c58fa255372adf7e7;
 I8297012f23a474aa863c56e6ab9f77f4 <= Ib6319f6f8e74409bd60d624b07fc75d2;
 I703fa28fdfb32f8e7fe5062a3332ff6a <= I344f88b13d6f536724dd33ed2d9fa07a;
 I4d60a4630a93dbf6460fc525f16fb69b <= Ia9c1251bf7d48ef32d67ee176ca55e07;
 If6a1f518420fbc246e2524469689a5e7 <= I8a885ced1613614d0bc3e1d2ce31cd34;
 I48c55cdc6c1e3bb5e36a5451cb43c5a9 <= I084e8923b177a76c4fbed301ae5f905f;
 I147accfb14f15341869779b74c8cadb6 <= I58d2c7aa1ec77bc041b6b1e2e4ad8277;
 I0d302535ee6928ed74d7b456efaf01e6 <= I9be477a653c8d0bd98ea404fa8876dd5;
 I0039a78cbf75de3d875c319e3bc08d22 <= Ifefb2b21271a5578ec1e1d9ddae2047c;
 I7a43154a62ef625844cda08b1dfc9c79 <= I708bb50785dd2710e712438dcfec5eb1;
 I8e05a477fab7c0c6f70c681626640b93 <= I12e20bdca30dd5a4695333353faaafe1;
 I51393ac63dc5f8c0898ffa6dd59ee183 <= I37da1f9f97e273359be9e4912f8a8ee7;
 Ib4f7dd6e43c7a291d753f96b1aac8ce6 <= I0df8e26f5e3a60744a02e8b50cff23a5;
 Ibf76adf5511e851727200f4fd60bf34b <= I0f005326cad2001188a9fc4b919bd19a;
 Id90de24703e5b15356a8ab3862612957 <= I1b7f0cb10a2a1c63083aa2e5d5fe84d8;
 I2b42badcbe3d18d033edbd6d4663fac6 <= I43240748b90a2f1b2738d7773256f36c;
 I72450aa2c2f2f501a5465f008e95ba4f <= I9d301fb4da56021d4bf0df8dd2719eb4;
 Ib802f2c9c1265a47e5acfc419034488d <= I50188fbeeabb5bbc1549229769cc58d3;
 Idb28449172f54add7ac6fd1287543a5b <= I85af941bfb4adc588579de64e51887bb;
 I6b33174bb2786da0ba9ba988a96aa5bf <= I6baa38fdfb9b81d807b09ca3b7cd5d32;
 Ib68892cce1de9f46fb391a7ee8a01afb <= Ica83cfc4696601a6936e577389a395cc;
 Ia0e39ef7db11ff2f95f50e6a912e945e <= I9ae9897faacb46733dcec0b985a590ce;
 I1f3153881fc6a7fc767a33253f80e06f <= Ibcf6f538d26631634b6ceafdd3ee991f;
 I994e4d13d16c12025cb60205b8f7559f <= Ia2d7c7007306e7b2ca65518fcc005588;
 I3e4b2dbb8f44350c5cff7430502401b7 <= I5db8abcf5c9f55ffbe360502c0acf592;
 Id1e6e9ac8ddad3aedd347aee9f615d9f <= Iebf161a4f32971bd911356670349e894;
 I5a6da3732e0f265ad95269f5a629c1e8 <= Iba78cb5ab1da071088bf8f924095d1dd;
 If8773fa380ec5c1199794d4128d443f1 <= Ib8bc0d119e76d93a801d9749ff205d30;
 I63283e5286a737d3ba1f99ae29902bb9 <= I7d760437e7830701c90db6653febff5a;
 Iedcc3a589dba858f1193b1be582db24b <= Ie7d3e4264ef52d194bcd054dc421e97e;
 I8a87d3adcb2989738d70db84c3b97a3a <= I2271582af0c776dadff851456aa6e4a7;
 I267e058f7db05744d80df6b52be83475 <= I851e3c75bf75803e1d745053721aa9ad;
 I5e121581d8a5f81fc84da2fa982d8fd6 <= Ifa32facd628d97fa55482c63464bbeed;
 I51f875fbf103d8b8093d73279f127843 <= I37a83fa1dac26d4614760db718790dfb;
 Ifcbf9c1d4d6f111f06212e58764d29ea <= Icdfa771d45c36fef80efda13b0481130;
 Ie0e816b57f511fc0479210deebbd9fc1 <= Ic72a44c59c204b5d5b77523429df133b;
 Ia7673dc1d477d486371935040ff7dce9 <= I1395b926b6d89fdfe41444e3a94d0d10;
 I7df5c4ad52bf35d254a4a14771a28fe7 <= I8393828bf7f4ce64ef97785fcd0d65fb;
 I9ae2d00bf699c7f12c3f5d78ad2c405c <= I2f6dc9f6f5d1316b9426bbe277b82427;
 Icb740a93e2adc0a9f18ac25d0c5d018c <= I60098787140a26167a69e135e08c6e8b;
 Ia9691e7c587528f3ca0d85d842225da4 <= Ice5b808b49ac5331f4fd6f36e74f0897;
 Iab732884bb2d4b1781e31c7a1c109000 <= I3480a29289d8eca6cbf762b798ec68fc;
 I67d8e4c822cc57b150a76dbb3478b5b5 <= Ie8718369d950a31dd1e9b307ce68984c;
 I3bb2f03bf7d2f7480187062b45c6fdd9 <= I954ad53f646754aa0c8db5073aff65fe;
 I8e57236f80078ae72706aa8102e1bf53 <= I8f9194a8b73a5008a74dfe09429e455b;
 I1732bcc59b7bad3d08b232d099fdefdc <= I9b0851ae1b88864bd086003066137b86;
 I4b568309171ac557250c2ec600b9d7b0 <= Ia8d552e62e3c642796936c2c4188f8a4;
 I886251a3307e5fe20788c8e947f4ef37 <= Idaffd115023b38f3f7e7cafe8e2cedb8;
 Ic0d064e8436ad001f7e9d97e800e5636 <= Id6ff758a9c646a75ea986fe323b91966;
 I9f2ba5b0600c5eb81cef40d0822d0aea <= Iabbe6a5d643c1d8c3f7e2c8ddb41f8f2;
 I2aaf6ff0daa3d3e26b197e6895cabf3c <= Id4b54da5ca05664d454c620a63622da2;
 I2e8c68a51f1f1f4e413897791a6823a0 <= I0e4e792c6af3f2575e3e36eed213e7bb;
 I1a318a04ba3cf92f4ba0dc132a564040 <= I2c7afb36c88b388e24d0edf20acf3bf5;
 Id32b88b33bfbcf79ff0a10d447f69619 <= Ibb053ae1486e202396d69ec80ceb37b5;
 Ia41215dbdcd4b27a8ab41f48d40d644a <= I88a88c8c4b3a9af4f49565aac9e5f248;
 I53c239961c5745db892194a0a62b5d57 <= I359e996afe4b35d29d9180b990a27fcd;
 I0ffed4dfc4e97bb477647e5eab3a18f3 <= I899a8e3a18bc3f9e4f3a5af73fa61dcb;
 I46fcaa5311cc831199bb4a5a3dba797e <= Ic124969a8cfb359b1ccc12c38b92f031;
 I69b693e03eccfe9a889894988c0c9a53 <= Ibd06fe0881c395a5e679d87fb9ffdef4;
 Id0ca109680ce0cb6603139baeebac59f <= I8d0c94e6e41f653eeefb5b911e56e229;
 I7bcf3409fb1f7bf880f945db8f2eb6c2 <= I06d6e9bf2bf5fe1d0d06a7a7bf9aef4a;
 I873254d95f4a9976acf9210228365521 <= I3df5795d906a0f00bf42bf6e3ea2da66;
 I2a437c10a562e8e7f4cef30bbfde2fd3 <= Idf0aba59612a66e3e74e0a90e1f24024;
 I50e26d2184d04613f297357308e7c91e <= I4ebe1cce938e487efd6289f437e5dc5a;
 I8b14ff6b303ae081ae414ca7a00da3eb <= Ia2818dffb7609ae601acc9bad920308c;
 Ibf3a99967d7cbab53676fed78da28eb8 <= I26a3e6a339b41ad00866844786681513;
 Ifb6cf60f578b5a5dd0c27da72408cbce <= I76b2e256804d1913c453dc19742869fb;
 I000bdba9ccdb068a02fd37d2991675b6 <= I2ff4e3eb141f0d9f284bab6b5c9eb9bc;
 I5110f5370812f6d0319c0f42a6638b5b <= Ife7243ad867ecc4e311906fc4ede4451;
 Ic36cb86884806afb677ac8fb42aead36 <= If65d250d229376f2091caa5d0eed8b8c;
 Ie4dba51278ebf8a9358c2019383fbaf8 <= Iab0e973383f884115980f16a6261ebfb;
 I96373fc8bdf40551ef8206b4ba38cd98 <= I2c4e82e4c7fe3917596e9dfe8f01f865;
 I7b8a50810f6a4c27a23c82330707c4b6 <= Ie17470e1d818de84c8e5e0269c5a18c3;
 Id84a4cc9f82244c2357edc537824eb30 <= I25a3a01cc23b7303e828c5a76d108335;
 I8866b1e80ead799943d3ad273ee0c97e <= I393c613e2dc208cf7724920ccf7da4a2;
 I33d92c1bdacf71fa60865f1741288cdf <= I6dcc14bced84384b08b054ad1ed5d6ba;
 I834a4a93056d8777cd2d4996ae33122a <= I93713849034deecf3189479b9012f123;
 I51bc583f480542f3f95241643bb39eee <= Ia20663615bcd8de7a403e368c23aa942;
 I35539407bedb7d43642e952787216ce6 <= I2623b7a7673b4061c0cfdd92e0119112;
 Ifa78beaa6ae7a7a32f4886a14e4d1532 <= I37517b2fa41b7fa2d25a45058b8369d1;
 Iae691c305b2fd52617ef92705568a8b8 <= I613289d33f6a2742ef380880a6e4fe0b;
 Ie87c6bd3452b53ef57df5f420f351434 <= I79d675be55634575c1ca36153e9b3637;
 I03106ddaebe00bc59e1611573835f727 <= I5a21a18c1e1992154869c922fa691c74;
 I8b947b6c3139066fbd5873d5b818183e <= If8be80c27161a6257e0f1d41359727e0;
 Ibb1c668cb8ad3eb49b9bff842d118aa7 <= I7991f753713b02ebd49178ca1ca2f1cc;
 I4c3bda40c1fe5dbacee1829e0d60bcab <= I040f9f3dc40e2bcc958191055ca6b6d2;
 I405504d762cd698722b183721df7243f <= I70a8f1f9966c63b414a3bb68e5e3972c;
 Iae9c6245aa98b5758df6d57f8c33ab31 <= Id8f36cdae93ca8a388aff8fb4806f4a3;
 I35f897e994d6fb9ae452bee5b423c4e9 <= I906be6a8bc43d22dd04b47c2bba5c2f9;
 I413a7fe2255064627ed283d35d910de4 <= Id4df0a1c44ea75f32970739cb4c5a2cc;
 Ic930f61e087bf2477712e8fef9c413d3 <= I971cb87b4023114252557346c9a07d0e;
 I61ce1d41fa5221c01f7e9571965eb3fe <= I6e1912c5b6a09ff090f2d49d51002030;
 Ic70b0be144931713bc160b7b4d8038e2 <= Ia276ca65e85b9ccd4a9553b970b418a9;
 Ic854870518bb942314f6269c6833ff5a <= Ia0b083b9bf3175a9961f79464d1b6bde;
 Ifdbf3e9abf7bff7ce4c689bb7e1226f4 <= I6aea13b6ec3703c9c919731b7c43e44f;
 I4576ad4e2708a5635d93b304f1f10677 <= Ieb8b3cb38d28c4357bbd35d485f66dfe;
 Ibe54160f877c63dfaace0fc2c41ff11e <= I25fcdd6fea9bc9d728e5b6dc28cabee4;
 I04e75fe6916169cea741152b9fc6600b <= I0ef97b8205f4a544cc31d1ab9fd62d90;
 I60fc524227900d3fcb19263336db4383 <= I157f4891b58262db67a57781e6789205;
 I11555ad63e8caa81cb02dd9264668a3d <= I0306b43f29eb07e97472616ba7516f54;
 Ie9feb0382e321c4cc1602c4fab33f939 <= Id8c72b2670ca8001c69b60551519f4b8;
 I21a1b05b4e659507fc3ff2077e7d2e8d <= If32e24d0be817c10df587ed0aac48af2;
 I5af0b1d227ed007db9cd98d8a93b89a6 <= I6c17cb40f5ab67595f89afc0aa3e570d;
 If9bdb9270926fe47e645cea702bf7775 <= I2789fbaed627ab6bea83080a0634f73d;
 Ie6694b28f83262c5051dd00e336eb8da <= Id4415bf69046a95359a7f23a0ec3d5a3;
 I500e2c4d34270abc5a6f51cec578a7b5 <= I25862ee3c8452b8f0d3187132477b77f;
 I4c4c87637fc7973a58e933ffa76e611e <= I5e8114931cbd9da66eec0a9e96b647b3;
 Id7d81b33ad4bd7ae9df6a69b8e1e3351 <= I01a946c09a7ce0b62c7ba805e301de52;
 I9eae9bcc567e9c051d268bd446b238ec <= Ice805f2d2607178baf73b8c8bdd1b725;
 I614d496a5262a7f6ebd9a2d078ad30ac <= I77767e8e8a46c270774c64d18eebca4c;
 Ifdde7e51b6c92f13208685e0dc05c95f <= Iac7d03545a18a22c01e97d9f8ca93e40;
 I0ce07744582a47bf9cfcbdb2776a04c3 <= I1a60f16daa4667129838097d94c932b2;
 I4b0ae6a7608a5ba8b1d66f7dac61bd11 <= I8f08550281859dc884c13197e046ef10;
 I6c2a048243ceddc9e31b7a37f74eeac1 <= I23978d82bd6e911f5366f97765be24aa;
 I461cf1d25b347dd378a48f0dd2f5c5ae <= Ib26450dc355c3ca34ba704abe7350e2d;
 If32b0bc17ee8e3a95335b09550f05167 <= I29c302625d14d028e34ae65f37961e3a;
 I2f751a32b067b688a98c0d98a8461265 <= Iede527989cec0a93d78423b7df14d707;
 Ib8528ee13f669ca3b7d0fddcc4fe697c <= Ic0b1d8a6c00df4a35e285accfd1d149b;
 Ic0698d2eab5cdc70666a51ac0962e5f4 <= Ic82e6892a22a0fd064bdfbe31cc171f3;
 I2ff4fa27b4aef5cca03eff8bb129a9eb <= Icd96d324832586b90e3d89709934fc9a;
 I7770f02fbe5d3c1c49b9d5a3ffe4cd24 <= I07aea291890873ea17e211143a7a8291;
 Ib731ae113881b22a9abea15970d8c906 <= I424af84f8e7d7f4c85fe9e4632d0a5b1;
 Iaef6a7213e546e24b635fd39c69b22a1 <= Ied903684ae1a9f6b1d39d3714b6db7d1;
 I5f2f0073edbf2de118fb329b9d2f6d2c <= I07e0123a7a61773a58a82d037140d1bc;
 Idf85836a87828a65b1a189608df72380 <= Ideeabf83d0b70f18efb7a46d88efc352;
 Ib3f304bc897f97659a51764e156f4002 <= I148d4ff69853a123a3c5a306e978d9a2;
 I02c642372452e4dc5069ceb96098ff71 <= If578b689c5609b11df900bf92d0a388a;
 Ie6a18db9c01142eb719b8426919a114d <= Ibc5a4c442eab539e5bb136a83112191f;
 Ia96c18f8eef3c498f310b2aace71b9cd <= Ia19a1d1736d5feb515750e680b83db4d;
 I94c6e4bc6b9ec661a6d76814aafa1e74 <= I98f9daa53631a03ce5f4d21fa499a734;
 I3c2369669172ef6a4f0a1b36916e4a34 <= I3a1a9a79b0dd6856b5d6ef8eda18c564;
 If22f0f17b0156ee153508c5e4c9742ff <= I9268175b692637227825c86f87dad083;
 Ife58da9674cbcfa416675f629c158399 <= I1571e04768855319692febc19c86f630;
 Iaefac912d485b61e57075ddb0212fc55 <= I382b613b4744799d708ecb0c361c7293;
 I4b044f5c58a7d4eab6a1d2735e997f44 <= I736ed9a09ea1b83b13fc3b53ded0c560;
 I805cf823cf1cc902fe63131647d582c5 <= I0e2430406a0c161380cfd60e7bbfa542;
 I468c07efbe31fa2f18ae967a769e5db0 <= Icfce7d26af22431c30d34d5738109a18;
 I68941b5c1b03152c7425aa0a1e347385 <= I070f6f095b8a43ed92048d9fcd6625b2;
 Iee2c7d458d2673fe0cd58bcae0eca7de <= I7b5d1412081b2bad3b5dd0cffe78238f;
 I49597f093b8baac9c769fce82f7ad0d3 <= I04e76b2c5bf274bc2d8b9862c3690980;
 I2f80f409a3c59f56aa230c393d6c4297 <= I7fdb420f639b22294c896a20c8036f02;
 I87fcfc6fe1957f42e271128cfa0be7e0 <= I7a40ef6e10e3406e1d8c57ae53c6c3a1;
 I37b6525d09e5cd2be4f64b64d380cf06 <= I2e3fbfe6dd237424289f6f4d00ad486e;
 Ib915a0bb2acae5abe82646277a50f211 <= I2cef2ca61302b60079b80fd9f252c56c;
 If7d1635e4aceeaeb897a2b9d03caaac6 <= Ib44222bf07803a788687a877f1491ef1;
 Ib8ef3c757de68cd0afc90a6786286248 <= Id5fbe2f0dbe2a2d864202212c5db88cc;
 I627418190ef1e1115d0346d2db6134ba <= I6f4cc724a3e77e3b282e08a162448b75;
 Id59e1e3a73e7db64fd4808fed9e3e173 <= I573fcd75e769729647bc1c5fc8e54852;
 Iad4c43fc6e3ea0cddeb3da00b8faab4f <= I806e05d43c46bf4f67ccf2f1afa2911e;
 I097da986a541504f1f641404c1749e43 <= Ia2f45ae7f344cf3de7a61fcc35ae4651;
 If307175952944fcf9053a4d0eed964c9 <= I3debb601b68a3cd58ecdaa7d78e66c7f;
 Ib834d61619c282eb6994727f4b1fe2dd <= I9bc3698d4111848c8ff7f5082b4e6f3f;
 I9c6851db428c373c2fd723c1a374795a <= I4f5449753716964b3600bbcbd44902f0;
 Ib815852a6d56c5ea21f7a23acb120f3b <= I39de7cf13d732f3d5c89eaa718407a97;
 If80d97d0c5785dd6a0cd9fd3c0a6f870 <= I1936f1a842424a3fdc777207a05433c7;
 Ifdff70e8ea00c64f13abd0d6da5bc11e <= I2b5d24b895e1386c5acec6ec51af70ee;
 I64fc41bf20b9f82b2bb86fc9f2438e81 <= I9cdec4376c54fd0d5892b20f7f3944e5;
 I303191eabaa2211774eb1341a7ce1d32 <= Ic3dc6389680526e4e9f3db1a31c4e954;
 Ief8d6b623591a56818c091c5f08e9bcb <= I6de265c429ab7ef182f2ed2b52f413b3;
 I4fa399fc2e70ae442ef421db22b5ea9c <= I17dd943cac50d93f041a310edf916616;
 I4580e224188f11052c47c9d7d81178ac <= I2a2db61ae5f793391b0388d1139c1003;
 I3c484edf6cf740303824b22ad09ecdf1 <= I3a4a24d886c2c06e283081c1b0079aff;
 Ic22fe13fadb6b0abb614918dd785552d <= I1ae5bf5c035790ca6279076719f7d218;
 I015c6af005c8eb5a6ccdf97fd0073bbd <= Ic98fdc1a35fc3c698dd9c5bfe2fdd1ac;
 Iee7fd00e1644e71903c0ca268ba813ec <= I0b771b927e8acb823e30239c89aafe9f;
 Ic9143d7200fec6ef38e6cde1fc13d859 <= Ic3caaaecbbca186ebf9cc35e554ff62e;
 I974755cb3f16a1db503e4d6658d1f4bd <= I33fc4ecd929152c59d62af65ecb38414;
 Ie7d8d3754dc7cc7ac9fc8ebcbd3bf82a <= I09a3008676f21e58545563dff1cc9328;
 I903284ce681f1526c56a4889306a65ec <= I566a0851428acd33e432b33fe3c42b4c;
 I2e1e3933f8ec5db47edbec59fd1772b5 <= I96884d5c0babd2437ec14429856c0414;
 Ieccf95256e095c0e79b8ac959cea7655 <= I6a3539539860b98d7a310f63314a2932;
 I5c9eba93bf9c01e161dd3bd508980acb <= Ice31c844af4b8c3b966b778cca601527;
 I8f66edb2bb1d6c6f228711fc27836a3d <= I8eec3d66ef763226b960a24192aafe27;
 I0be6fa3f4ae264a84a3b241edd706034 <= I093a0ecd0a1aaea8a97d08d54cd37fec;
 I7fa9026688537d119b6997572564584d <= I3b2708fccba619958a392242efbbeea7;
 I501a61dbbe9a6edfbf51d18b14d96f10 <= I543deb703bb9eb808f4381f543e408de;
 I4fc839b634aaa2e0b5775984e0dbf6ae <= I0e0c7e753509c664971fd12be9183537;
 I9a432f4a190d752c5e723107243daa1d <= I68577e7dec24946ec0745c5d4255795f;
 I23a1b8a01fbaa3122ef3d1efe362a3ff <= If53e38b5b6031a7e927a65f90acf5120;
 I97a78caa8c75ef80934e8d013fee43a4 <= I372a38a8675f65c5257b645fb5d809af;
 I72d4a7275ddf3d5d41149fbc6e6cce23 <= I0d37309bb37b707e10a4e12425157fe3;
 Iaf87541d81d0e3cefb78aecf3ae9c92f <= I5935a4ee604a8c6259d88bd4b679babf;
 I55ebb5c7ded985c8911629524e62aa16 <= If4ed201fbbaa5ce9bfd05d65d79458d0;
 I19a49d3680e5786fad7060cbc4be4a16 <= I9b11c7aa2d35ee4589dec055ab0df2ca;
 I60e4a3789fb3df162298306c815259b2 <= I45a6d3691aef6c693ae6ee25c25a4b24;
 I25054529bc0fe35bd08f6294a2d51f5e <= Ia15364dea1e0f0243204b4bc4c9b8bb9;
 I8a471bd6f3fd220a34d9cc870eaeafe4 <= I2f31acde416c079c48ce54697eac5e60;
 I12d2ea504991199ca905ca91925f2d26 <= Idab577631403b170aa07d02c7d455315;
 If93a23874096c597803aa347c0900cd2 <= I36b79e4befc1673140076d2f9cbc9d82;
 I5f3af0ef6d4722a508201707b6994fed <= I9f263275a24efe9297aa995282c48360;
 Ib88cf5d737b09afb18cbce8072be2ea0 <= I7915e8a9a775ea1bc1bf7fe71648303d;
 I626fef2cd9d071cb8c797471055cf245 <= I4a7ac8c9709967341ededa935aa65581;
 I723088e5c9b31e731220874d2f27f195 <= Ibd7437a655d4985728ce070004e3b419;
 Iacdb27c060a48b7ade76d256e858b314 <= I8a834fd9d1425a79f7ff0713777fcdcc;
 I3719da3863fb069e898484ce997c2f40 <= Ia60cc135f03b89516e61d52335e69674;
 I3dfcd0d247d56f8167bcbc6aea6e3504 <= Ia1b1f012b02265afed03cb146e88f2a0;
 I477e8f9e2ac8c5d142856ec6787e28ac <= I6095ee8675c10be082abccd7cef7ceeb;
 I2865e7f35c36e2cd4a4e3435aa8c7c14 <= I2be07fc5652209f0e8eda31090dbb162;
 I4d83852d202e9f1c49955b59d183cc07 <= Ic60fc4bb6e7ccb8bee260e5b982bc5a1;
 I7d5b2a7bca99f2164a7ba2cfe46b20e1 <= I217d1876f768c7dd3eed096e2de59dfd;
 I3c7c5071212ff5db857e3f84f6131391 <= Ibb297f22ba2e0d4786042f7503ff3f61;
 I6296deff598d27ebc1a06cb1316a3eb4 <= I8d917a51d32729f4a5a98b5d3a40f947;
 Ie6acf5390a3487fca3f8e4b66a640da3 <= I08213a1a86aa27e3d3ed2d294d972ea7;
 I6a993db6733d3efe90511bbe7f4d5654 <= I271dfdeef4359fa9b2ebf80ca950a08e;
 I3ba62f936f0832ff2ebed33f862286ff <= Iff44a32b2e9a1a65d820b0839313015e;
 I0f8f8ce5dfbc020b547758c239f923c4 <= I2882587956babd713eb3a53af6afe389;
 Ife2ceb6bb50cdc7adb4a20e1851d54c5 <= I4f1ca888cae3ee3efeefafcfb12e16b3;
 I361c911024ff757958306a38c4bf4465 <= Icff2aa823d2f0e9421f3fbce6d21f510;
 I8ca3c12dd3e04f05ca52ebd1ea32cfee <= I2cd19bf0afc4563ea24619849ab7d8b7;
 I56a419f6f3b841e7e5dbbbcc0e6af190 <= I80cae65874911e05bc77db3e5fe0fcd2;
 I5ee41fe39af22ebe82e91a1dee0b7221 <= I18c43491892bd258dfd07aa0263c5479;
 I807e19c30c0328199d5ab2d64593d509 <= If322bf2a59be9bf7b33a49a6baf72ed7;
 Id4a5425f6a2a8a689eb1e5e25131fa0c <= I2bb21cbf03db27c0b9d814517033b56e;
 I2ba381005b1ffbcf163c40f2dd92d2f9 <= Ib408b39624c6576c228f32eed26ccf8b;
 I2a48609c13ebc0cc9a8551fdf244a2d8 <= Ib6dee36145f77a6f1364c218140266b4;
 Ib0db88e9d645459a03e908dbbf6b5803 <= Iafa25738d96fb115c78d8d295902c263;
 I9170cf346273d705158f36c2a9e59961 <= Ie7cb395e7ce65ca399d99a5e62a7efad;
 Iec7ceaf0d09a3629dbe42f8926383e83 <= I1bee0c6e3a24ee319d219799ce58f13e;
 I9d738422a85fb3cd648444a039b96e9d <= I7fcbf3d532ed0c810cdc1c5be536d263;
 Iece0c68af7dff6bbe73e9e2d468585c2 <= Ied7f9cbbcacc43332f1219e8bd0a07bb;
 I66f0d7b1c32cba28b55806d443090f9f <= I491888fefe23bb0bef60f293668491af;
 I3d2bc0bd4abfa1286242b841ef4f04ba <= I1b9368c7a0d236ed73a6783281144bca;
 If83620428cf14f11cbd5eb3584a0e877 <= I2adf1f34eb55f6f7e5f37b328b2bcf21;
 Ib9161bcd780dcb77507b4851bb21193d <= Iaa61cf5ca911de351708963438768cee;
 I584c580e66ed2d89371a7a1a4fd59599 <= Iacba64081faa56ef9190aa65fc89ae7f;
 Ie3ac6cf6fedf997b6839abbcee584fce <= I5d41596aeb3aeb4f07dbc0c995b5f4a3;
 I3a67256306c29f917d28ff55be76d4bc <= I1c01c903faacd546e44a6fd6564ef3bd;
 I8506a14aacf97d360aa4c10a91ef184f <= I3e3195b93f03e3c8c24655259f745374;
 I6751092e3a762e4f0ac88e02e8d145df <= Ie229e972daab0a41969c5cc066e52e61;
 Iaf3e9f18da33e20e42838b4467d9741c <= I5a646f85f9e6d52063b0c0e6f479f6f1;
 I83649a386aab66f1c0774263a77831c7 <= I01a50cb46ae1b229eda9094867090aae;
 I8ff4739a83ed374704f039515b99162f <= I68026b1eb748133551563bea029c3488;
 I9851d75a6dcdb74212fd0146a9aa49f7 <= I726047b0a4d45f8ad1f394301dbfb78d;
 I9653890e840ec994e81844c9a34b10ba <= I2cddfa0b89e0aececac2dd7d983beb26;
 I1322f065e413aef275747decaa48d550 <= Ic5e1dd806582ee08eb6d1048d6617b13;
 Iad493aff89cf569ffcc57b8f204c11ad <= I9040f68430c75ce7527990dd702b7feb;
 I99928f669eb8b23feb022a8fb39ef5f6 <= I40ebb4eb571f18c2fb810daab0d5770f;
 I98207474d16dc958a7e695a56a81b614 <= Ia4738ee511867aa46e0e92f3d86c4ccf;
 I422a5ea4034e59d308907e5684f8ad8e <= Ic10326eae7434399af6e611e31389963;
 I2911a1c5c49beebcd2fe684678ab89ca <= I8fafe7fe582d027b97dbf2cc58763096;
 I0a3206015f8d35fafd10bd4709b95faf <= I8a329168f83731c15dbedb1f1f966d78;
 I10d423113bbfd394aca2695798b2d4ad <= I603a5f82891f62b59f7890d631d0b6df;
 I596999303fc894014a5ae6ba2f09f143 <= I620517db078658289fcde4200f15ac06;
 I1e24b9c9e023b6f0b00cdeaa071366a2 <= I51271c02c6fd9cbda153c9b28aa099e3;
 I6983ea7dcebc925bd95ee96457a2de66 <= I8def31183d1a648a6a50245eeb6b57a1;
 I3d0c2d0d76d54c59e1d282a37e0aeae8 <= I0c3a1185a9fbb05c0dcec0d655068786;
 I6f6c9a635c0ad62e7687a666f98ca4d1 <= Icf0284aeb5d603e893733d2139a79ef3;
 I929ddfd7ec9bf7b7c2dd2378395a403a <= I3d0e6fa7f7edbd105fd8f7823722bcf0;
 I6fce04d1f8c9975afa3e6abb203b13db <= I55e28dff0ebd1007f4f00c512f1df1b7;
 I88d063cb6f169e9f1ae067641fc0d802 <= I2b33fef3c83dab2f2d254cb295264482;
 I2adbad4296c06db0ef231d53e6516986 <= I1689bfa3340ff4798ef7eb160714ede5;
 I4b139847ca9cce5281ceb1d63a453d05 <= I1b5deee5754dcc0762ca2691fd927056;
 If9c81e3f27ee171ff282cc7fe18947ed <= I1e63fce77120b91dc6195d2febce4d42;
 I7648b4562836acb77aebba8b19dc62e8 <= I1d3f5624cb6f217fac422833ed8b7195;
 I9f2892cd4e16b8719b5ffcb4b051ac0f <= I1fde6652c1fb298d84e88620edc9e91a;
 I159acdea94fb6185fccd6310e9d1b071 <= Iffd2d0fd17d604ddadcfc2dd9e46276a;
 I7a19ff6c711f9ed53df05a4999041a70 <= I8295b6fa92e241d4b689ad0e26f6a2db;
 Ifa65fb0d14e454b62f138630d2f9f370 <= I8573b3db0d36442c2f233d12586d82f5;
 I0f24875d6dcbc0c7c83602f50ee3a8f5 <= I5319144e65be1e69c9ef767bfecd4ea3;
 Ic888c593409b429e20523b414861da69 <= Ie7da9e9fdd626504cb2f00a3ec899718;
 Ic10e70c69f2401950c31aeaaa1600ed5 <= I8293d7dc145b31d28c05c02677760e9a;
 I3c6576aed9ae9c1a1e86afdc00082fc0 <= Ia372f6e388ed5cf8e9810c52d3749136;
 If710661738ba49d8040a1aaa6c4a0dfe <= Ibd959e3bf9ef7ee76ec2754a06926d9a;
 Ic6e2dd06abadb6b0613d8be1d3e91da7 <= I8f03815159c11486a4805e7f72c84a38;
 I6e72837b363b91f0a1301ccc2c3a9e32 <= I15e5e06b7dcf6616094faeb798a0fdc8;
 Ieb48cc2ae37e2d9dd9144b587cce78da <= If23f4bc5d45a3e7a22a9e8596b99c575;
 I0c2ea6ea58ccc53502b8765d9ab08a56 <= I70afe2bb83173aa96269271270d03f2e;
 I2590acd159fd90fe367126ce432e39e8 <=  start_d_flogtanh0x00000;
end
