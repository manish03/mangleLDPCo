parameter n_minus_m = 'd40;
parameter n_int = 'd208;
parameter m_int = 'd168;



parameter z_int = 'd4;



wire I6f1a75e774a70c6b59279764b820c455; 
assign I6f1a75e774a70c6b59279764b820c455 = 
        y_nr_in[1] ^ 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[14] ^ 
        y_nr_in[25] ^ 
0; 



wire I6cac6b878889968e94101cb5f36d695d; 
assign I6cac6b878889968e94101cb5f36d695d = 
        y_nr_in[37] ^ 
        y_nr_in[40] ^ 
        y_nr_in[44] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[0] = 
I6f1a75e774a70c6b59279764b820c455 ^ 
I6cac6b878889968e94101cb5f36d695d ^ 
0; 



wire I7a5dae8d8ca069078ba2d63900ac5b86; 
assign I7a5dae8d8ca069078ba2d63900ac5b86 = 
        y_nr_in[2] ^ 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[15] ^ 
        y_nr_in[26] ^ 
0; 



wire I02eeb7b4d4ec59ae0aeb59b87e7d9e77; 
assign I02eeb7b4d4ec59ae0aeb59b87e7d9e77 = 
        y_nr_in[38] ^ 
        y_nr_in[41] ^ 
        y_nr_in[45] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[1] = 
I7a5dae8d8ca069078ba2d63900ac5b86 ^ 
I02eeb7b4d4ec59ae0aeb59b87e7d9e77 ^ 
0; 



wire I0928decc55b7e882ab070edd079aaeba; 
assign I0928decc55b7e882ab070edd079aaeba = 
        y_nr_in[3] ^ 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[12] ^ 
        y_nr_in[27] ^ 
0; 



wire Ib688d0f14e5c3e856f7fa73809f0f2a4; 
assign Ib688d0f14e5c3e856f7fa73809f0f2a4 = 
        y_nr_in[39] ^ 
        y_nr_in[42] ^ 
        y_nr_in[46] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[2] = 
I0928decc55b7e882ab070edd079aaeba ^ 
Ib688d0f14e5c3e856f7fa73809f0f2a4 ^ 
0; 



wire I6f65c0d31734679921529495ea3772af; 
assign I6f65c0d31734679921529495ea3772af = 
        y_nr_in[0] ^ 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[13] ^ 
        y_nr_in[24] ^ 
0; 



wire I0186182b974c898821bd080775fca83b; 
assign I0186182b974c898821bd080775fca83b = 
        y_nr_in[36] ^ 
        y_nr_in[43] ^ 
        y_nr_in[47] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[3] = 
I6f65c0d31734679921529495ea3772af ^ 
I0186182b974c898821bd080775fca83b ^ 
0; 



wire I3e87075c14fd49a26c9e10b1cdd0daf6; 
assign I3e87075c14fd49a26c9e10b1cdd0daf6 = 
        y_nr_in[3] ^ 
        y_nr_in[14] ^ 
        y_nr_in[17] ^ 
        y_nr_in[21] ^ 
        y_nr_in[26] ^ 
0; 



wire Id7605657f7b356d38c15a612f29ca630; 
assign Id7605657f7b356d38c15a612f29ca630 = 
        y_nr_in[28] ^ 
        y_nr_in[32] ^ 
        y_nr_in[36] ^ 
        y_nr_in[44] ^ 
        y_nr_in[48] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[4] = 
I3e87075c14fd49a26c9e10b1cdd0daf6 ^ 
Id7605657f7b356d38c15a612f29ca630 ^ 
0; 



wire I3858b188811df9290d0ae4e1af7eebdb; 
assign I3858b188811df9290d0ae4e1af7eebdb = 
        y_nr_in[0] ^ 
        y_nr_in[15] ^ 
        y_nr_in[18] ^ 
        y_nr_in[22] ^ 
        y_nr_in[27] ^ 
0; 



wire I2a643f1ae9595a2834b7b4efb3fe1751; 
assign I2a643f1ae9595a2834b7b4efb3fe1751 = 
        y_nr_in[29] ^ 
        y_nr_in[33] ^ 
        y_nr_in[37] ^ 
        y_nr_in[45] ^ 
        y_nr_in[49] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[5] = 
I3858b188811df9290d0ae4e1af7eebdb ^ 
I2a643f1ae9595a2834b7b4efb3fe1751 ^ 
0; 



wire I57824975e3f21fc32f30355cc50b281c; 
assign I57824975e3f21fc32f30355cc50b281c = 
        y_nr_in[1] ^ 
        y_nr_in[12] ^ 
        y_nr_in[19] ^ 
        y_nr_in[23] ^ 
        y_nr_in[24] ^ 
0; 



wire I4b74027daab9b73a87ea34f841520c87; 
assign I4b74027daab9b73a87ea34f841520c87 = 
        y_nr_in[30] ^ 
        y_nr_in[34] ^ 
        y_nr_in[38] ^ 
        y_nr_in[46] ^ 
        y_nr_in[50] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[6] = 
I57824975e3f21fc32f30355cc50b281c ^ 
I4b74027daab9b73a87ea34f841520c87 ^ 
0; 



wire I27f049f03d2e955683a43486c1d9cc6a; 
assign I27f049f03d2e955683a43486c1d9cc6a = 
        y_nr_in[2] ^ 
        y_nr_in[13] ^ 
        y_nr_in[16] ^ 
        y_nr_in[20] ^ 
        y_nr_in[25] ^ 
0; 



wire I5b6a2a50df56add8a025dd2f2ea5efe3; 
assign I5b6a2a50df56add8a025dd2f2ea5efe3 = 
        y_nr_in[31] ^ 
        y_nr_in[35] ^ 
        y_nr_in[39] ^ 
        y_nr_in[47] ^ 
        y_nr_in[51] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[7] = 
I27f049f03d2e955683a43486c1d9cc6a ^ 
I5b6a2a50df56add8a025dd2f2ea5efe3 ^ 
0; 



wire Ia67c51a12204e65ba3bd8578ae7c9e23; 
assign Ia67c51a12204e65ba3bd8578ae7c9e23 = 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
        y_nr_in[12] ^ 
        y_nr_in[16] ^ 
        y_nr_in[32] ^ 
0; 



wire Ie2e4b274b6bc6fea073b4a39f318838d; 
assign Ie2e4b274b6bc6fea073b4a39f318838d = 
        y_nr_in[40] ^ 
        y_nr_in[48] ^ 
        y_nr_in[52] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[8] = 
Ia67c51a12204e65ba3bd8578ae7c9e23 ^ 
Ie2e4b274b6bc6fea073b4a39f318838d ^ 
0; 



wire I28f13c8d2c5c324a981ae667f99d1268; 
assign I28f13c8d2c5c324a981ae667f99d1268 = 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
        y_nr_in[13] ^ 
        y_nr_in[17] ^ 
        y_nr_in[33] ^ 
0; 



wire I82bc2997b68a0cdba7c9697aad8d67ea; 
assign I82bc2997b68a0cdba7c9697aad8d67ea = 
        y_nr_in[41] ^ 
        y_nr_in[49] ^ 
        y_nr_in[53] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[9] = 
I28f13c8d2c5c324a981ae667f99d1268 ^ 
I82bc2997b68a0cdba7c9697aad8d67ea ^ 
0; 



wire Iacce51ad287ecdd51e65b15b7c9f61ca; 
assign Iacce51ad287ecdd51e65b15b7c9f61ca = 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
        y_nr_in[14] ^ 
        y_nr_in[18] ^ 
        y_nr_in[34] ^ 
0; 



wire Ic9bb4be8798f9b593215b2287553daeb; 
assign Ic9bb4be8798f9b593215b2287553daeb = 
        y_nr_in[42] ^ 
        y_nr_in[50] ^ 
        y_nr_in[54] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[10] = 
Iacce51ad287ecdd51e65b15b7c9f61ca ^ 
Ic9bb4be8798f9b593215b2287553daeb ^ 
0; 



wire I4f47f7c1a721275e7adf311eda66444e; 
assign I4f47f7c1a721275e7adf311eda66444e = 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
        y_nr_in[15] ^ 
        y_nr_in[19] ^ 
        y_nr_in[35] ^ 
0; 



wire I73646f40cd547b9ca1769ee7a042b88a; 
assign I73646f40cd547b9ca1769ee7a042b88a = 
        y_nr_in[43] ^ 
        y_nr_in[51] ^ 
        y_nr_in[55] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[11] = 
I4f47f7c1a721275e7adf311eda66444e ^ 
I73646f40cd547b9ca1769ee7a042b88a ^ 
0; 



wire I1575f4a29affe00dcc863457fcebd435; 
assign I1575f4a29affe00dcc863457fcebd435 = 
        y_nr_in[4] ^ 
        y_nr_in[10] ^ 
        y_nr_in[18] ^ 
        y_nr_in[20] ^ 
        y_nr_in[25] ^ 
0; 



wire Id94abdd3f0fe21eba8b25a4aae15e1fb; 
assign Id94abdd3f0fe21eba8b25a4aae15e1fb = 
        y_nr_in[30] ^ 
        y_nr_in[34] ^ 
        y_nr_in[36] ^ 
        y_nr_in[40] ^ 
        y_nr_in[52] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[12] = 
I1575f4a29affe00dcc863457fcebd435 ^ 
Id94abdd3f0fe21eba8b25a4aae15e1fb ^ 
0; 



wire Ifde44d59cfcd9b6210df197b5568c133; 
assign Ifde44d59cfcd9b6210df197b5568c133 = 
        y_nr_in[5] ^ 
        y_nr_in[11] ^ 
        y_nr_in[19] ^ 
        y_nr_in[21] ^ 
        y_nr_in[26] ^ 
0; 



wire I082d600f71c54f7ab2658e3764206bbc; 
assign I082d600f71c54f7ab2658e3764206bbc = 
        y_nr_in[31] ^ 
        y_nr_in[35] ^ 
        y_nr_in[37] ^ 
        y_nr_in[41] ^ 
        y_nr_in[53] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[13] = 
Ifde44d59cfcd9b6210df197b5568c133 ^ 
I082d600f71c54f7ab2658e3764206bbc ^ 
0; 



wire If1618f3776387e59d5e95808a9f350a0; 
assign If1618f3776387e59d5e95808a9f350a0 = 
        y_nr_in[6] ^ 
        y_nr_in[8] ^ 
        y_nr_in[16] ^ 
        y_nr_in[22] ^ 
        y_nr_in[27] ^ 
0; 



wire Ic36348bc39d3601846b9fb1867b514e1; 
assign Ic36348bc39d3601846b9fb1867b514e1 = 
        y_nr_in[28] ^ 
        y_nr_in[32] ^ 
        y_nr_in[38] ^ 
        y_nr_in[42] ^ 
        y_nr_in[54] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[14] = 
If1618f3776387e59d5e95808a9f350a0 ^ 
Ic36348bc39d3601846b9fb1867b514e1 ^ 
0; 



wire I5d3f90fb97d3baa54c8e6e1a9c78592c; 
assign I5d3f90fb97d3baa54c8e6e1a9c78592c = 
        y_nr_in[7] ^ 
        y_nr_in[9] ^ 
        y_nr_in[17] ^ 
        y_nr_in[23] ^ 
        y_nr_in[24] ^ 
0; 



wire Ic33e43c8c227d597550b6b84cbc90ad9; 
assign Ic33e43c8c227d597550b6b84cbc90ad9 = 
        y_nr_in[29] ^ 
        y_nr_in[33] ^ 
        y_nr_in[39] ^ 
        y_nr_in[43] ^ 
        y_nr_in[55] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[15] = 
I5d3f90fb97d3baa54c8e6e1a9c78592c ^ 
Ic33e43c8c227d597550b6b84cbc90ad9 ^ 
0; 



wire If8a63370a226423e4a1fac7f5707ed24; 
assign If8a63370a226423e4a1fac7f5707ed24 = 
        y_nr_in[3] ^ 
        y_nr_in[6] ^ 
        y_nr_in[47] ^ 
        y_nr_in[56] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[16] = 
If8a63370a226423e4a1fac7f5707ed24 ^ 
0; 



wire I8bb7c789a604fbc4e6e0f18cc7ac7e8c; 
assign I8bb7c789a604fbc4e6e0f18cc7ac7e8c = 
        y_nr_in[0] ^ 
        y_nr_in[7] ^ 
        y_nr_in[44] ^ 
        y_nr_in[57] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[17] = 
I8bb7c789a604fbc4e6e0f18cc7ac7e8c ^ 
0; 



wire I411ca96a0fab2fc3567676c79c37db3b; 
assign I411ca96a0fab2fc3567676c79c37db3b = 
        y_nr_in[1] ^ 
        y_nr_in[4] ^ 
        y_nr_in[45] ^ 
        y_nr_in[58] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[18] = 
I411ca96a0fab2fc3567676c79c37db3b ^ 
0; 



wire Idcaabb5c30032343892ff44ed2c12149; 
assign Idcaabb5c30032343892ff44ed2c12149 = 
        y_nr_in[2] ^ 
        y_nr_in[5] ^ 
        y_nr_in[46] ^ 
        y_nr_in[59] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[19] = 
Idcaabb5c30032343892ff44ed2c12149 ^ 
0; 



wire Id0a7516377a8704a17006e040ac2c260; 
assign Id0a7516377a8704a17006e040ac2c260 = 
        y_nr_in[3] ^ 
        y_nr_in[5] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
        y_nr_in[47] ^ 
0; 



wire I509fda348d96588af57fac13ce87a464; 
assign I509fda348d96588af57fac13ce87a464 = 
        y_nr_in[60] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[20] = 
Id0a7516377a8704a17006e040ac2c260 ^ 
I509fda348d96588af57fac13ce87a464 ^ 
0; 



wire I7729a9afa2264d4707ecbc78b11ddc61; 
assign I7729a9afa2264d4707ecbc78b11ddc61 = 
        y_nr_in[0] ^ 
        y_nr_in[6] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
        y_nr_in[44] ^ 
0; 



wire Ie17136a034aa20fa1f2dc9c0134bf3be; 
assign Ie17136a034aa20fa1f2dc9c0134bf3be = 
        y_nr_in[61] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[21] = 
I7729a9afa2264d4707ecbc78b11ddc61 ^ 
Ie17136a034aa20fa1f2dc9c0134bf3be ^ 
0; 



wire Ic677b8f221359b4b05b114e760088026; 
assign Ic677b8f221359b4b05b114e760088026 = 
        y_nr_in[1] ^ 
        y_nr_in[7] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
        y_nr_in[45] ^ 
0; 



wire I65ba49fe883c3799a2bb0c4b9c721d9a; 
assign I65ba49fe883c3799a2bb0c4b9c721d9a = 
        y_nr_in[62] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[22] = 
Ic677b8f221359b4b05b114e760088026 ^ 
I65ba49fe883c3799a2bb0c4b9c721d9a ^ 
0; 



wire Ic7d0f4caa039b2afeb85d8fb2076370f; 
assign Ic7d0f4caa039b2afeb85d8fb2076370f = 
        y_nr_in[2] ^ 
        y_nr_in[4] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
        y_nr_in[46] ^ 
0; 



wire Ie2707d69382156df60f572f42fef6d82; 
assign Ie2707d69382156df60f572f42fef6d82 = 
        y_nr_in[63] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[23] = 
Ic7d0f4caa039b2afeb85d8fb2076370f ^ 
Ie2707d69382156df60f572f42fef6d82 ^ 
0; 



wire Ic3eccf6c7eca6c5e359fad33ea91c2f6; 
assign Ic3eccf6c7eca6c5e359fad33ea91c2f6 = 
        y_nr_in[3] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
        y_nr_in[36] ^ 
        y_nr_in[46] ^ 
0; 



wire I8e466d425aaf25aa381d135c1c0e15bb; 
assign I8e466d425aaf25aa381d135c1c0e15bb = 
        y_nr_in[64] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[24] = 
Ic3eccf6c7eca6c5e359fad33ea91c2f6 ^ 
I8e466d425aaf25aa381d135c1c0e15bb ^ 
0; 



wire Ie7a7f6d008bab98310894fefe850f9f2; 
assign Ie7a7f6d008bab98310894fefe850f9f2 = 
        y_nr_in[0] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
        y_nr_in[37] ^ 
        y_nr_in[47] ^ 
0; 



wire I1eb9e6ded618528afb132c0fb1d0c693; 
assign I1eb9e6ded618528afb132c0fb1d0c693 = 
        y_nr_in[65] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[25] = 
Ie7a7f6d008bab98310894fefe850f9f2 ^ 
I1eb9e6ded618528afb132c0fb1d0c693 ^ 
0; 



wire I32b9dea9070f1dde87ba8f0f85522fe8; 
assign I32b9dea9070f1dde87ba8f0f85522fe8 = 
        y_nr_in[1] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
        y_nr_in[38] ^ 
        y_nr_in[44] ^ 
0; 



wire I49feeb0e192ad2bd21922b53d5a7934f; 
assign I49feeb0e192ad2bd21922b53d5a7934f = 
        y_nr_in[66] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[26] = 
I32b9dea9070f1dde87ba8f0f85522fe8 ^ 
I49feeb0e192ad2bd21922b53d5a7934f ^ 
0; 



wire I60c9aa445b88a587ac9d690a6d461fb0; 
assign I60c9aa445b88a587ac9d690a6d461fb0 = 
        y_nr_in[2] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
        y_nr_in[39] ^ 
        y_nr_in[45] ^ 
0; 



wire Ic687128ec1afce062367ea23d2443dbf; 
assign Ic687128ec1afce062367ea23d2443dbf = 
        y_nr_in[67] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[27] = 
I60c9aa445b88a587ac9d690a6d461fb0 ^ 
Ic687128ec1afce062367ea23d2443dbf ^ 
0; 



wire I58ab5a30327f79a04753ef0a898f8d61; 
assign I58ab5a30327f79a04753ef0a898f8d61 = 
        y_nr_in[5] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
        y_nr_in[47] ^ 
        y_nr_in[52] ^ 
0; 



wire I737fb7996b130ed186f11f93f757a2c3; 
assign I737fb7996b130ed186f11f93f757a2c3 = 
        y_nr_in[68] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[28] = 
I58ab5a30327f79a04753ef0a898f8d61 ^ 
I737fb7996b130ed186f11f93f757a2c3 ^ 
0; 



wire I79f33d19781dda0516767ab237d2e5b5; 
assign I79f33d19781dda0516767ab237d2e5b5 = 
        y_nr_in[6] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
        y_nr_in[44] ^ 
        y_nr_in[53] ^ 
0; 



wire I26a5712a6166f08c0ece9115cc2b4217; 
assign I26a5712a6166f08c0ece9115cc2b4217 = 
        y_nr_in[69] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[29] = 
I79f33d19781dda0516767ab237d2e5b5 ^ 
I26a5712a6166f08c0ece9115cc2b4217 ^ 
0; 



wire I999b8fea9de99304c0f32ccf85e8fe35; 
assign I999b8fea9de99304c0f32ccf85e8fe35 = 
        y_nr_in[7] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
        y_nr_in[45] ^ 
        y_nr_in[54] ^ 
0; 



wire I9ed433f3241bd10fd8e845ea9fbbbaf1; 
assign I9ed433f3241bd10fd8e845ea9fbbbaf1 = 
        y_nr_in[70] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[30] = 
I999b8fea9de99304c0f32ccf85e8fe35 ^ 
I9ed433f3241bd10fd8e845ea9fbbbaf1 ^ 
0; 



wire I8133c1f62bebb9a28addbaebd3d64928; 
assign I8133c1f62bebb9a28addbaebd3d64928 = 
        y_nr_in[4] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
        y_nr_in[46] ^ 
        y_nr_in[55] ^ 
0; 



wire I6e79baebb440527a660a6a84d5d0aede; 
assign I6e79baebb440527a660a6a84d5d0aede = 
        y_nr_in[71] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[31] = 
I8133c1f62bebb9a28addbaebd3d64928 ^ 
I6e79baebb440527a660a6a84d5d0aede ^ 
0; 



wire I0a4e21b1e023bb1edb52d2ff7d1da294; 
assign I0a4e21b1e023bb1edb52d2ff7d1da294 = 
        y_nr_in[2] ^ 
        y_nr_in[6] ^ 
        y_nr_in[50] ^ 
        y_nr_in[72] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[32] = 
I0a4e21b1e023bb1edb52d2ff7d1da294 ^ 
0; 



wire I2b6d676d44737efc41dd40dcac0419e6; 
assign I2b6d676d44737efc41dd40dcac0419e6 = 
        y_nr_in[3] ^ 
        y_nr_in[7] ^ 
        y_nr_in[51] ^ 
        y_nr_in[73] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[33] = 
I2b6d676d44737efc41dd40dcac0419e6 ^ 
0; 



wire I92b61b2776bf0f9c25a28925f8d7b977; 
assign I92b61b2776bf0f9c25a28925f8d7b977 = 
        y_nr_in[0] ^ 
        y_nr_in[4] ^ 
        y_nr_in[48] ^ 
        y_nr_in[74] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[34] = 
I92b61b2776bf0f9c25a28925f8d7b977 ^ 
0; 



wire If70b9fb4df54006b0cd207ef0494ff34; 
assign If70b9fb4df54006b0cd207ef0494ff34 = 
        y_nr_in[1] ^ 
        y_nr_in[5] ^ 
        y_nr_in[49] ^ 
        y_nr_in[75] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[35] = 
If70b9fb4df54006b0cd207ef0494ff34 ^ 
0; 



wire I8d794790ffdcbf7953586b3eb99358f5; 
assign I8d794790ffdcbf7953586b3eb99358f5 = 
        y_nr_in[7] ^ 
        y_nr_in[33] ^ 
        y_nr_in[41] ^ 
        y_nr_in[47] ^ 
        y_nr_in[76] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[36] = 
I8d794790ffdcbf7953586b3eb99358f5 ^ 
0; 



wire Ib08d9fde464d1fa679ec711509c4dfd4; 
assign Ib08d9fde464d1fa679ec711509c4dfd4 = 
        y_nr_in[4] ^ 
        y_nr_in[34] ^ 
        y_nr_in[42] ^ 
        y_nr_in[44] ^ 
        y_nr_in[77] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[37] = 
Ib08d9fde464d1fa679ec711509c4dfd4 ^ 
0; 



wire I5205a99fc8c12ff619a1f282f4ca3377; 
assign I5205a99fc8c12ff619a1f282f4ca3377 = 
        y_nr_in[5] ^ 
        y_nr_in[35] ^ 
        y_nr_in[43] ^ 
        y_nr_in[45] ^ 
        y_nr_in[78] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[38] = 
I5205a99fc8c12ff619a1f282f4ca3377 ^ 
0; 



wire Icfb334e065bf257c870f207e495ac5f4; 
assign Icfb334e065bf257c870f207e495ac5f4 = 
        y_nr_in[6] ^ 
        y_nr_in[32] ^ 
        y_nr_in[40] ^ 
        y_nr_in[46] ^ 
        y_nr_in[79] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[39] = 
Icfb334e065bf257c870f207e495ac5f4 ^ 
0; 



wire I4404102e5bf39203979d969c30a30b08; 
assign I4404102e5bf39203979d969c30a30b08 = 
        y_nr_in[3] ^ 
        y_nr_in[5] ^ 
        y_nr_in[24] ^ 
        y_nr_in[29] ^ 
        y_nr_in[80] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[40] = 
I4404102e5bf39203979d969c30a30b08 ^ 
0; 



wire I93296f6aa6d631cbe0d2f8e1b0c7e080; 
assign I93296f6aa6d631cbe0d2f8e1b0c7e080 = 
        y_nr_in[0] ^ 
        y_nr_in[6] ^ 
        y_nr_in[25] ^ 
        y_nr_in[30] ^ 
        y_nr_in[81] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[41] = 
I93296f6aa6d631cbe0d2f8e1b0c7e080 ^ 
0; 



wire I2180ac538cb197b0cf0c4705b0ddecf4; 
assign I2180ac538cb197b0cf0c4705b0ddecf4 = 
        y_nr_in[1] ^ 
        y_nr_in[7] ^ 
        y_nr_in[26] ^ 
        y_nr_in[31] ^ 
        y_nr_in[82] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[42] = 
I2180ac538cb197b0cf0c4705b0ddecf4 ^ 
0; 



wire I8d51ab0cca28a45d30149217fe0a81e4; 
assign I8d51ab0cca28a45d30149217fe0a81e4 = 
        y_nr_in[2] ^ 
        y_nr_in[4] ^ 
        y_nr_in[27] ^ 
        y_nr_in[28] ^ 
        y_nr_in[83] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[43] = 
I8d51ab0cca28a45d30149217fe0a81e4 ^ 
0; 



wire I9f830d3f7bdd988590974d2408c85a2a; 
assign I9f830d3f7bdd988590974d2408c85a2a = 
        y_nr_in[3] ^ 
        y_nr_in[28] ^ 
        y_nr_in[38] ^ 
        y_nr_in[52] ^ 
        y_nr_in[84] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[44] = 
I9f830d3f7bdd988590974d2408c85a2a ^ 
0; 



wire I58631a056b50ae0f45852849cfd5ae0c; 
assign I58631a056b50ae0f45852849cfd5ae0c = 
        y_nr_in[0] ^ 
        y_nr_in[29] ^ 
        y_nr_in[39] ^ 
        y_nr_in[53] ^ 
        y_nr_in[85] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[45] = 
I58631a056b50ae0f45852849cfd5ae0c ^ 
0; 



wire Ibae0f4738d52d9236789e9a624a549fe; 
assign Ibae0f4738d52d9236789e9a624a549fe = 
        y_nr_in[1] ^ 
        y_nr_in[30] ^ 
        y_nr_in[36] ^ 
        y_nr_in[54] ^ 
        y_nr_in[86] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[46] = 
Ibae0f4738d52d9236789e9a624a549fe ^ 
0; 



wire I7e54959fb12dfe41d92a70d5d5ab5f3a; 
assign I7e54959fb12dfe41d92a70d5d5ab5f3a = 
        y_nr_in[2] ^ 
        y_nr_in[31] ^ 
        y_nr_in[37] ^ 
        y_nr_in[55] ^ 
        y_nr_in[87] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[47] = 
I7e54959fb12dfe41d92a70d5d5ab5f3a ^ 
0; 



wire Iad6a3ea7209fd923008860221631b0d4; 
assign Iad6a3ea7209fd923008860221631b0d4 = 
        y_nr_in[7] ^ 
        y_nr_in[15] ^ 
        y_nr_in[46] ^ 
        y_nr_in[88] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[48] = 
Iad6a3ea7209fd923008860221631b0d4 ^ 
0; 



wire I929b2b75e148c3e735bc3ffd0c735c4c; 
assign I929b2b75e148c3e735bc3ffd0c735c4c = 
        y_nr_in[4] ^ 
        y_nr_in[12] ^ 
        y_nr_in[47] ^ 
        y_nr_in[89] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[49] = 
I929b2b75e148c3e735bc3ffd0c735c4c ^ 
0; 



wire I889ca4e5a809c19e1c0c366c763c6dff; 
assign I889ca4e5a809c19e1c0c366c763c6dff = 
        y_nr_in[5] ^ 
        y_nr_in[13] ^ 
        y_nr_in[44] ^ 
        y_nr_in[90] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[50] = 
I889ca4e5a809c19e1c0c366c763c6dff ^ 
0; 



wire I90556dfbde663aefa9c004e080bc5ebc; 
assign I90556dfbde663aefa9c004e080bc5ebc = 
        y_nr_in[6] ^ 
        y_nr_in[14] ^ 
        y_nr_in[45] ^ 
        y_nr_in[91] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[51] = 
I90556dfbde663aefa9c004e080bc5ebc ^ 
0; 



wire Idef9c3d3b6b9dc9d75d4b2d70756a014; 
assign Idef9c3d3b6b9dc9d75d4b2d70756a014 = 
        y_nr_in[3] ^ 
        y_nr_in[6] ^ 
        y_nr_in[34] ^ 
        y_nr_in[54] ^ 
        y_nr_in[92] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[52] = 
Idef9c3d3b6b9dc9d75d4b2d70756a014 ^ 
0; 



wire I59e33a88645895fa470fd8b5f8e3d1cc; 
assign I59e33a88645895fa470fd8b5f8e3d1cc = 
        y_nr_in[0] ^ 
        y_nr_in[7] ^ 
        y_nr_in[35] ^ 
        y_nr_in[55] ^ 
        y_nr_in[93] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[53] = 
I59e33a88645895fa470fd8b5f8e3d1cc ^ 
0; 



wire I228b7aed69ff4ffb5d1f5133f4c11e10; 
assign I228b7aed69ff4ffb5d1f5133f4c11e10 = 
        y_nr_in[1] ^ 
        y_nr_in[4] ^ 
        y_nr_in[32] ^ 
        y_nr_in[52] ^ 
        y_nr_in[94] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[54] = 
I228b7aed69ff4ffb5d1f5133f4c11e10 ^ 
0; 



wire I41785b0035f0bb83aea0b6cebd41962f; 
assign I41785b0035f0bb83aea0b6cebd41962f = 
        y_nr_in[2] ^ 
        y_nr_in[5] ^ 
        y_nr_in[33] ^ 
        y_nr_in[53] ^ 
        y_nr_in[95] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[55] = 
I41785b0035f0bb83aea0b6cebd41962f ^ 
0; 



wire If3ab999799a1eba48193657f6a470f44; 
assign If3ab999799a1eba48193657f6a470f44 = 
        y_nr_in[7] ^ 
        y_nr_in[25] ^ 
        y_nr_in[47] ^ 
        y_nr_in[52] ^ 
        y_nr_in[96] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[56] = 
If3ab999799a1eba48193657f6a470f44 ^ 
0; 



wire I98295432b77f6baf07da6c5d54a6bf85; 
assign I98295432b77f6baf07da6c5d54a6bf85 = 
        y_nr_in[4] ^ 
        y_nr_in[26] ^ 
        y_nr_in[44] ^ 
        y_nr_in[53] ^ 
        y_nr_in[97] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[57] = 
I98295432b77f6baf07da6c5d54a6bf85 ^ 
0; 



wire Ia5599d3d02f47feddf15cac50efc11ac; 
assign Ia5599d3d02f47feddf15cac50efc11ac = 
        y_nr_in[5] ^ 
        y_nr_in[27] ^ 
        y_nr_in[45] ^ 
        y_nr_in[54] ^ 
        y_nr_in[98] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[58] = 
Ia5599d3d02f47feddf15cac50efc11ac ^ 
0; 



wire I5a77920d43f226b7ab7aaf1053363aba; 
assign I5a77920d43f226b7ab7aaf1053363aba = 
        y_nr_in[6] ^ 
        y_nr_in[24] ^ 
        y_nr_in[46] ^ 
        y_nr_in[55] ^ 
        y_nr_in[99] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[59] = 
I5a77920d43f226b7ab7aaf1053363aba ^ 
0; 



wire I8d99e973e3d281fad7037214dcfa04fe; 
assign I8d99e973e3d281fad7037214dcfa04fe = 
        y_nr_in[3] ^ 
        y_nr_in[43] ^ 
        y_nr_in[45] ^ 
        y_nr_in[100] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[60] = 
I8d99e973e3d281fad7037214dcfa04fe ^ 
0; 



wire Ida129ff582ace5f9691c239858fbab4c; 
assign Ida129ff582ace5f9691c239858fbab4c = 
        y_nr_in[0] ^ 
        y_nr_in[40] ^ 
        y_nr_in[46] ^ 
        y_nr_in[101] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[61] = 
Ida129ff582ace5f9691c239858fbab4c ^ 
0; 



wire I412e480850ab5d1ccd3ccbf4306bfe05; 
assign I412e480850ab5d1ccd3ccbf4306bfe05 = 
        y_nr_in[1] ^ 
        y_nr_in[41] ^ 
        y_nr_in[47] ^ 
        y_nr_in[102] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[62] = 
I412e480850ab5d1ccd3ccbf4306bfe05 ^ 
0; 



wire Icc2d8eb756016564495467427ac1bb1c; 
assign Icc2d8eb756016564495467427ac1bb1c = 
        y_nr_in[2] ^ 
        y_nr_in[42] ^ 
        y_nr_in[44] ^ 
        y_nr_in[103] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[63] = 
Icc2d8eb756016564495467427ac1bb1c ^ 
0; 



wire Iafdddb183bf157e29ed9c4323987304b; 
assign Iafdddb183bf157e29ed9c4323987304b = 
        y_nr_in[7] ^ 
        y_nr_in[38] ^ 
        y_nr_in[44] ^ 
        y_nr_in[50] ^ 
        y_nr_in[104] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[64] = 
Iafdddb183bf157e29ed9c4323987304b ^ 
0; 



wire Iad54e785c16eb6c2b8b9712e1fe9bc32; 
assign Iad54e785c16eb6c2b8b9712e1fe9bc32 = 
        y_nr_in[4] ^ 
        y_nr_in[39] ^ 
        y_nr_in[45] ^ 
        y_nr_in[51] ^ 
        y_nr_in[105] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[65] = 
Iad54e785c16eb6c2b8b9712e1fe9bc32 ^ 
0; 



wire I7afbdbb080d3398ffdb66312340bb529; 
assign I7afbdbb080d3398ffdb66312340bb529 = 
        y_nr_in[5] ^ 
        y_nr_in[36] ^ 
        y_nr_in[46] ^ 
        y_nr_in[48] ^ 
        y_nr_in[106] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[66] = 
I7afbdbb080d3398ffdb66312340bb529 ^ 
0; 



wire I4f3f8325af4f5d639c72c0368b0906b8; 
assign I4f3f8325af4f5d639c72c0368b0906b8 = 
        y_nr_in[6] ^ 
        y_nr_in[37] ^ 
        y_nr_in[47] ^ 
        y_nr_in[49] ^ 
        y_nr_in[107] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[67] = 
I4f3f8325af4f5d639c72c0368b0906b8 ^ 
0; 



wire I17397105dd7c843430a11c1354eec772; 
assign I17397105dd7c843430a11c1354eec772 = 
        y_nr_in[6] ^ 
        y_nr_in[20] ^ 
        y_nr_in[46] ^ 
        y_nr_in[48] ^ 
        y_nr_in[108] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[68] = 
I17397105dd7c843430a11c1354eec772 ^ 
0; 



wire Ib838d5bbc18e72e791bf34bed1e3375b; 
assign Ib838d5bbc18e72e791bf34bed1e3375b = 
        y_nr_in[7] ^ 
        y_nr_in[21] ^ 
        y_nr_in[47] ^ 
        y_nr_in[49] ^ 
        y_nr_in[109] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[69] = 
Ib838d5bbc18e72e791bf34bed1e3375b ^ 
0; 



wire I69c3dd09a1a064e92fd5ec315e100e00; 
assign I69c3dd09a1a064e92fd5ec315e100e00 = 
        y_nr_in[4] ^ 
        y_nr_in[22] ^ 
        y_nr_in[44] ^ 
        y_nr_in[50] ^ 
        y_nr_in[110] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[70] = 
I69c3dd09a1a064e92fd5ec315e100e00 ^ 
0; 



wire I18aa40d35da802303236196a5177d333; 
assign I18aa40d35da802303236196a5177d333 = 
        y_nr_in[5] ^ 
        y_nr_in[23] ^ 
        y_nr_in[45] ^ 
        y_nr_in[51] ^ 
        y_nr_in[111] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[71] = 
I18aa40d35da802303236196a5177d333 ^ 
0; 



wire I81781416a91b3cae8dead2fc966b5baa; 
assign I81781416a91b3cae8dead2fc966b5baa = 
        y_nr_in[0] ^ 
        y_nr_in[26] ^ 
        y_nr_in[30] ^ 
        y_nr_in[112] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[72] = 
I81781416a91b3cae8dead2fc966b5baa ^ 
0; 



wire Ie3def9ad89d976bc39eae9bb13cc710b; 
assign Ie3def9ad89d976bc39eae9bb13cc710b = 
        y_nr_in[1] ^ 
        y_nr_in[27] ^ 
        y_nr_in[31] ^ 
        y_nr_in[113] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[73] = 
Ie3def9ad89d976bc39eae9bb13cc710b ^ 
0; 



wire I8f69316d0b78574f5dfa08c70875442a; 
assign I8f69316d0b78574f5dfa08c70875442a = 
        y_nr_in[2] ^ 
        y_nr_in[24] ^ 
        y_nr_in[28] ^ 
        y_nr_in[114] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[74] = 
I8f69316d0b78574f5dfa08c70875442a ^ 
0; 



wire I17230e178a47c5138b98e398ba6e7c8b; 
assign I17230e178a47c5138b98e398ba6e7c8b = 
        y_nr_in[3] ^ 
        y_nr_in[25] ^ 
        y_nr_in[29] ^ 
        y_nr_in[115] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[75] = 
I17230e178a47c5138b98e398ba6e7c8b ^ 
0; 



wire I1dbf2ce97a856912e1520b954179e523; 
assign I1dbf2ce97a856912e1520b954179e523 = 
        y_nr_in[3] ^ 
        y_nr_in[4] ^ 
        y_nr_in[41] ^ 
        y_nr_in[116] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[76] = 
I1dbf2ce97a856912e1520b954179e523 ^ 
0; 



wire I4555e8bbe7220ef88a4b7c99ab747c06; 
assign I4555e8bbe7220ef88a4b7c99ab747c06 = 
        y_nr_in[0] ^ 
        y_nr_in[5] ^ 
        y_nr_in[42] ^ 
        y_nr_in[117] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[77] = 
I4555e8bbe7220ef88a4b7c99ab747c06 ^ 
0; 



wire Ic312ea4981841bfb8c45afde83c3408c; 
assign Ic312ea4981841bfb8c45afde83c3408c = 
        y_nr_in[1] ^ 
        y_nr_in[6] ^ 
        y_nr_in[43] ^ 
        y_nr_in[118] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[78] = 
Ic312ea4981841bfb8c45afde83c3408c ^ 
0; 



wire I6030957820002aa576f92acfd56391fa; 
assign I6030957820002aa576f92acfd56391fa = 
        y_nr_in[2] ^ 
        y_nr_in[7] ^ 
        y_nr_in[40] ^ 
        y_nr_in[119] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[79] = 
I6030957820002aa576f92acfd56391fa ^ 
0; 



wire I1c32e62de8804d077d57d03d02c79cb3; 
assign I1c32e62de8804d077d57d03d02c79cb3 = 
        y_nr_in[6] ^ 
        y_nr_in[17] ^ 
        y_nr_in[45] ^ 
        y_nr_in[120] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[80] = 
I1c32e62de8804d077d57d03d02c79cb3 ^ 
0; 



wire I338a51204679def922c0cfb9231f7037; 
assign I338a51204679def922c0cfb9231f7037 = 
        y_nr_in[7] ^ 
        y_nr_in[18] ^ 
        y_nr_in[46] ^ 
        y_nr_in[121] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[81] = 
I338a51204679def922c0cfb9231f7037 ^ 
0; 



wire I6a8ea57981879d3ef59eb44ad7794f46; 
assign I6a8ea57981879d3ef59eb44ad7794f46 = 
        y_nr_in[4] ^ 
        y_nr_in[19] ^ 
        y_nr_in[47] ^ 
        y_nr_in[122] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[82] = 
I6a8ea57981879d3ef59eb44ad7794f46 ^ 
0; 



wire I3b16e5275a15e94b36df84e4dde0c841; 
assign I3b16e5275a15e94b36df84e4dde0c841 = 
        y_nr_in[5] ^ 
        y_nr_in[16] ^ 
        y_nr_in[44] ^ 
        y_nr_in[123] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[83] = 
I3b16e5275a15e94b36df84e4dde0c841 ^ 
0; 



wire Ibdadb99746c7b49d48cac8789bf7e150; 
assign Ibdadb99746c7b49d48cac8789bf7e150 = 
        y_nr_in[0] ^ 
        y_nr_in[34] ^ 
        y_nr_in[54] ^ 
        y_nr_in[124] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[84] = 
Ibdadb99746c7b49d48cac8789bf7e150 ^ 
0; 



wire Ifc8e81bc5164edc24bb598e85f6e6f9d; 
assign Ifc8e81bc5164edc24bb598e85f6e6f9d = 
        y_nr_in[1] ^ 
        y_nr_in[35] ^ 
        y_nr_in[55] ^ 
        y_nr_in[125] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[85] = 
Ifc8e81bc5164edc24bb598e85f6e6f9d ^ 
0; 



wire I93dd82883fcab2cc199de5b04e0daa65; 
assign I93dd82883fcab2cc199de5b04e0daa65 = 
        y_nr_in[2] ^ 
        y_nr_in[32] ^ 
        y_nr_in[52] ^ 
        y_nr_in[126] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[86] = 
I93dd82883fcab2cc199de5b04e0daa65 ^ 
0; 



wire I0df496d01c662296bf9c8285dc76355f; 
assign I0df496d01c662296bf9c8285dc76355f = 
        y_nr_in[3] ^ 
        y_nr_in[33] ^ 
        y_nr_in[53] ^ 
        y_nr_in[127] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[87] = 
I0df496d01c662296bf9c8285dc76355f ^ 
0; 



wire Ie568d06d2b66ced1be7d951b479fbf9b; 
assign Ie568d06d2b66ced1be7d951b479fbf9b = 
        y_nr_in[6] ^ 
        y_nr_in[11] ^ 
        y_nr_in[128] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[88] = 
Ie568d06d2b66ced1be7d951b479fbf9b ^ 
0; 



wire I652145e8d8909699cf2e62012f2888a1; 
assign I652145e8d8909699cf2e62012f2888a1 = 
        y_nr_in[7] ^ 
        y_nr_in[8] ^ 
        y_nr_in[129] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[89] = 
I652145e8d8909699cf2e62012f2888a1 ^ 
0; 



wire Ibc157aaf0ab31bae42517726c57f6822; 
assign Ibc157aaf0ab31bae42517726c57f6822 = 
        y_nr_in[4] ^ 
        y_nr_in[9] ^ 
        y_nr_in[130] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[90] = 
Ibc157aaf0ab31bae42517726c57f6822 ^ 
0; 



wire I99b784aa0f76968cd7f1c5aa3585f01c; 
assign I99b784aa0f76968cd7f1c5aa3585f01c = 
        y_nr_in[5] ^ 
        y_nr_in[10] ^ 
        y_nr_in[131] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[91] = 
I99b784aa0f76968cd7f1c5aa3585f01c ^ 
0; 



wire I987e716719b1ee4fae7a4cf87443693d; 
assign I987e716719b1ee4fae7a4cf87443693d = 
        y_nr_in[3] ^ 
        y_nr_in[15] ^ 
        y_nr_in[22] ^ 
        y_nr_in[132] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[92] = 
I987e716719b1ee4fae7a4cf87443693d ^ 
0; 



wire Ia5e8b3f8cbec23457548ca09840bdb2e; 
assign Ia5e8b3f8cbec23457548ca09840bdb2e = 
        y_nr_in[0] ^ 
        y_nr_in[12] ^ 
        y_nr_in[23] ^ 
        y_nr_in[133] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[93] = 
Ia5e8b3f8cbec23457548ca09840bdb2e ^ 
0; 



wire I48848ec661e0f6d8a2916f0fa5e2c317; 
assign I48848ec661e0f6d8a2916f0fa5e2c317 = 
        y_nr_in[1] ^ 
        y_nr_in[13] ^ 
        y_nr_in[20] ^ 
        y_nr_in[134] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[94] = 
I48848ec661e0f6d8a2916f0fa5e2c317 ^ 
0; 



wire Ibe1d577080dafadb1d35924d8328dcbf; 
assign Ibe1d577080dafadb1d35924d8328dcbf = 
        y_nr_in[2] ^ 
        y_nr_in[14] ^ 
        y_nr_in[21] ^ 
        y_nr_in[135] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[95] = 
Ibe1d577080dafadb1d35924d8328dcbf ^ 
0; 



wire Ifa3b588c73b1d3f0f7a3b77f3bedd969; 
assign Ifa3b588c73b1d3f0f7a3b77f3bedd969 = 
        y_nr_in[6] ^ 
        y_nr_in[11] ^ 
        y_nr_in[36] ^ 
        y_nr_in[136] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[96] = 
Ifa3b588c73b1d3f0f7a3b77f3bedd969 ^ 
0; 



wire I74d793aaedd2d17ca1ac5c28d8e00ddc; 
assign I74d793aaedd2d17ca1ac5c28d8e00ddc = 
        y_nr_in[7] ^ 
        y_nr_in[8] ^ 
        y_nr_in[37] ^ 
        y_nr_in[137] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[97] = 
I74d793aaedd2d17ca1ac5c28d8e00ddc ^ 
0; 



wire I89d73c6136fc7cf9bef28b54bce4448d; 
assign I89d73c6136fc7cf9bef28b54bce4448d = 
        y_nr_in[4] ^ 
        y_nr_in[9] ^ 
        y_nr_in[38] ^ 
        y_nr_in[138] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[98] = 
I89d73c6136fc7cf9bef28b54bce4448d ^ 
0; 



wire I82a05805c0383b4b7e9d18984b5bcd3a; 
assign I82a05805c0383b4b7e9d18984b5bcd3a = 
        y_nr_in[5] ^ 
        y_nr_in[10] ^ 
        y_nr_in[39] ^ 
        y_nr_in[139] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[99] = 
I82a05805c0383b4b7e9d18984b5bcd3a ^ 
0; 



wire I9128871fae777e06bbb350a72e6f9e4f; 
assign I9128871fae777e06bbb350a72e6f9e4f = 
        y_nr_in[0] ^ 
        y_nr_in[20] ^ 
        y_nr_in[140] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[100] = 
I9128871fae777e06bbb350a72e6f9e4f ^ 
0; 



wire Ic50a2c7df181f1045665db84f646594f; 
assign Ic50a2c7df181f1045665db84f646594f = 
        y_nr_in[1] ^ 
        y_nr_in[21] ^ 
        y_nr_in[141] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[101] = 
Ic50a2c7df181f1045665db84f646594f ^ 
0; 



wire If347375c829c8b65105d9248d021d5b8; 
assign If347375c829c8b65105d9248d021d5b8 = 
        y_nr_in[2] ^ 
        y_nr_in[22] ^ 
        y_nr_in[142] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[102] = 
If347375c829c8b65105d9248d021d5b8 ^ 
0; 



wire I4ae6273b0782c4c1ec5c0c50bf65f1bc; 
assign I4ae6273b0782c4c1ec5c0c50bf65f1bc = 
        y_nr_in[3] ^ 
        y_nr_in[23] ^ 
        y_nr_in[143] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[103] = 
I4ae6273b0782c4c1ec5c0c50bf65f1bc ^ 
0; 



wire I874aaaaaf5989e844a752550d5745ad9; 
assign I874aaaaaf5989e844a752550d5745ad9 = 
        y_nr_in[9] ^ 
        y_nr_in[31] ^ 
        y_nr_in[48] ^ 
        y_nr_in[54] ^ 
        y_nr_in[144] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[104] = 
I874aaaaaf5989e844a752550d5745ad9 ^ 
0; 



wire Iada01caae18d74509024f59711ccc9f2; 
assign Iada01caae18d74509024f59711ccc9f2 = 
        y_nr_in[10] ^ 
        y_nr_in[28] ^ 
        y_nr_in[49] ^ 
        y_nr_in[55] ^ 
        y_nr_in[145] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[105] = 
Iada01caae18d74509024f59711ccc9f2 ^ 
0; 



wire I0e529a3e23121b53803627cb083b838a; 
assign I0e529a3e23121b53803627cb083b838a = 
        y_nr_in[11] ^ 
        y_nr_in[29] ^ 
        y_nr_in[50] ^ 
        y_nr_in[52] ^ 
        y_nr_in[146] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[106] = 
I0e529a3e23121b53803627cb083b838a ^ 
0; 



wire I2863b9ccaca74b299d63ccb3aa1008c3; 
assign I2863b9ccaca74b299d63ccb3aa1008c3 = 
        y_nr_in[8] ^ 
        y_nr_in[30] ^ 
        y_nr_in[51] ^ 
        y_nr_in[53] ^ 
        y_nr_in[147] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[107] = 
I2863b9ccaca74b299d63ccb3aa1008c3 ^ 
0; 



wire Ia5b2fbfa58545fac2334f4f3d43b403c; 
assign Ia5b2fbfa58545fac2334f4f3d43b403c = 
        y_nr_in[0] ^ 
        y_nr_in[27] ^ 
        y_nr_in[148] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[108] = 
Ia5b2fbfa58545fac2334f4f3d43b403c ^ 
0; 



wire I177e7f6095ad2c5a43168aa37d4aa977; 
assign I177e7f6095ad2c5a43168aa37d4aa977 = 
        y_nr_in[1] ^ 
        y_nr_in[24] ^ 
        y_nr_in[149] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[109] = 
I177e7f6095ad2c5a43168aa37d4aa977 ^ 
0; 



wire I992dff0e62ca4039f019a31daa95ae09; 
assign I992dff0e62ca4039f019a31daa95ae09 = 
        y_nr_in[2] ^ 
        y_nr_in[25] ^ 
        y_nr_in[150] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[110] = 
I992dff0e62ca4039f019a31daa95ae09 ^ 
0; 



wire Ib2cbff7b947445399e30aefa3f01a6c5; 
assign Ib2cbff7b947445399e30aefa3f01a6c5 = 
        y_nr_in[3] ^ 
        y_nr_in[26] ^ 
        y_nr_in[151] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[111] = 
Ib2cbff7b947445399e30aefa3f01a6c5 ^ 
0; 



wire I9c2ba3d90c02993ad371600f7c01a4e5; 
assign I9c2ba3d90c02993ad371600f7c01a4e5 = 
        y_nr_in[6] ^ 
        y_nr_in[9] ^ 
        y_nr_in[23] ^ 
        y_nr_in[152] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[112] = 
I9c2ba3d90c02993ad371600f7c01a4e5 ^ 
0; 



wire I8a89007134bcb3bec1d4715e2515b9fe; 
assign I8a89007134bcb3bec1d4715e2515b9fe = 
        y_nr_in[7] ^ 
        y_nr_in[10] ^ 
        y_nr_in[20] ^ 
        y_nr_in[153] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[113] = 
I8a89007134bcb3bec1d4715e2515b9fe ^ 
0; 



wire I84a2bfe393b23e3c218f3b8a268fcc40; 
assign I84a2bfe393b23e3c218f3b8a268fcc40 = 
        y_nr_in[4] ^ 
        y_nr_in[11] ^ 
        y_nr_in[21] ^ 
        y_nr_in[154] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[114] = 
I84a2bfe393b23e3c218f3b8a268fcc40 ^ 
0; 



wire I17adba6aa9d903b7961ca91a44456b86; 
assign I17adba6aa9d903b7961ca91a44456b86 = 
        y_nr_in[5] ^ 
        y_nr_in[8] ^ 
        y_nr_in[22] ^ 
        y_nr_in[155] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[115] = 
I17adba6aa9d903b7961ca91a44456b86 ^ 
0; 



wire Id72f6ff2b857eccbeb2d68cdb48b565e; 
assign Id72f6ff2b857eccbeb2d68cdb48b565e = 
        y_nr_in[2] ^ 
        y_nr_in[16] ^ 
        y_nr_in[156] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[116] = 
Id72f6ff2b857eccbeb2d68cdb48b565e ^ 
0; 



wire I09d47b16a82326c3ca630fc2f95fe003; 
assign I09d47b16a82326c3ca630fc2f95fe003 = 
        y_nr_in[3] ^ 
        y_nr_in[17] ^ 
        y_nr_in[157] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[117] = 
I09d47b16a82326c3ca630fc2f95fe003 ^ 
0; 



wire Ifeb5ad5815b4cab0cdec106d941b2bc3; 
assign Ifeb5ad5815b4cab0cdec106d941b2bc3 = 
        y_nr_in[0] ^ 
        y_nr_in[18] ^ 
        y_nr_in[158] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[118] = 
Ifeb5ad5815b4cab0cdec106d941b2bc3 ^ 
0; 



wire Ie5a64dc98a03056cd6d4d689e75cda62; 
assign Ie5a64dc98a03056cd6d4d689e75cda62 = 
        y_nr_in[1] ^ 
        y_nr_in[19] ^ 
        y_nr_in[159] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[119] = 
Ie5a64dc98a03056cd6d4d689e75cda62 ^ 
0; 



wire I6d78420ca46fc92155be2d1351b7f11a; 
assign I6d78420ca46fc92155be2d1351b7f11a = 
        y_nr_in[11] ^ 
        y_nr_in[20] ^ 
        y_nr_in[29] ^ 
        y_nr_in[36] ^ 
        y_nr_in[160] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[120] = 
I6d78420ca46fc92155be2d1351b7f11a ^ 
0; 



wire Ic5308709c54362a205dbbd582a32955b; 
assign Ic5308709c54362a205dbbd582a32955b = 
        y_nr_in[8] ^ 
        y_nr_in[21] ^ 
        y_nr_in[30] ^ 
        y_nr_in[37] ^ 
        y_nr_in[161] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[121] = 
Ic5308709c54362a205dbbd582a32955b ^ 
0; 



wire Ieae049479d0089894db606d224ec1bb3; 
assign Ieae049479d0089894db606d224ec1bb3 = 
        y_nr_in[9] ^ 
        y_nr_in[22] ^ 
        y_nr_in[31] ^ 
        y_nr_in[38] ^ 
        y_nr_in[162] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[122] = 
Ieae049479d0089894db606d224ec1bb3 ^ 
0; 



wire I53e13f817c31e7378aa87943111141b1; 
assign I53e13f817c31e7378aa87943111141b1 = 
        y_nr_in[10] ^ 
        y_nr_in[23] ^ 
        y_nr_in[28] ^ 
        y_nr_in[39] ^ 
        y_nr_in[163] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[123] = 
I53e13f817c31e7378aa87943111141b1 ^ 
0; 



wire If0151dacb1b207313fbd59cfbce132f7; 
assign If0151dacb1b207313fbd59cfbce132f7 = 
        y_nr_in[6] ^ 
        y_nr_in[53] ^ 
        y_nr_in[164] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[124] = 
If0151dacb1b207313fbd59cfbce132f7 ^ 
0; 



wire I0e5f8f249f721e14c07e013b3c3a9a87; 
assign I0e5f8f249f721e14c07e013b3c3a9a87 = 
        y_nr_in[7] ^ 
        y_nr_in[54] ^ 
        y_nr_in[165] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[125] = 
I0e5f8f249f721e14c07e013b3c3a9a87 ^ 
0; 



wire I9a26ba97b1ab3a558151e9158f1ace2c; 
assign I9a26ba97b1ab3a558151e9158f1ace2c = 
        y_nr_in[4] ^ 
        y_nr_in[55] ^ 
        y_nr_in[166] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[126] = 
I9a26ba97b1ab3a558151e9158f1ace2c ^ 
0; 



wire I5319fae71e5b003b59ca762f730c8e19; 
assign I5319fae71e5b003b59ca762f730c8e19 = 
        y_nr_in[5] ^ 
        y_nr_in[52] ^ 
        y_nr_in[167] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[127] = 
I5319fae71e5b003b59ca762f730c8e19 ^ 
0; 



wire I3818c5a025045b67cec952da32991301; 
assign I3818c5a025045b67cec952da32991301 = 
        y_nr_in[2] ^ 
        y_nr_in[20] ^ 
        y_nr_in[50] ^ 
        y_nr_in[168] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[128] = 
I3818c5a025045b67cec952da32991301 ^ 
0; 



wire Ia1101d7b28acfef186a853cb29ac4c25; 
assign Ia1101d7b28acfef186a853cb29ac4c25 = 
        y_nr_in[3] ^ 
        y_nr_in[21] ^ 
        y_nr_in[51] ^ 
        y_nr_in[169] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[129] = 
Ia1101d7b28acfef186a853cb29ac4c25 ^ 
0; 



wire Ib3ffea5f22173fe649225d6ab1299efd; 
assign Ib3ffea5f22173fe649225d6ab1299efd = 
        y_nr_in[0] ^ 
        y_nr_in[22] ^ 
        y_nr_in[48] ^ 
        y_nr_in[170] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[130] = 
Ib3ffea5f22173fe649225d6ab1299efd ^ 
0; 



wire I152e78d206482446d9e0349d109db9bb; 
assign I152e78d206482446d9e0349d109db9bb = 
        y_nr_in[1] ^ 
        y_nr_in[23] ^ 
        y_nr_in[49] ^ 
        y_nr_in[171] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[131] = 
I152e78d206482446d9e0349d109db9bb ^ 
0; 



wire I07188611a6e2b9c4860060582f799fc6; 
assign I07188611a6e2b9c4860060582f799fc6 = 
        y_nr_in[8] ^ 
        y_nr_in[28] ^ 
        y_nr_in[43] ^ 
        y_nr_in[172] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[132] = 
I07188611a6e2b9c4860060582f799fc6 ^ 
0; 



wire I18105f6686e85f7d8d0c595d26a0b104; 
assign I18105f6686e85f7d8d0c595d26a0b104 = 
        y_nr_in[9] ^ 
        y_nr_in[29] ^ 
        y_nr_in[40] ^ 
        y_nr_in[173] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[133] = 
I18105f6686e85f7d8d0c595d26a0b104 ^ 
0; 



wire I5902f1dd3b50ab4d94f70cadccdf134e; 
assign I5902f1dd3b50ab4d94f70cadccdf134e = 
        y_nr_in[10] ^ 
        y_nr_in[30] ^ 
        y_nr_in[41] ^ 
        y_nr_in[174] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[134] = 
I5902f1dd3b50ab4d94f70cadccdf134e ^ 
0; 



wire I9cd3ebd61d954b09977f08a24aaad472; 
assign I9cd3ebd61d954b09977f08a24aaad472 = 
        y_nr_in[11] ^ 
        y_nr_in[31] ^ 
        y_nr_in[42] ^ 
        y_nr_in[175] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[135] = 
I9cd3ebd61d954b09977f08a24aaad472 ^ 
0; 



wire I027661fa4b20baf06ed6dd5817aa20f8; 
assign I027661fa4b20baf06ed6dd5817aa20f8 = 
        y_nr_in[3] ^ 
        y_nr_in[49] ^ 
        y_nr_in[52] ^ 
        y_nr_in[176] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[136] = 
I027661fa4b20baf06ed6dd5817aa20f8 ^ 
0; 



wire I9b09625d5954214d3154e7200129e318; 
assign I9b09625d5954214d3154e7200129e318 = 
        y_nr_in[0] ^ 
        y_nr_in[50] ^ 
        y_nr_in[53] ^ 
        y_nr_in[177] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[137] = 
I9b09625d5954214d3154e7200129e318 ^ 
0; 



wire Ie261f34f64899da2fbe8ceea78b5b4f0; 
assign Ie261f34f64899da2fbe8ceea78b5b4f0 = 
        y_nr_in[1] ^ 
        y_nr_in[51] ^ 
        y_nr_in[54] ^ 
        y_nr_in[178] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[138] = 
Ie261f34f64899da2fbe8ceea78b5b4f0 ^ 
0; 



wire I4adc3b50f0aa3586b3f78bf410a5ccfc; 
assign I4adc3b50f0aa3586b3f78bf410a5ccfc = 
        y_nr_in[2] ^ 
        y_nr_in[48] ^ 
        y_nr_in[55] ^ 
        y_nr_in[179] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[139] = 
I4adc3b50f0aa3586b3f78bf410a5ccfc ^ 
0; 



wire Ic3e50a904a86df001cf063d99e8436ca; 
assign Ic3e50a904a86df001cf063d99e8436ca = 
        y_nr_in[5] ^ 
        y_nr_in[20] ^ 
        y_nr_in[47] ^ 
        y_nr_in[180] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[140] = 
Ic3e50a904a86df001cf063d99e8436ca ^ 
0; 



wire Id91b187f81a3aa7914bc33fd2f3ea369; 
assign Id91b187f81a3aa7914bc33fd2f3ea369 = 
        y_nr_in[6] ^ 
        y_nr_in[21] ^ 
        y_nr_in[44] ^ 
        y_nr_in[181] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[141] = 
Id91b187f81a3aa7914bc33fd2f3ea369 ^ 
0; 



wire I9bce0668c89d26094a58fc55008293e0; 
assign I9bce0668c89d26094a58fc55008293e0 = 
        y_nr_in[7] ^ 
        y_nr_in[22] ^ 
        y_nr_in[45] ^ 
        y_nr_in[182] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[142] = 
I9bce0668c89d26094a58fc55008293e0 ^ 
0; 



wire Ia707df27cd9e632d430e530c71077452; 
assign Ia707df27cd9e632d430e530c71077452 = 
        y_nr_in[4] ^ 
        y_nr_in[23] ^ 
        y_nr_in[46] ^ 
        y_nr_in[183] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[143] = 
Ia707df27cd9e632d430e530c71077452 ^ 
0; 



wire I5a2bc1ba5f9d9062636fa7efaf27a615; 
assign I5a2bc1ba5f9d9062636fa7efaf27a615 = 
        y_nr_in[0] ^ 
        y_nr_in[10] ^ 
        y_nr_in[30] ^ 
        y_nr_in[184] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[144] = 
I5a2bc1ba5f9d9062636fa7efaf27a615 ^ 
0; 



wire Ibed44a0faea14928275cdbbda91f750e; 
assign Ibed44a0faea14928275cdbbda91f750e = 
        y_nr_in[1] ^ 
        y_nr_in[11] ^ 
        y_nr_in[31] ^ 
        y_nr_in[185] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[145] = 
Ibed44a0faea14928275cdbbda91f750e ^ 
0; 



wire I0ea35c7ecd2931f713239f6c18874ff7; 
assign I0ea35c7ecd2931f713239f6c18874ff7 = 
        y_nr_in[2] ^ 
        y_nr_in[8] ^ 
        y_nr_in[28] ^ 
        y_nr_in[186] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[146] = 
I0ea35c7ecd2931f713239f6c18874ff7 ^ 
0; 



wire If6b7aee9fd2617639a1b21a8efafd064; 
assign If6b7aee9fd2617639a1b21a8efafd064 = 
        y_nr_in[3] ^ 
        y_nr_in[9] ^ 
        y_nr_in[29] ^ 
        y_nr_in[187] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[147] = 
If6b7aee9fd2617639a1b21a8efafd064 ^ 
0; 



wire I1b52246a6bd429a323a690084ff1adbf; 
assign I1b52246a6bd429a323a690084ff1adbf = 
        y_nr_in[43] ^ 
        y_nr_in[55] ^ 
        y_nr_in[188] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[148] = 
I1b52246a6bd429a323a690084ff1adbf ^ 
0; 



wire I7f63e70637cc82703e7139451514fc34; 
assign I7f63e70637cc82703e7139451514fc34 = 
        y_nr_in[40] ^ 
        y_nr_in[52] ^ 
        y_nr_in[189] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[149] = 
I7f63e70637cc82703e7139451514fc34 ^ 
0; 



wire I9c55c7a8703858d14b92d362a121a529; 
assign I9c55c7a8703858d14b92d362a121a529 = 
        y_nr_in[41] ^ 
        y_nr_in[53] ^ 
        y_nr_in[190] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[150] = 
I9c55c7a8703858d14b92d362a121a529 ^ 
0; 



wire I73242a04195961520de17bb831a67340; 
assign I73242a04195961520de17bb831a67340 = 
        y_nr_in[42] ^ 
        y_nr_in[54] ^ 
        y_nr_in[191] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[151] = 
I73242a04195961520de17bb831a67340 ^ 
0; 



wire Ie9c09569e6b80fcbb527d196856a2311; 
assign Ie9c09569e6b80fcbb527d196856a2311 = 
        y_nr_in[7] ^ 
        y_nr_in[22] ^ 
        y_nr_in[46] ^ 
        y_nr_in[192] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[152] = 
Ie9c09569e6b80fcbb527d196856a2311 ^ 
0; 



wire Iace7382cabbec56b98dfbb7b74558d5a; 
assign Iace7382cabbec56b98dfbb7b74558d5a = 
        y_nr_in[4] ^ 
        y_nr_in[23] ^ 
        y_nr_in[47] ^ 
        y_nr_in[193] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[153] = 
Iace7382cabbec56b98dfbb7b74558d5a ^ 
0; 



wire I0c3eb9bb0a70fdbc1f4bd86ea5687afc; 
assign I0c3eb9bb0a70fdbc1f4bd86ea5687afc = 
        y_nr_in[5] ^ 
        y_nr_in[20] ^ 
        y_nr_in[44] ^ 
        y_nr_in[194] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[154] = 
I0c3eb9bb0a70fdbc1f4bd86ea5687afc ^ 
0; 



wire Iec5145499f910e94d8fea9af1b69b6fe; 
assign Iec5145499f910e94d8fea9af1b69b6fe = 
        y_nr_in[6] ^ 
        y_nr_in[21] ^ 
        y_nr_in[45] ^ 
        y_nr_in[195] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[155] = 
Iec5145499f910e94d8fea9af1b69b6fe ^ 
0; 



wire Iccd2984043aa17d5d5bd1bb142412c92; 
assign Iccd2984043aa17d5d5bd1bb142412c92 = 
        y_nr_in[3] ^ 
        y_nr_in[28] ^ 
        y_nr_in[50] ^ 
        y_nr_in[196] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[156] = 
Iccd2984043aa17d5d5bd1bb142412c92 ^ 
0; 



wire I9c615aa98d0ba18438612332a02f3b4f; 
assign I9c615aa98d0ba18438612332a02f3b4f = 
        y_nr_in[0] ^ 
        y_nr_in[29] ^ 
        y_nr_in[51] ^ 
        y_nr_in[197] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[157] = 
I9c615aa98d0ba18438612332a02f3b4f ^ 
0; 



wire I2d3103a2a93572b8cee6b5df58103c8b; 
assign I2d3103a2a93572b8cee6b5df58103c8b = 
        y_nr_in[1] ^ 
        y_nr_in[30] ^ 
        y_nr_in[48] ^ 
        y_nr_in[198] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[158] = 
I2d3103a2a93572b8cee6b5df58103c8b ^ 
0; 



wire Ic2e109b0711c2c271e6d5fb8bb9d5618; 
assign Ic2e109b0711c2c271e6d5fb8bb9d5618 = 
        y_nr_in[2] ^ 
        y_nr_in[31] ^ 
        y_nr_in[49] ^ 
        y_nr_in[199] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[159] = 
Ic2e109b0711c2c271e6d5fb8bb9d5618 ^ 
0; 



wire Id4121884b2a4dbae3ac5f125810c6fe3; 
assign Id4121884b2a4dbae3ac5f125810c6fe3 = 
        y_nr_in[8] ^ 
        y_nr_in[43] ^ 
        y_nr_in[52] ^ 
        y_nr_in[200] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[160] = 
Id4121884b2a4dbae3ac5f125810c6fe3 ^ 
0; 



wire Icf8e93bc13888b236df96d117d5d8a43; 
assign Icf8e93bc13888b236df96d117d5d8a43 = 
        y_nr_in[9] ^ 
        y_nr_in[40] ^ 
        y_nr_in[53] ^ 
        y_nr_in[201] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[161] = 
Icf8e93bc13888b236df96d117d5d8a43 ^ 
0; 



wire If44976055a3682505dfa69367e519577; 
assign If44976055a3682505dfa69367e519577 = 
        y_nr_in[10] ^ 
        y_nr_in[41] ^ 
        y_nr_in[54] ^ 
        y_nr_in[202] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[162] = 
If44976055a3682505dfa69367e519577 ^ 
0; 



wire Id41eef9050d65e401f1ae40027ce52d2; 
assign Id41eef9050d65e401f1ae40027ce52d2 = 
        y_nr_in[11] ^ 
        y_nr_in[42] ^ 
        y_nr_in[55] ^ 
        y_nr_in[203] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[163] = 
Id41eef9050d65e401f1ae40027ce52d2 ^ 
0; 



wire Ia571e9d90d1840625dda701118990ff0; 
assign Ia571e9d90d1840625dda701118990ff0 = 
        y_nr_in[5] ^ 
        y_nr_in[21] ^ 
        y_nr_in[46] ^ 
        y_nr_in[204] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[164] = 
Ia571e9d90d1840625dda701118990ff0 ^ 
0; 



wire Ieaaf8a003c240b7649420f309bd36445; 
assign Ieaaf8a003c240b7649420f309bd36445 = 
        y_nr_in[6] ^ 
        y_nr_in[22] ^ 
        y_nr_in[47] ^ 
        y_nr_in[205] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[165] = 
Ieaaf8a003c240b7649420f309bd36445 ^ 
0; 



wire I102e12bfca09b1adbb0a4098432726e2; 
assign I102e12bfca09b1adbb0a4098432726e2 = 
        y_nr_in[7] ^ 
        y_nr_in[23] ^ 
        y_nr_in[44] ^ 
        y_nr_in[206] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[166] = 
I102e12bfca09b1adbb0a4098432726e2 ^ 
0; 



wire I98f435952752e1e6a9c7f0909227fdac; 
assign I98f435952752e1e6a9c7f0909227fdac = 
        y_nr_in[4] ^ 
        y_nr_in[20] ^ 
        y_nr_in[45] ^ 
        y_nr_in[207] ^ 
0; 



assign Icab1e6ce3154e84b7ea0d3d9c82bcdc1[167] = 
I98f435952752e1e6a9c7f0909227fdac ^ 
0; 



