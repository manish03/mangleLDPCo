//`include "GF2_LDPC_flogtanh_0x00012_assign_inc.sv"
//always_comb begin
              Ia9be81772a42d1908d7f14f7ec313644['h00000] = 
          (!flogtanh_sel['h00012]) ? 
                       Ic7e91188980d728ad34dbe693d9a6e04['h00000] : //%
                       Ic7e91188980d728ad34dbe693d9a6e04['h00001] ;
//end
