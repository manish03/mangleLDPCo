//`include "GF2_LDPC_flogtanh_0x0000a_assign_inc.sv"
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00000] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h00000] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h00001] ;
//end
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00001] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h00002] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h00003] ;
//end
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00002] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h00004] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h00005] ;
//end
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00003] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h00006] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h00007] ;
//end
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00004] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h00008] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h00009] ;
//end
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00005] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h0000a] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h0000b] ;
//end
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00006] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h0000c] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h0000d] ;
//end
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00007] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h0000e] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h0000f] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00008] =  I986ccea2f9226242e2772b9c3af42d87['h00010] ;
//end
//always_comb begin
              I1a62004aa5608ddf7a551106f9a8a7ac['h00009] = 
          (!flogtanh_sel['h0000a]) ? 
                       I986ccea2f9226242e2772b9c3af42d87['h00012] : //%
                       I986ccea2f9226242e2772b9c3af42d87['h00013] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0000a] =  I986ccea2f9226242e2772b9c3af42d87['h00014] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0000b] =  I986ccea2f9226242e2772b9c3af42d87['h00016] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0000c] =  I986ccea2f9226242e2772b9c3af42d87['h00018] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0000d] =  I986ccea2f9226242e2772b9c3af42d87['h0001a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0000e] =  I986ccea2f9226242e2772b9c3af42d87['h0001c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0000f] =  I986ccea2f9226242e2772b9c3af42d87['h0001e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00010] =  I986ccea2f9226242e2772b9c3af42d87['h00020] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00011] =  I986ccea2f9226242e2772b9c3af42d87['h00022] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00012] =  I986ccea2f9226242e2772b9c3af42d87['h00024] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00013] =  I986ccea2f9226242e2772b9c3af42d87['h00026] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00014] =  I986ccea2f9226242e2772b9c3af42d87['h00028] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00015] =  I986ccea2f9226242e2772b9c3af42d87['h0002a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00016] =  I986ccea2f9226242e2772b9c3af42d87['h0002c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00017] =  I986ccea2f9226242e2772b9c3af42d87['h0002e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00018] =  I986ccea2f9226242e2772b9c3af42d87['h00030] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00019] =  I986ccea2f9226242e2772b9c3af42d87['h00032] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0001a] =  I986ccea2f9226242e2772b9c3af42d87['h00034] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0001b] =  I986ccea2f9226242e2772b9c3af42d87['h00036] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0001c] =  I986ccea2f9226242e2772b9c3af42d87['h00038] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0001d] =  I986ccea2f9226242e2772b9c3af42d87['h0003a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0001e] =  I986ccea2f9226242e2772b9c3af42d87['h0003c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0001f] =  I986ccea2f9226242e2772b9c3af42d87['h0003e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00020] =  I986ccea2f9226242e2772b9c3af42d87['h00040] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00021] =  I986ccea2f9226242e2772b9c3af42d87['h00042] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00022] =  I986ccea2f9226242e2772b9c3af42d87['h00044] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00023] =  I986ccea2f9226242e2772b9c3af42d87['h00046] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00024] =  I986ccea2f9226242e2772b9c3af42d87['h00048] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00025] =  I986ccea2f9226242e2772b9c3af42d87['h0004a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00026] =  I986ccea2f9226242e2772b9c3af42d87['h0004c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00027] =  I986ccea2f9226242e2772b9c3af42d87['h0004e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00028] =  I986ccea2f9226242e2772b9c3af42d87['h00050] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00029] =  I986ccea2f9226242e2772b9c3af42d87['h00052] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0002a] =  I986ccea2f9226242e2772b9c3af42d87['h00054] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0002b] =  I986ccea2f9226242e2772b9c3af42d87['h00056] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0002c] =  I986ccea2f9226242e2772b9c3af42d87['h00058] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0002d] =  I986ccea2f9226242e2772b9c3af42d87['h0005a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0002e] =  I986ccea2f9226242e2772b9c3af42d87['h0005c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0002f] =  I986ccea2f9226242e2772b9c3af42d87['h0005e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00030] =  I986ccea2f9226242e2772b9c3af42d87['h00060] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00031] =  I986ccea2f9226242e2772b9c3af42d87['h00062] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00032] =  I986ccea2f9226242e2772b9c3af42d87['h00064] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00033] =  I986ccea2f9226242e2772b9c3af42d87['h00066] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00034] =  I986ccea2f9226242e2772b9c3af42d87['h00068] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00035] =  I986ccea2f9226242e2772b9c3af42d87['h0006a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00036] =  I986ccea2f9226242e2772b9c3af42d87['h0006c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00037] =  I986ccea2f9226242e2772b9c3af42d87['h0006e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00038] =  I986ccea2f9226242e2772b9c3af42d87['h00070] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00039] =  I986ccea2f9226242e2772b9c3af42d87['h00072] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0003a] =  I986ccea2f9226242e2772b9c3af42d87['h00074] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0003b] =  I986ccea2f9226242e2772b9c3af42d87['h00076] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0003c] =  I986ccea2f9226242e2772b9c3af42d87['h00078] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0003d] =  I986ccea2f9226242e2772b9c3af42d87['h0007a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0003e] =  I986ccea2f9226242e2772b9c3af42d87['h0007c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0003f] =  I986ccea2f9226242e2772b9c3af42d87['h0007e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00040] =  I986ccea2f9226242e2772b9c3af42d87['h00080] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00041] =  I986ccea2f9226242e2772b9c3af42d87['h00082] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00042] =  I986ccea2f9226242e2772b9c3af42d87['h00084] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00043] =  I986ccea2f9226242e2772b9c3af42d87['h00086] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00044] =  I986ccea2f9226242e2772b9c3af42d87['h00088] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00045] =  I986ccea2f9226242e2772b9c3af42d87['h0008a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00046] =  I986ccea2f9226242e2772b9c3af42d87['h0008c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00047] =  I986ccea2f9226242e2772b9c3af42d87['h0008e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00048] =  I986ccea2f9226242e2772b9c3af42d87['h00090] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00049] =  I986ccea2f9226242e2772b9c3af42d87['h00092] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0004a] =  I986ccea2f9226242e2772b9c3af42d87['h00094] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0004b] =  I986ccea2f9226242e2772b9c3af42d87['h00096] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0004c] =  I986ccea2f9226242e2772b9c3af42d87['h00098] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0004d] =  I986ccea2f9226242e2772b9c3af42d87['h0009a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0004e] =  I986ccea2f9226242e2772b9c3af42d87['h0009c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0004f] =  I986ccea2f9226242e2772b9c3af42d87['h0009e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00050] =  I986ccea2f9226242e2772b9c3af42d87['h000a0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00051] =  I986ccea2f9226242e2772b9c3af42d87['h000a2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00052] =  I986ccea2f9226242e2772b9c3af42d87['h000a4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00053] =  I986ccea2f9226242e2772b9c3af42d87['h000a6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00054] =  I986ccea2f9226242e2772b9c3af42d87['h000a8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00055] =  I986ccea2f9226242e2772b9c3af42d87['h000aa] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00056] =  I986ccea2f9226242e2772b9c3af42d87['h000ac] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00057] =  I986ccea2f9226242e2772b9c3af42d87['h000ae] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00058] =  I986ccea2f9226242e2772b9c3af42d87['h000b0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00059] =  I986ccea2f9226242e2772b9c3af42d87['h000b2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0005a] =  I986ccea2f9226242e2772b9c3af42d87['h000b4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0005b] =  I986ccea2f9226242e2772b9c3af42d87['h000b6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0005c] =  I986ccea2f9226242e2772b9c3af42d87['h000b8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0005d] =  I986ccea2f9226242e2772b9c3af42d87['h000ba] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0005e] =  I986ccea2f9226242e2772b9c3af42d87['h000bc] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0005f] =  I986ccea2f9226242e2772b9c3af42d87['h000be] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00060] =  I986ccea2f9226242e2772b9c3af42d87['h000c0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00061] =  I986ccea2f9226242e2772b9c3af42d87['h000c2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00062] =  I986ccea2f9226242e2772b9c3af42d87['h000c4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00063] =  I986ccea2f9226242e2772b9c3af42d87['h000c6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00064] =  I986ccea2f9226242e2772b9c3af42d87['h000c8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00065] =  I986ccea2f9226242e2772b9c3af42d87['h000ca] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00066] =  I986ccea2f9226242e2772b9c3af42d87['h000cc] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00067] =  I986ccea2f9226242e2772b9c3af42d87['h000ce] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00068] =  I986ccea2f9226242e2772b9c3af42d87['h000d0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00069] =  I986ccea2f9226242e2772b9c3af42d87['h000d2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0006a] =  I986ccea2f9226242e2772b9c3af42d87['h000d4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0006b] =  I986ccea2f9226242e2772b9c3af42d87['h000d6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0006c] =  I986ccea2f9226242e2772b9c3af42d87['h000d8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0006d] =  I986ccea2f9226242e2772b9c3af42d87['h000da] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0006e] =  I986ccea2f9226242e2772b9c3af42d87['h000dc] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0006f] =  I986ccea2f9226242e2772b9c3af42d87['h000de] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00070] =  I986ccea2f9226242e2772b9c3af42d87['h000e0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00071] =  I986ccea2f9226242e2772b9c3af42d87['h000e2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00072] =  I986ccea2f9226242e2772b9c3af42d87['h000e4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00073] =  I986ccea2f9226242e2772b9c3af42d87['h000e6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00074] =  I986ccea2f9226242e2772b9c3af42d87['h000e8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00075] =  I986ccea2f9226242e2772b9c3af42d87['h000ea] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00076] =  I986ccea2f9226242e2772b9c3af42d87['h000ec] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00077] =  I986ccea2f9226242e2772b9c3af42d87['h000ee] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00078] =  I986ccea2f9226242e2772b9c3af42d87['h000f0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00079] =  I986ccea2f9226242e2772b9c3af42d87['h000f2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0007a] =  I986ccea2f9226242e2772b9c3af42d87['h000f4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0007b] =  I986ccea2f9226242e2772b9c3af42d87['h000f6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0007c] =  I986ccea2f9226242e2772b9c3af42d87['h000f8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0007d] =  I986ccea2f9226242e2772b9c3af42d87['h000fa] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0007e] =  I986ccea2f9226242e2772b9c3af42d87['h000fc] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0007f] =  I986ccea2f9226242e2772b9c3af42d87['h000fe] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00080] =  I986ccea2f9226242e2772b9c3af42d87['h00100] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00081] =  I986ccea2f9226242e2772b9c3af42d87['h00102] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00082] =  I986ccea2f9226242e2772b9c3af42d87['h00104] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00083] =  I986ccea2f9226242e2772b9c3af42d87['h00106] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00084] =  I986ccea2f9226242e2772b9c3af42d87['h00108] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00085] =  I986ccea2f9226242e2772b9c3af42d87['h0010a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00086] =  I986ccea2f9226242e2772b9c3af42d87['h0010c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00087] =  I986ccea2f9226242e2772b9c3af42d87['h0010e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00088] =  I986ccea2f9226242e2772b9c3af42d87['h00110] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00089] =  I986ccea2f9226242e2772b9c3af42d87['h00112] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0008a] =  I986ccea2f9226242e2772b9c3af42d87['h00114] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0008b] =  I986ccea2f9226242e2772b9c3af42d87['h00116] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0008c] =  I986ccea2f9226242e2772b9c3af42d87['h00118] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0008d] =  I986ccea2f9226242e2772b9c3af42d87['h0011a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0008e] =  I986ccea2f9226242e2772b9c3af42d87['h0011c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0008f] =  I986ccea2f9226242e2772b9c3af42d87['h0011e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00090] =  I986ccea2f9226242e2772b9c3af42d87['h00120] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00091] =  I986ccea2f9226242e2772b9c3af42d87['h00122] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00092] =  I986ccea2f9226242e2772b9c3af42d87['h00124] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00093] =  I986ccea2f9226242e2772b9c3af42d87['h00126] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00094] =  I986ccea2f9226242e2772b9c3af42d87['h00128] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00095] =  I986ccea2f9226242e2772b9c3af42d87['h0012a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00096] =  I986ccea2f9226242e2772b9c3af42d87['h0012c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00097] =  I986ccea2f9226242e2772b9c3af42d87['h0012e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00098] =  I986ccea2f9226242e2772b9c3af42d87['h00130] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h00099] =  I986ccea2f9226242e2772b9c3af42d87['h00132] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0009a] =  I986ccea2f9226242e2772b9c3af42d87['h00134] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0009b] =  I986ccea2f9226242e2772b9c3af42d87['h00136] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0009c] =  I986ccea2f9226242e2772b9c3af42d87['h00138] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0009d] =  I986ccea2f9226242e2772b9c3af42d87['h0013a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0009e] =  I986ccea2f9226242e2772b9c3af42d87['h0013c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h0009f] =  I986ccea2f9226242e2772b9c3af42d87['h0013e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a0] =  I986ccea2f9226242e2772b9c3af42d87['h00140] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a1] =  I986ccea2f9226242e2772b9c3af42d87['h00142] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a2] =  I986ccea2f9226242e2772b9c3af42d87['h00144] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a3] =  I986ccea2f9226242e2772b9c3af42d87['h00146] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a4] =  I986ccea2f9226242e2772b9c3af42d87['h00148] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a5] =  I986ccea2f9226242e2772b9c3af42d87['h0014a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a6] =  I986ccea2f9226242e2772b9c3af42d87['h0014c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a7] =  I986ccea2f9226242e2772b9c3af42d87['h0014e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a8] =  I986ccea2f9226242e2772b9c3af42d87['h00150] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000a9] =  I986ccea2f9226242e2772b9c3af42d87['h00152] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000aa] =  I986ccea2f9226242e2772b9c3af42d87['h00154] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ab] =  I986ccea2f9226242e2772b9c3af42d87['h00156] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ac] =  I986ccea2f9226242e2772b9c3af42d87['h00158] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ad] =  I986ccea2f9226242e2772b9c3af42d87['h0015a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ae] =  I986ccea2f9226242e2772b9c3af42d87['h0015c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000af] =  I986ccea2f9226242e2772b9c3af42d87['h0015e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b0] =  I986ccea2f9226242e2772b9c3af42d87['h00160] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b1] =  I986ccea2f9226242e2772b9c3af42d87['h00162] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b2] =  I986ccea2f9226242e2772b9c3af42d87['h00164] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b3] =  I986ccea2f9226242e2772b9c3af42d87['h00166] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b4] =  I986ccea2f9226242e2772b9c3af42d87['h00168] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b5] =  I986ccea2f9226242e2772b9c3af42d87['h0016a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b6] =  I986ccea2f9226242e2772b9c3af42d87['h0016c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b7] =  I986ccea2f9226242e2772b9c3af42d87['h0016e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b8] =  I986ccea2f9226242e2772b9c3af42d87['h00170] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000b9] =  I986ccea2f9226242e2772b9c3af42d87['h00172] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ba] =  I986ccea2f9226242e2772b9c3af42d87['h00174] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000bb] =  I986ccea2f9226242e2772b9c3af42d87['h00176] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000bc] =  I986ccea2f9226242e2772b9c3af42d87['h00178] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000bd] =  I986ccea2f9226242e2772b9c3af42d87['h0017a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000be] =  I986ccea2f9226242e2772b9c3af42d87['h0017c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000bf] =  I986ccea2f9226242e2772b9c3af42d87['h0017e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c0] =  I986ccea2f9226242e2772b9c3af42d87['h00180] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c1] =  I986ccea2f9226242e2772b9c3af42d87['h00182] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c2] =  I986ccea2f9226242e2772b9c3af42d87['h00184] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c3] =  I986ccea2f9226242e2772b9c3af42d87['h00186] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c4] =  I986ccea2f9226242e2772b9c3af42d87['h00188] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c5] =  I986ccea2f9226242e2772b9c3af42d87['h0018a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c6] =  I986ccea2f9226242e2772b9c3af42d87['h0018c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c7] =  I986ccea2f9226242e2772b9c3af42d87['h0018e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c8] =  I986ccea2f9226242e2772b9c3af42d87['h00190] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000c9] =  I986ccea2f9226242e2772b9c3af42d87['h00192] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ca] =  I986ccea2f9226242e2772b9c3af42d87['h00194] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000cb] =  I986ccea2f9226242e2772b9c3af42d87['h00196] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000cc] =  I986ccea2f9226242e2772b9c3af42d87['h00198] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000cd] =  I986ccea2f9226242e2772b9c3af42d87['h0019a] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ce] =  I986ccea2f9226242e2772b9c3af42d87['h0019c] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000cf] =  I986ccea2f9226242e2772b9c3af42d87['h0019e] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d0] =  I986ccea2f9226242e2772b9c3af42d87['h001a0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d1] =  I986ccea2f9226242e2772b9c3af42d87['h001a2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d2] =  I986ccea2f9226242e2772b9c3af42d87['h001a4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d3] =  I986ccea2f9226242e2772b9c3af42d87['h001a6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d4] =  I986ccea2f9226242e2772b9c3af42d87['h001a8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d5] =  I986ccea2f9226242e2772b9c3af42d87['h001aa] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d6] =  I986ccea2f9226242e2772b9c3af42d87['h001ac] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d7] =  I986ccea2f9226242e2772b9c3af42d87['h001ae] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d8] =  I986ccea2f9226242e2772b9c3af42d87['h001b0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000d9] =  I986ccea2f9226242e2772b9c3af42d87['h001b2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000da] =  I986ccea2f9226242e2772b9c3af42d87['h001b4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000db] =  I986ccea2f9226242e2772b9c3af42d87['h001b6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000dc] =  I986ccea2f9226242e2772b9c3af42d87['h001b8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000dd] =  I986ccea2f9226242e2772b9c3af42d87['h001ba] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000de] =  I986ccea2f9226242e2772b9c3af42d87['h001bc] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000df] =  I986ccea2f9226242e2772b9c3af42d87['h001be] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e0] =  I986ccea2f9226242e2772b9c3af42d87['h001c0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e1] =  I986ccea2f9226242e2772b9c3af42d87['h001c2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e2] =  I986ccea2f9226242e2772b9c3af42d87['h001c4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e3] =  I986ccea2f9226242e2772b9c3af42d87['h001c6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e4] =  I986ccea2f9226242e2772b9c3af42d87['h001c8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e5] =  I986ccea2f9226242e2772b9c3af42d87['h001ca] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e6] =  I986ccea2f9226242e2772b9c3af42d87['h001cc] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e7] =  I986ccea2f9226242e2772b9c3af42d87['h001ce] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e8] =  I986ccea2f9226242e2772b9c3af42d87['h001d0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000e9] =  I986ccea2f9226242e2772b9c3af42d87['h001d2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ea] =  I986ccea2f9226242e2772b9c3af42d87['h001d4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000eb] =  I986ccea2f9226242e2772b9c3af42d87['h001d6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ec] =  I986ccea2f9226242e2772b9c3af42d87['h001d8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ed] =  I986ccea2f9226242e2772b9c3af42d87['h001da] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ee] =  I986ccea2f9226242e2772b9c3af42d87['h001dc] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ef] =  I986ccea2f9226242e2772b9c3af42d87['h001de] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f0] =  I986ccea2f9226242e2772b9c3af42d87['h001e0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f1] =  I986ccea2f9226242e2772b9c3af42d87['h001e2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f2] =  I986ccea2f9226242e2772b9c3af42d87['h001e4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f3] =  I986ccea2f9226242e2772b9c3af42d87['h001e6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f4] =  I986ccea2f9226242e2772b9c3af42d87['h001e8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f5] =  I986ccea2f9226242e2772b9c3af42d87['h001ea] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f6] =  I986ccea2f9226242e2772b9c3af42d87['h001ec] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f7] =  I986ccea2f9226242e2772b9c3af42d87['h001ee] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f8] =  I986ccea2f9226242e2772b9c3af42d87['h001f0] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000f9] =  I986ccea2f9226242e2772b9c3af42d87['h001f2] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000fa] =  I986ccea2f9226242e2772b9c3af42d87['h001f4] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000fb] =  I986ccea2f9226242e2772b9c3af42d87['h001f6] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000fc] =  I986ccea2f9226242e2772b9c3af42d87['h001f8] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000fd] =  I986ccea2f9226242e2772b9c3af42d87['h001fa] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000fe] =  I986ccea2f9226242e2772b9c3af42d87['h001fc] ;
//end
//always_comb begin // 
               I1a62004aa5608ddf7a551106f9a8a7ac['h000ff] =  I986ccea2f9226242e2772b9c3af42d87['h001fe] ;
//end
