              I9c9ab24ecd80ca61b89534e3e5adfca8 = 
          (!fgallag_sel[0]) ? 
                       I53846946a877f30f72076ee6f633a0e5: 
                       I5d219e3294f2763bc17209a55758ab54;
              Ie92d645c17dda47f594bc34b0937caac = 
          (!fgallag_sel[0]) ? 
                       I6273ee09aacad20f733530af1a987ff3: 
                       Ie0f63a67c0a6ec07e7bcb943e7804f9a;
              Ieb8b25a5f6d3cc4cead3f3845234d1d3 = 
          (!fgallag_sel[0]) ? 
                       I7b83ef4e45fe20e023e08aa3e56bb21e: 
                       Ibc8f334cefc147e5c58e7542d26fbe2b;
              Ibcbdbe8034a373448800d1b745cb5849 = 
          (!fgallag_sel[0]) ? 
                       I662a566f576ee431bced6f852294713e: 
                       I2a4bc966b71864a79f582727f122ab60;
              Ibd0769c69670150d8263d9873cbf668f = 
          (!fgallag_sel[0]) ? 
                       I23d9f47edf51ff1c2a6275531a1f66be: 
                       Id46ae2d16f43af3529d91eb4d6bd098e;
              I2010cff1e77f9706d8c659482f51c898 = 
          (!fgallag_sel[0]) ? 
                       I51298122656d9b893c1dbb33a281f134: 
                       I22e0a22ed1768671dbe3caef8ac499cb;
              I4183447a1a1727e91b0fcabb9bec1963 = 
          (!fgallag_sel[0]) ? 
                       Ifb9327c663379f77471d460eced9c1b7: 
                       Id6080749dda3cd29c1ce36ab39759709;
              I780bea956f609c6f3cd0ffd126f99316 = 
          (!fgallag_sel[0]) ? 
                       I532fd8f9065e524727e276a1a8408008: 
                       I1f0b23c673ff55115f55c80a970172fc;
              I349cff38817dd1607e798b9a2ae6fb8b = 
          (!fgallag_sel[0]) ? 
                       I9f99ad4587fb6907b3804c11125f738f: 
                       I719bd7e94d4289c6fd59bb91ee559980;
              I3ff605a8af8eceb2c055e842e6208958 = 
          (!fgallag_sel[0]) ? 
                       I9103b57e3550cb68266ba8b102e50dfd: 
                       I89fca1c1832813b84cafe145377d7b5e;
              Ib53b2b0d39dbe6d09f51e0af27e5986f = 
          (!fgallag_sel[0]) ? 
                       Ie17de6e388779502a143212813a50317: 
                       Ifcc046128364b8da7bc3d9ddab96a061;
              I343242367c13febc05ee63f57dd4f754 = 
          (!fgallag_sel[0]) ? 
                       Iabe4b7a23f682ed62162dfde9e15d6cf: 
                       I734eaef0b7d7f6ae5d668ac9b374ff51;
              Ibde6749f31c571c5209a8b36c1c8f4da = 
          (!fgallag_sel[0]) ? 
                       I0e0e9fdfeb3e2115deb903b973217384: 
                       Ibfd2fd7aa2426054706d0c4e4c0a7cba;
              Ib735324969bc744cc0ab8c2b3a7c5561 = 
          (!fgallag_sel[0]) ? 
                       I0906247e3ba96971232bc42185c9a9b8: 
                       Ia3908fda391d7caf1b479d9655164c30;
              If53ed28774233bca87090e799465e3a5 = 
          (!fgallag_sel[0]) ? 
                       I820e95cdc583108195e8dd0e2d1f4b7f: 
                       Ibdf5c2c57269da1b04748a59802c8e2a;
              Ib5017be08e079fe946c365fc01461d11 = 
          (!fgallag_sel[0]) ? 
                       Idd85c8c853438679d99bed4d0ba46af7: 
                       I4d617d0b669b3ff1b08dcd4b7440af33;
              I0f24b1ca1d272d4971cde83a2acfe5ac = 
          (!fgallag_sel[0]) ? 
                       I60d579b60b02f9fc14e98d7d0eb54c18: 
                       Ic1a37750fc3d7eb08ad649de157f45a9;
              I1d1f2f5dd46b3f89c5a614ebad298d13 = 
          (!fgallag_sel[0]) ? 
                       I0c13ec63e7208b35a1d4511e1da29fa3: 
                       If10c9545a713996735934c5f15cf5365;
              I09dbcf2140141aaa400ad52408f8ab41 = 
          (!fgallag_sel[0]) ? 
                       Ic475963164a956dd24ede91e9d61003d: 
                       I42001c4b6ab9fb03489ca25defb6c222;
              I8315726dd19b5074a78796ee704d7108 = 
          (!fgallag_sel[0]) ? 
                       Idcfb16adf2996c8cb51e402daafd1734: 
                       I924108a2723afd07735574a6f4ebe671;
              Idb03654ee570200d2fe82907af7095d7 = 
          (!fgallag_sel[0]) ? 
                       If9fd9ae380997e75ebed2ddd3f93e76f: 
                       Ief876b7b2af1fbed4d3f457cdb46e0d9;
              I9a5f25915425b586c1c3979240ff1a54 = 
          (!fgallag_sel[0]) ? 
                       Id2bd196ca25e1a077fb2a9207f143c01: 
                       I926e2a038d48db29b5ce215cd6cf6a04;
              I259241ceeda0568e6c10162cd43ca1dc = 
          (!fgallag_sel[0]) ? 
                       I4ba2cfd94590dee1723ce63afd0926ab: 
                       I0d42326464ae4c3a55038e0343cebf5a;
              I66d1b07d77d2fe21d535920b30e176ff = 
          (!fgallag_sel[0]) ? 
                       If05fde321fd1456422550f5c3903b826: 
                       I41ec48a5a1d657a6266b8f845550d0c2;
              I135dcccb8e63f697fe4559b964322345 = 
          (!fgallag_sel[0]) ? 
                       I76473b4885d423029324fe74ed13d6ed: 
                       I8ef2366947e3f1352f3874e4ac58d7b2;
              Ic37c4058485edfc0ca4f12fd7a97bf93 = 
          (!fgallag_sel[0]) ? 
                       I874c1e455f85e617a5032ec230fdfdc5: 
                       I16d6b6b19890a6bbdf15ddc27717aa30;
              I1400488e51bbe6c921439713342d39f8 = 
          (!fgallag_sel[0]) ? 
                       I6af6d04126eec9eb91e5653cc95c9ef3: 
                       If501a668f24fd62a69d0e3c253739c79;
              Iaa8359974e7a41f754b38d6a232c5e72 = 
          (!fgallag_sel[0]) ? 
                       I9b70e215a2a1578811b40c669826d41a: 
                       I26d82966efbe51e03edcd66a5a507ebb;
              Ie99b9c10b4b5208374b9f4ba1bd3eeab = 
          (!fgallag_sel[0]) ? 
                       I2e4afb94e4af76b4e3d859815bb338fb: 
                       Ie19faf5d037b74974102c386a13f4946;
              I54462091230adebf4bf4ec0cea25e374 = 
          (!fgallag_sel[0]) ? 
                       I2d56338af0755ae5c4ef71ddad3112b1: 
                       I99ab212db901b0e65eb33be27c46bd19;
              Iba9e737dd791a2ee966dbf6958339d65 = 
          (!fgallag_sel[0]) ? 
                       If8c09c14d78b1deaf76df6f4de910c64: 
                       I1b0ccac0f5cc741403fd6e680899f96f;
               Ib205f5f9a6005baa465f1b254e4014d0 =  I38153cd88e8b2452977d7dc9b9f44a74 ;
              I5ea13e282884d2343e8fdbe17d7ee058 = 
          (!fgallag_sel[0]) ? 
                       Ic10eb104fe38a176a51507e748406958: 
                       I979fd1b01c99b76a4ff2d0abfb0c2ae9;
              I6d8ed091d5f44b3b49e8b0eb63f0d106 = 
          (!fgallag_sel[0]) ? 
                       Ibe530a86c501fbc8dba64ed24806bdf4: 
                       If03531315c68272f7de2b0e969770f48;
               I4109473d968250506e17f8227bc55d06 =  I20160f4e380b0920bcb30a0321b7bfa8 ;
              Ia7da78b0d37028fcd34d3d39c7e36596 = 
          (!fgallag_sel[0]) ? 
                       I70f4396800d2cb065ad5fe655bacbfd0: 
                       If27a0187d1188cf7a8aba100a90cb069;
               I034454a1608fbde69fffb6b28e685f9f =  I8994866d080b1befe414fea347e7e74a ;
              I6e487d671a19855fd1eae42664d9c57f = 
          (!fgallag_sel[0]) ? 
                       I8730924fec54ffaa78a0ffea7e8386ba: 
                       I338fb9183219691c6b50e6a824fcb14c;
              Ib49b6b6895bd7200dc9e026584bea017 = 
          (!fgallag_sel[0]) ? 
                       I1a3d82eaf2fc9235163c0a50765f4ef5: 
                       I922539f8d9ffc119ed3a5c92a21f149e;
               I220ce4284bf6adf0e46cf524b04a0e1b =  I3bc0f1eaad327d5990adb826e54c6d2f ;
              I64586e3b7241a57c2e887b651819c7f9 = 
          (!fgallag_sel[0]) ? 
                       I2e0ae02d7a3cdfa36e8645cc7dd0bce6: 
                       If2c59f326f3658dee0fd3b048af14cb7;
              Ifad0bf7a3d7d334b5f8ea0d1a973fd39 = 
          (!fgallag_sel[0]) ? 
                       I04431bd4be4601d3cb700c0cd6d9fd24: 
                       I7a6fe8c804087a19e32e760f50e3edfa;
              If060b99963382d16c1f779faf00a7128 = 
          (!fgallag_sel[0]) ? 
                       I979817e250e46dcc05f8a6690c2380f9: 
                       I3bbb836eee6b5e10fe55879f8620b888;
               Ie80ad5b1c3c4046c80e6cb96ee51e5c0 =  I8bc5128382cbffa289caec56f9b4a3f3 ;
               I4fe400daeacdfbebafcdf7e753af2787 =  I4ea5b39ed827d8d4618bcfd9283dfa83 ;
               I5c1ec1001d1ea61ab7198336742ed99d =  I0653a9ef861e5d8af22d120172c2dc03 ;
               If50cfdca6c9b8000665da2513244ff24 =  I1583cdcd13120f953691a5a60ee72b11 ;
               I4367feaf57687befa18bc6a902573bb9 =  I9bd98a9d18ce7c07e85287f6b80bfd31 ;
               I8f2820928683d8d88d41b80a9d9832dd =  I11f2e4eafc706b43c10a26edc8567052 ;
               Id980002a738b3ab2a4c2ccb9d232d141 =  I75705fa2cc0ac0577570501510e4e0fc ;
               Ib1db1798d076dc0a6fa322c47e0ac062 =  I8cefcac1f7fa2df45bb8a2f3d64f99c3 ;
              Iba73f7b76a2e16d7d84cfbab4473143d = 
          (!fgallag_sel[0]) ? 
                       I71a33ca1c7d18d5089d08a8476c8baf7: 
                       Ic85b012b9fa77becd419cac0f3692aed;
              Iad0a6e20283bbf4bd4114a0c70c0685e = 
          (!fgallag_sel[0]) ? 
                       I0ae9b4ca5ebb5f3d2e8b02884069e4e7: 
                       Ief312304eec0415d1ab208ed6726dd12;
              Ic772211084626d2ed3ddc4f32b467c6c = 
          (!fgallag_sel[0]) ? 
                       Icb9ebf1f5becaede273da59f466506ac: 
                       I465b9607a8dad0f1c499318d04f42aea;
               Ifcba38a9a6ca0931ba9d86396f257929 =  I2523c109974807b3b1c0f4b34693e255 ;
               I3ae9dbf37dbadabaf8a56188eae40288 =  Ibfb66b89c59008f3d4497ee16dad6712 ;
              Iae4d59e569911a81bb653cdb58c65137 = 
          (!fgallag_sel[0]) ? 
                       I489d1b46970800e9684c68b439c15be1: 
                       I835143e23243f3fd25cc1ab0ba5c123a;
               I9b12cb33d0f37813bd735c14d8be517e =  I028ef05ea84be3bc45c518f4f45653d2 ;
               Ifab01268c2a1f0385dc4b18a9d488321 =  If5a85945ad1f8d9bdc9213c5ae2c890f ;
              Ie0f0a8cf008e6a10d1698c11c380df97 = 
          (!fgallag_sel[0]) ? 
                       Ie703b5f1eeedaaaddf56ded14b1765bc: 
                       I21f34fbc269f5424ea30334ff7ab54f5;
               I99aa62ad841c5bd5b1f2b6758d046784 =  I07b47fce56edeb30319038e3a093efd7 ;
               I3fc64e5c431cd64d48f3cc5c9c86f342 =  Iee1b23b99f7de56829706633297a0513 ;
              I65a139ae2fa69f57c3a8ed35e00e29ae = 
          (!fgallag_sel[0]) ? 
                       Ifd5fcb1552fb372ae203fd0166d3df2c: 
                       Ibb2fb63aef1d336dfa829cd5ab3675b7;
               I628bc7c30b5e896c2b8f4af752b44637 =  I1672371cf33b259cf87210cc49aa35c8 ;
              I5c7ed27126a8097481ab5f966867783b = 
          (!fgallag_sel[0]) ? 
                       I2372d0a72998f0630e994aa3e1c20ff4: 
                       I8e363e0bd65cae9725cdd70e46778fee;
               I686481757183441e45d85fece1a7b514 =  Id6af962a16ff79ac6e9da3b4518b80b2 ;
               I10929316643f6670bedc63e77b293c97 =  I693f2c9a5d4da90c3105876991c4f4ba ;
               Ia66d818d01365175f416a4de87a281bb =  Id6561e53aa8f9fd116159969afaa20ae ;
               I7711386635a1760e7976d0947e0a5f8a =  I567872d8892064b62caeb3dcdc39e89c ;
               I4b2cc8ae58d2fb89bd9095b2bb688cbe =  Ia4e5d30bc160c1f72c8f39cdcd13e5a4 ;
               Ied1035a697824a18281435fe2b7f1f56 =  Ifdd13523ba0ce3329e3aca49a0a36385 ;
               I3e9ecaf8da044766c57685a1065ce10a =  I134d223e71b68cc9c76379f1368fb0f1 ;
              Ibebda2f9816088ea15cd5b4f555c5d33 = 
          (!fgallag_sel[0]) ? 
                       Ie501d0f392be1309df48c1616ace5a27: 
                       I29468f8318cd5bebb5cea27e1ee57b7f;
               I6043631f93e2c514d5ed6e86beffa7c6 =  Ie3f06a529d5f22198b3b33d649b740e1 ;
               Ibc084904fb63bb24102789357ce2cd76 =  I0456541b6e82ffeb05fc4052fafc41f7 ;
               I9e82413dca68de150b81bd27ab180980 =  Iabe05603679da24a44565e756adc0881 ;
               I4992c306a07d2e104a72dfcc37968e8c =  I98805e117c2f4ba4a8f6c2755ebe1fee ;
              I637c0445b26879a0fb9d7d94baef55e4 = 
          (!fgallag_sel[0]) ? 
                       Ia82b6e01034a63c2a1a446029f58f1c6: 
                       I05de7fd67a0e226201b563fa6c50f362;
               I3f1f9cecc45287a2c9487c04d8430b5b =  I8df8f128712fe5445a97566f8f29ecd4 ;
               Ife3d2f48786c2e11f7c4f8b4a7bb829e =  Ibcab213dbb173403005b3d65f780fa2d ;
              I0a019e2861b41f395bd12b43cd978e59 = 
          (!fgallag_sel[0]) ? 
                       Ide1a993a1dfca37107fc81e985714d93: 
                       I7004a1bc0ec2272163d33907d21616ea;
               I34fcd098fa2b426f98542121dae204fc =  I4ac93ed29241fee9390fd824452e6632 ;
               I8c9a0911720c403f2794fa5662a31207 =  I21281177f31dc70c65db2e9a3aa72392 ;
              I11af377ea2ae07f2249042a6daeef846 = 
          (!fgallag_sel[0]) ? 
                       I4cebb1a21b9c76387237fe8784f97ac1: 
                       I3b8cbc445627a75cc4b05aafc8a23cc5;
               Ib5d6d77cf92f29c1b498252859ec19ff =  I46c35e4856fb0288a23d9c4c68290ee9 ;
               I1d6100bd00e7e46af792dd99286391a5 =  I86454d943e7ff4b244882b0f6955d9df ;
               Ia6e85ec8c498ed70cb4a4e01bf8d1530 =  Id34d6ac40408151f201a8b3131463b3b ;
               Icc6d40c383e5580bbac65b6c77da6528 =  I3ffe132daa39f108095cd1fd5c38c6d6 ;
               Id939e83f81205a66485908e0bba8504d =  I080d693c8cdddee8f9c80ad68d1db1fe ;
               Ie709765eec241ae95c588fbfed18a87e =  I30ce714aeca130dc1978c6eda3ec0e11 ;
               I497fb247a6572f689aea3e595e657fdb =  Icd76d18cf8b38caaafc592047ff3b48c ;
               I659b78a601b47941441dc1debcae4d46 =  Ia29e3ba7f03b070d4381093dcafcdeb9 ;
               Ibed2d1ab1707ca759a8b09a5147a4268 =  I49dd3ecb280e2ea8639a2397343f1700 ;
               I23c058e418bad060fb1404b248782705 =  Iecf3c7051c364595cb29b47e8ceae9d7 ;
               I95f73f2e7a5268d25f4fcaa53339c2fc =  I1623b3a676440bab948f5f01c31c87a2 ;
               I90b927c01ca8d69239141958db410c54 =  I858523451a6554f7bc0238638450bb3d ;
               I79c64b98cdd4f4a1b41ddd2480c5d62a =  I88222b3d351f2f7334c9f3f22d3f0255 ;
               I76071439d501dfac67b1355c33f04c79 =  I2347ec4791ee62d976d13c7c6319e16a ;
               I3bed56f31105c1dd5524f2e04a6cdc0f =  I4c48730b147596406983412e0e6ae556 ;
               I1ca06bac6a4d082efeed13d0448630fb =  I70281a4f7bfe2fc5e4a0b91b4194d286 ;
               Iefd7ba660203932e953d509b10032e4d =  Ib9d8fdfe03633433eab48b80f9d4bae8 ;
               I76b3bd4ded426c469b208f83f7bb1781 =  I69f8f0b916f8d0b4d146e839c19a0756 ;
               I36261da4cc2946a22e80fb6f2a394753 =  Ic31af45750c67aca08c2af5f1fdc52d4 ;
               Iaa84b434bf0040f25a2dd6af77d90df4 =  Idec985d498536ef129885e9baaa69be5 ;
               I1a314b0ac2b2897b23d2e9fd3e5e63f0 =  I64c48585300f968447198fd11396fd71 ;
               I64eff7490d835e24cf4e5f4d0c60e18e =  I8d49cc394888a3e49b8e5cd72f2877e5 ;
               I95c886a9726c33f2a8f2f9413c9486cb =  I80802c2f239fbc3ed9bff61e9c873550 ;
              Ie2fbf1593b8aa394377ccc4ef0f705b6 = 
          (!fgallag_sel[0]) ? 
                       Ib8b1376de13c22be5126d585890438d7: 
                       I0a617772f4b574bc44555b85eb425b3a;
               I124a5e6d2c3103fbb4699cc2f7528a48 =  I3a9c038e7e278e6630b3defab662e10c ;
               I3625276282d727c6510f5123ee467e73 =  I878e4888b177aa7880c8ab11384db32a ;
               I771e25faed091d437e00dae0e66d088b =  If808ebd32478faac57b26b5306292dc4 ;
               Iad7a84f48832522261c3495844b19dde =  I88320212337ea2d63720b17e98675475 ;
               I8de675a8e37ed2b30a82e49ff6d510a0 =  I20f9fe0be090aee8bf1dcc46f806d73c ;
               I4bbc70e0a3a56eeb62af73e6c80006b4 =  I47c779e7352c5c5f13cccdd737dc994b ;
               I5c97bebf3cd2472e43ae7312d3956bb5 =  I7ae4796f21cd658ec17c8ff97f369784 ;
              I527847fbb55900e97761446b030ed540 = 
          (!fgallag_sel[0]) ? 
                       Idc1a3fedeccab7f0ee34f79366f5c4e5: 
                       Ie8117cdb093d8606a07c83ee8e80b388;
               Ie707c8b057532a88aff15ca43d1a4cef =  I0a65eb60e084d42aa5f5d9d6803068df ;
               I41708d131f34ee41b74f571661e751c6 =  Ia45d63e797413cb23c429c7d7a1eef02 ;
               I410af2866a81357ed84738c1800ee8e2 =  Ib89de4c510d53bd06fe0f10c7513de04 ;
               Iae78b53a85d3b3441bb251688c85fe66 =  I8b7353fd85fd2ee67a1df24a9f239f50 ;
               I1c4646eab74db4876187e2e87d861e4d =  I3ceb68a7f17d021fb3ce01821a19e7d8 ;
               Idb04b139376a9fd83c6f921b02c31849 =  Ia67f20bc0f3e32bf1e443bae34efc4b0 ;
               I64c0c3c0d18d18ed62b2b2910930f8a0 =  I6631364f87a3c0d43c4e1e433b61a132 ;
               I0c622446a77fe077062fd87448e11fec =  Ief1269d4009e33d56efce8d693d3588c ;
               Ie69cbbb6131f04ccf84db28990b4dbdd =  If36edf1833e16bf79b7ea16dcc551d2d ;
               Id0b467dbeaa2b30126ed60489530e29f =  I1cc0a80d74fe4b030cd838bd32b3cb20 ;
              Idac7b0bec594eccd74ac2d944da4484e = 
          (!fgallag_sel[0]) ? 
                       I4566be9ae01ab539195295433536bb4e: 
                       I9ba42ab3f14a648fa7ba73189a272474;
               I4ddb027f246fb2b145bba7b01687d39b =  I735b9bdb73b8701ec3181c5c08f9637c ;
               I754ff7341b379de55d5facc6fcc9f874 =  I78d31cfda6c9de83fbee1581d2cf4330 ;
               Ia7a71696b5ebed6c80cafb33a031626e =  Ie29fc0c82ccfe2e936226bbf8a22aa93 ;
               I542db58e949d7d1c542c075005fb065c =  I3b383604747befb7811e7cbda19108f2 ;
               I28aaa9370cb22a81b7c8d20fe7e1d347 =  I6e38e23fc4b5a6d9f5990d7f82f6a0c7 ;
               If4abfdcd468d4d98db5f32bb99303035 =  Id5737f058ffd0a11b2d29f088cf7591b ;
               Idfc14e592719d57828f8e6dc2130e270 =  Ib906993ed1101ad0992f24c4dae29370 ;
               Ia51b4598ba3f6c128ffcd421a3ba7309 =  I4c6811b2d28239598a23f790a03326fc ;
               Iee935e25f9fe5c7844bb0c0490cbb90f =  I9ac5de9728a0349bdb44341a68adeeec ;
               I05d0b3631f8501ecafcbb321c15be5f1 =  I969fc047ddc46bca31190e0d7f435bd9 ;
               I7ea9adf8dba141eef7a08d76105580ec =  I38083dfdf321de81daef5771d0546525 ;
               Ifa4cd939b137dc050f675a493546ddf6 =  I9d6d3cf2eccd6cba144db2459967a901 ;
               I7a6215a05dd8dbdcb421d7df535c5b67 =  I1cbd09f17301a0bee1cd695a2bde4e1c ;
               Ibd0c06d4190a37b90c51d562c6019551 =  I54b29fec4a88bc1e03197a0c55b875db ;
               I75b4b57cf9d7400feec38e037c948352 =  Ib4dee5c8efd8022bd9c3f9bf8d5e328b ;
              I14a4e51be5aa98fa28cc4740e6446747 = 
          (!fgallag_sel[0]) ? 
                       I3ae123c41c91d9b53a70aa3e4793be9b: 
                       If4ccd39857a7317488e9215271db7210;
               I43196769a96d15dd03318e43b48a6b4d =  Ief6d7060558cf2ccd8d561ec17b846d5 ;
               I8494b9c75594140fabc1158bacf4438a =  Ie03342fcc484bd9f1c934e675c9f6ec4 ;
               I931bf44a358d9fd91d31aa78d3e16312 =  Idb2832cb2e894a8c02e7dab1dccdef87 ;
               I5355f3939098f1ae0aa0f254b8e7e163 =  I8f9db21a5dea66f9865796d164f689ea ;
               I6228ab1c737aec5845684c0eff41dac4 =  I2135e15ed882d1293741fd593369f88d ;
               I9034255c2128aa8c4d707bf003a57e86 =  I5e298171856ae5526301f6d5084f2796 ;
               Ia9bc32f3ef4f4681782fec452e572cf2 =  I1b7e4002a74d5f33e7d0168ed06aaa2d ;
               I9791a65b490a63c3c201409a30b86199 =  Ibe26ea03448b95798236cf228817dfd0 ;
               Id5297cb2f91d5b3e67c4bd97a8c05401 =  I21d9dac9d09da39f435c7082dca90127 ;
               Ibc826b606b10904061b2666eb204469e =  I8546eab32336885c49882f192be9904c ;
               I06dabbc9dc6fb6b8fa517e188ee74208 =  I8c50bd38d4339a6ae19e13db1a1994e9 ;
               I4d3607d7cd13b86ae4a22bebaf65ef0e =  Ia98d1ff0d0dac6a253cf48ab85e0eb75 ;
               Ia974eebd7b7563b2f0822f538c13a911 =  I0b963cc516bb0de18221dd724864d795 ;
               I191470ccfa2c2838a34aceb571582bb4 =  I7f856b89e8b206458e96335076d80c69 ;
               I01714219c84cfbfd7ff940108ddbb6b3 =  I72569b57d65e91bcea79d0682c51c4a7 ;
               I118d11a015af5944d64290a46bf49c09 =  Iad3645f6fa7141133b12534c70efc80c ;
               Ib878ef5592b0bf1af247ede54fe13a45 =  Id7216252c1febf54691e626861f6215c ;
               I7686f623f51c5a9f8f3f8d143ed8bcb5 =  Id25c2945168c44ec9f0a4bb2dc6aaf68 ;
               I4d48fc8081756af036b8f1b1b9e56051 =  I2b3c4fca6b0feb6fd829e9cbbe9d7142 ;
               Ia1d93d4bbc6b1e73dbb0c6c26d102f10 =  I7858226bb4feb944c5feaa52f2b51034 ;
               Ifb7d0d12a916fc3f2f9c0341f27ef53f =  I1201c86e1f6f9e890181790896c4afa4 ;
               I4ee596c96f91a18ef1ebb0ee6de285ae =  I3920223ae6d1a6d2ff327f53933ecad4 ;
               I5aeda0b5dc8459d86e9ab5082bf9fed8 =  Id23811d7cf32f6c5c63ce2782da15720 ;
               I7b6ff145fa076d152af672e0c3a062bc =  I7a01b2b85d70a35d44836e181a22b322 ;
               I3929cfb9fb8795d4dd9f54f9c4a2fa02 =  I45b1d972b2a5028cc340988f7c37f2e0 ;
               If33f043047ad17b323733a201aa649da =  I389856ba7ca6568e4ead3483c3e52353 ;
               Icfb9314b47604c3b065ffdd5d9042682 =  I591624fd56ff315e0084af5af206cf8e ;
               I5cd61f07b490ca79f1ec069ed2d47528 =  I92793401ab28d5ed265775c0d165dfe5 ;
               I1bace448ce54ae41e9e8d27acf548338 =  I3c28bfe18fb1543683ae264c396a0207 ;
               I692bf3f934f0ee8fbf02c7dce98f924c =  I2fd3c0dfd43b65e2fe8afd3368a50fc5 ;
               Ifb3af535b42775dae1e0ade2d8bf79df =  I22bbdf426df953feb5acede78c31b9b2 ;
               I569a621522dd636df609f60c1b22d7f7 =  I687ab1878d38c7c988507163c8a60070 ;
               Ic651187a36eb89eaf129a368af3474ee =  Id7f7499e9b3f529781f4aba6e63490ac ;
               Ib120bd9cfec97e7956bb64f8e4527caf =  I730aeccac38e1622c684c468f8cb29f4 ;
               I41e452eee26c8ede812d3ca957488aec =  Iba910435a91ee873f76fa3ec9ac9c3d3 ;
