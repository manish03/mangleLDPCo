//`include "GF2_LDPC_fgallag_0x0000b_assign_inc.sv"
//always_comb begin
              Ibbc4b022828a232d4b3d3eccc478fd3f['h00000] = 
          (!fgallag_sel['h0000b]) ? 
                       I45c1a80dd59b47025bbf3f233589964b['h00000] : //%
                       I45c1a80dd59b47025bbf3f233589964b['h00001] ;
//end
//always_comb begin
              Ibbc4b022828a232d4b3d3eccc478fd3f['h00001] = 
          (!fgallag_sel['h0000b]) ? 
                       I45c1a80dd59b47025bbf3f233589964b['h00002] : //%
                       I45c1a80dd59b47025bbf3f233589964b['h00003] ;
//end
//always_comb begin
              Ibbc4b022828a232d4b3d3eccc478fd3f['h00002] = 
          (!fgallag_sel['h0000b]) ? 
                       I45c1a80dd59b47025bbf3f233589964b['h00004] : //%
                       I45c1a80dd59b47025bbf3f233589964b['h00005] ;
//end
//always_comb begin
              Ibbc4b022828a232d4b3d3eccc478fd3f['h00003] = 
          (!fgallag_sel['h0000b]) ? 
                       I45c1a80dd59b47025bbf3f233589964b['h00006] : //%
                       I45c1a80dd59b47025bbf3f233589964b['h00007] ;
//end
//always_comb begin
              Ibbc4b022828a232d4b3d3eccc478fd3f['h00004] = 
          (!fgallag_sel['h0000b]) ? 
                       I45c1a80dd59b47025bbf3f233589964b['h00008] : //%
                       I45c1a80dd59b47025bbf3f233589964b['h00009] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00005] =  I45c1a80dd59b47025bbf3f233589964b['h0000a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00006] =  I45c1a80dd59b47025bbf3f233589964b['h0000c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00007] =  I45c1a80dd59b47025bbf3f233589964b['h0000e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00008] =  I45c1a80dd59b47025bbf3f233589964b['h00010] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00009] =  I45c1a80dd59b47025bbf3f233589964b['h00012] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0000a] =  I45c1a80dd59b47025bbf3f233589964b['h00014] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0000b] =  I45c1a80dd59b47025bbf3f233589964b['h00016] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0000c] =  I45c1a80dd59b47025bbf3f233589964b['h00018] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0000d] =  I45c1a80dd59b47025bbf3f233589964b['h0001a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0000e] =  I45c1a80dd59b47025bbf3f233589964b['h0001c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0000f] =  I45c1a80dd59b47025bbf3f233589964b['h0001e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00010] =  I45c1a80dd59b47025bbf3f233589964b['h00020] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00011] =  I45c1a80dd59b47025bbf3f233589964b['h00022] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00012] =  I45c1a80dd59b47025bbf3f233589964b['h00024] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00013] =  I45c1a80dd59b47025bbf3f233589964b['h00026] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00014] =  I45c1a80dd59b47025bbf3f233589964b['h00028] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00015] =  I45c1a80dd59b47025bbf3f233589964b['h0002a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00016] =  I45c1a80dd59b47025bbf3f233589964b['h0002c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00017] =  I45c1a80dd59b47025bbf3f233589964b['h0002e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00018] =  I45c1a80dd59b47025bbf3f233589964b['h00030] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00019] =  I45c1a80dd59b47025bbf3f233589964b['h00032] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0001a] =  I45c1a80dd59b47025bbf3f233589964b['h00034] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0001b] =  I45c1a80dd59b47025bbf3f233589964b['h00036] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0001c] =  I45c1a80dd59b47025bbf3f233589964b['h00038] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0001d] =  I45c1a80dd59b47025bbf3f233589964b['h0003a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0001e] =  I45c1a80dd59b47025bbf3f233589964b['h0003c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0001f] =  I45c1a80dd59b47025bbf3f233589964b['h0003e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00020] =  I45c1a80dd59b47025bbf3f233589964b['h00040] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00021] =  I45c1a80dd59b47025bbf3f233589964b['h00042] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00022] =  I45c1a80dd59b47025bbf3f233589964b['h00044] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00023] =  I45c1a80dd59b47025bbf3f233589964b['h00046] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00024] =  I45c1a80dd59b47025bbf3f233589964b['h00048] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00025] =  I45c1a80dd59b47025bbf3f233589964b['h0004a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00026] =  I45c1a80dd59b47025bbf3f233589964b['h0004c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00027] =  I45c1a80dd59b47025bbf3f233589964b['h0004e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00028] =  I45c1a80dd59b47025bbf3f233589964b['h00050] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00029] =  I45c1a80dd59b47025bbf3f233589964b['h00052] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0002a] =  I45c1a80dd59b47025bbf3f233589964b['h00054] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0002b] =  I45c1a80dd59b47025bbf3f233589964b['h00056] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0002c] =  I45c1a80dd59b47025bbf3f233589964b['h00058] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0002d] =  I45c1a80dd59b47025bbf3f233589964b['h0005a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0002e] =  I45c1a80dd59b47025bbf3f233589964b['h0005c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0002f] =  I45c1a80dd59b47025bbf3f233589964b['h0005e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00030] =  I45c1a80dd59b47025bbf3f233589964b['h00060] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00031] =  I45c1a80dd59b47025bbf3f233589964b['h00062] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00032] =  I45c1a80dd59b47025bbf3f233589964b['h00064] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00033] =  I45c1a80dd59b47025bbf3f233589964b['h00066] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00034] =  I45c1a80dd59b47025bbf3f233589964b['h00068] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00035] =  I45c1a80dd59b47025bbf3f233589964b['h0006a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00036] =  I45c1a80dd59b47025bbf3f233589964b['h0006c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00037] =  I45c1a80dd59b47025bbf3f233589964b['h0006e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00038] =  I45c1a80dd59b47025bbf3f233589964b['h00070] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00039] =  I45c1a80dd59b47025bbf3f233589964b['h00072] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0003a] =  I45c1a80dd59b47025bbf3f233589964b['h00074] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0003b] =  I45c1a80dd59b47025bbf3f233589964b['h00076] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0003c] =  I45c1a80dd59b47025bbf3f233589964b['h00078] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0003d] =  I45c1a80dd59b47025bbf3f233589964b['h0007a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0003e] =  I45c1a80dd59b47025bbf3f233589964b['h0007c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0003f] =  I45c1a80dd59b47025bbf3f233589964b['h0007e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00040] =  I45c1a80dd59b47025bbf3f233589964b['h00080] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00041] =  I45c1a80dd59b47025bbf3f233589964b['h00082] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00042] =  I45c1a80dd59b47025bbf3f233589964b['h00084] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00043] =  I45c1a80dd59b47025bbf3f233589964b['h00086] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00044] =  I45c1a80dd59b47025bbf3f233589964b['h00088] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00045] =  I45c1a80dd59b47025bbf3f233589964b['h0008a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00046] =  I45c1a80dd59b47025bbf3f233589964b['h0008c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00047] =  I45c1a80dd59b47025bbf3f233589964b['h0008e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00048] =  I45c1a80dd59b47025bbf3f233589964b['h00090] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00049] =  I45c1a80dd59b47025bbf3f233589964b['h00092] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0004a] =  I45c1a80dd59b47025bbf3f233589964b['h00094] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0004b] =  I45c1a80dd59b47025bbf3f233589964b['h00096] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0004c] =  I45c1a80dd59b47025bbf3f233589964b['h00098] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0004d] =  I45c1a80dd59b47025bbf3f233589964b['h0009a] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0004e] =  I45c1a80dd59b47025bbf3f233589964b['h0009c] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0004f] =  I45c1a80dd59b47025bbf3f233589964b['h0009e] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00050] =  I45c1a80dd59b47025bbf3f233589964b['h000a0] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00051] =  I45c1a80dd59b47025bbf3f233589964b['h000a2] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00052] =  I45c1a80dd59b47025bbf3f233589964b['h000a4] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00053] =  I45c1a80dd59b47025bbf3f233589964b['h000a6] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00054] =  I45c1a80dd59b47025bbf3f233589964b['h000a8] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00055] =  I45c1a80dd59b47025bbf3f233589964b['h000aa] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00056] =  I45c1a80dd59b47025bbf3f233589964b['h000ac] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00057] =  I45c1a80dd59b47025bbf3f233589964b['h000ae] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00058] =  I45c1a80dd59b47025bbf3f233589964b['h000b0] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00059] =  I45c1a80dd59b47025bbf3f233589964b['h000b2] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0005a] =  I45c1a80dd59b47025bbf3f233589964b['h000b4] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0005b] =  I45c1a80dd59b47025bbf3f233589964b['h000b6] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0005c] =  I45c1a80dd59b47025bbf3f233589964b['h000b8] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0005d] =  I45c1a80dd59b47025bbf3f233589964b['h000ba] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0005e] =  I45c1a80dd59b47025bbf3f233589964b['h000bc] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0005f] =  I45c1a80dd59b47025bbf3f233589964b['h000be] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00060] =  I45c1a80dd59b47025bbf3f233589964b['h000c0] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00061] =  I45c1a80dd59b47025bbf3f233589964b['h000c2] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00062] =  I45c1a80dd59b47025bbf3f233589964b['h000c4] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00063] =  I45c1a80dd59b47025bbf3f233589964b['h000c6] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00064] =  I45c1a80dd59b47025bbf3f233589964b['h000c8] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00065] =  I45c1a80dd59b47025bbf3f233589964b['h000ca] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00066] =  I45c1a80dd59b47025bbf3f233589964b['h000cc] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00067] =  I45c1a80dd59b47025bbf3f233589964b['h000ce] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00068] =  I45c1a80dd59b47025bbf3f233589964b['h000d0] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00069] =  I45c1a80dd59b47025bbf3f233589964b['h000d2] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0006a] =  I45c1a80dd59b47025bbf3f233589964b['h000d4] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0006b] =  I45c1a80dd59b47025bbf3f233589964b['h000d6] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0006c] =  I45c1a80dd59b47025bbf3f233589964b['h000d8] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0006d] =  I45c1a80dd59b47025bbf3f233589964b['h000da] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0006e] =  I45c1a80dd59b47025bbf3f233589964b['h000dc] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0006f] =  I45c1a80dd59b47025bbf3f233589964b['h000de] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00070] =  I45c1a80dd59b47025bbf3f233589964b['h000e0] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00071] =  I45c1a80dd59b47025bbf3f233589964b['h000e2] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00072] =  I45c1a80dd59b47025bbf3f233589964b['h000e4] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00073] =  I45c1a80dd59b47025bbf3f233589964b['h000e6] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00074] =  I45c1a80dd59b47025bbf3f233589964b['h000e8] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00075] =  I45c1a80dd59b47025bbf3f233589964b['h000ea] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00076] =  I45c1a80dd59b47025bbf3f233589964b['h000ec] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00077] =  I45c1a80dd59b47025bbf3f233589964b['h000ee] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00078] =  I45c1a80dd59b47025bbf3f233589964b['h000f0] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h00079] =  I45c1a80dd59b47025bbf3f233589964b['h000f2] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0007a] =  I45c1a80dd59b47025bbf3f233589964b['h000f4] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0007b] =  I45c1a80dd59b47025bbf3f233589964b['h000f6] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0007c] =  I45c1a80dd59b47025bbf3f233589964b['h000f8] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0007d] =  I45c1a80dd59b47025bbf3f233589964b['h000fa] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0007e] =  I45c1a80dd59b47025bbf3f233589964b['h000fc] ;
//end
//always_comb begin // 
               Ibbc4b022828a232d4b3d3eccc478fd3f['h0007f] =  I45c1a80dd59b47025bbf3f233589964b['h000fe] ;
//end
