 reg  ['h7f:0] [$clog2('h7000+1)-1:0] I9b3a227f14d8af7af837f644f90f9897fc24e24ae598906ef48809ee1fccd211 ;
