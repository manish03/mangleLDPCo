 reg  ['h3ff:0] [$clog2('h7000+1)-1:0] Icff8af1f5c3ae89ef95ed8451273154b ;
