//`include "GF2_LDPC_fgallag_0x0000b_assign_inc.sv"
//always_comb begin
              Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00000] = 
          (!fgallag_sel['h0000b]) ? 
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00000] : //%
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00001] ;
//end
//always_comb begin
              Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00001] = 
          (!fgallag_sel['h0000b]) ? 
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00002] : //%
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00003] ;
//end
//always_comb begin
              Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00002] = 
          (!fgallag_sel['h0000b]) ? 
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00004] : //%
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00005] ;
//end
//always_comb begin
              Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00003] = 
          (!fgallag_sel['h0000b]) ? 
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00006] : //%
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00007] ;
//end
//always_comb begin
              Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00004] = 
          (!fgallag_sel['h0000b]) ? 
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00008] : //%
                       Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00009] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00005] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00006] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00007] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0000e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00008] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00010] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00009] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00012] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0000a] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00014] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0000b] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00016] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0000c] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00018] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0000d] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0000e] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0000f] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0001e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00010] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00020] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00011] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00022] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00012] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00024] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00013] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00026] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00014] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00028] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00015] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00016] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00017] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0002e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00018] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00030] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00019] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00032] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0001a] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00034] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0001b] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00036] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0001c] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00038] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0001d] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0001e] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0001f] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0003e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00020] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00040] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00021] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00042] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00022] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00044] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00023] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00046] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00024] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00048] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00025] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00026] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00027] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0004e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00028] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00050] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00029] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00052] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0002a] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00054] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0002b] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00056] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0002c] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00058] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0002d] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0002e] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0002f] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0005e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00030] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00060] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00031] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00062] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00032] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00064] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00033] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00066] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00034] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00068] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00035] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00036] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00037] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0006e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00038] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00070] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00039] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00072] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0003a] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00074] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0003b] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00076] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0003c] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00078] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0003d] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0003e] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0003f] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0007e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00040] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00080] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00041] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00082] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00042] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00084] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00043] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00086] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00044] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00088] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00045] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00046] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00047] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0008e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00048] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00090] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00049] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00092] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0004a] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00094] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0004b] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00096] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0004c] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h00098] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0004d] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009a] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0004e] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009c] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0004f] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h0009e] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00050] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a0] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00051] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a2] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00052] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a4] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00053] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a6] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00054] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000a8] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00055] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000aa] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00056] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ac] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00057] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ae] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00058] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b0] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00059] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b2] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0005a] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b4] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0005b] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b6] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0005c] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000b8] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0005d] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ba] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0005e] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000bc] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0005f] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000be] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00060] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c0] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00061] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c2] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00062] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c4] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00063] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c6] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00064] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000c8] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00065] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ca] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00066] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000cc] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00067] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ce] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00068] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d0] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00069] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d2] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0006a] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d4] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0006b] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d6] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0006c] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000d8] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0006d] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000da] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0006e] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000dc] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0006f] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000de] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00070] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e0] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00071] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e2] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00072] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e4] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00073] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e6] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00074] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000e8] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00075] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ea] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00076] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ec] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00077] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000ee] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00078] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f0] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h00079] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f2] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0007a] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f4] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0007b] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f6] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0007c] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000f8] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0007d] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000fa] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0007e] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000fc] ;
//end
//always_comb begin // 
               Iab9b2227df9be85847d2443b8646d4fc421de8fd5d60f08364bd1704f7631d96['h0007f] =  Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765['h000fe] ;
//end
