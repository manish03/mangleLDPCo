//`include "GF2_LDPC_fgallag_0x0000f_assign_inc.sv"
//always_comb begin
              I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00000] = 
          (!fgallag_sel['h0000f]) ? 
                       I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00000] : //%
                       I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00001] ;
//end
//always_comb begin // 
               I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00001] =  I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00002] ;
//end
//always_comb begin // 
               I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00002] =  I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00004] ;
//end
//always_comb begin // 
               I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00003] =  I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00006] ;
//end
//always_comb begin // 
               I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00004] =  I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h00008] ;
//end
//always_comb begin // 
               I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00005] =  I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000a] ;
//end
//always_comb begin // 
               I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00006] =  I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000c] ;
//end
//always_comb begin // 
               I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00007] =  I333510d8572134ddfb62c52fc8869a236241ec893f038dd668e3222609245de0['h0000e] ;
//end
