//`include "GF2_LDPC_flogtanh_0x0000e_assign_inc.sv"
//always_comb begin
              Iaf491f5f8d1574e1cb610cbd3edeca68['h00000] = 
          (!flogtanh_sel['h0000e]) ? 
                       If72de6675c42172560d5d150642f3da8['h00000] : //%
                       If72de6675c42172560d5d150642f3da8['h00001] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00001] =  If72de6675c42172560d5d150642f3da8['h00002] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00002] =  If72de6675c42172560d5d150642f3da8['h00004] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00003] =  If72de6675c42172560d5d150642f3da8['h00006] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00004] =  If72de6675c42172560d5d150642f3da8['h00008] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00005] =  If72de6675c42172560d5d150642f3da8['h0000a] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00006] =  If72de6675c42172560d5d150642f3da8['h0000c] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00007] =  If72de6675c42172560d5d150642f3da8['h0000e] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00008] =  If72de6675c42172560d5d150642f3da8['h00010] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h00009] =  If72de6675c42172560d5d150642f3da8['h00012] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h0000a] =  If72de6675c42172560d5d150642f3da8['h00014] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h0000b] =  If72de6675c42172560d5d150642f3da8['h00016] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h0000c] =  If72de6675c42172560d5d150642f3da8['h00018] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h0000d] =  If72de6675c42172560d5d150642f3da8['h0001a] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h0000e] =  If72de6675c42172560d5d150642f3da8['h0001c] ;
//end
//always_comb begin // 
               Iaf491f5f8d1574e1cb610cbd3edeca68['h0000f] =  If72de6675c42172560d5d150642f3da8['h0001e] ;
//end
