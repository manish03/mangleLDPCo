 reg  ['h3:0] [$clog2('h7000+1)-1:0] I3bcb7ea9f76eac891526e809fd382eaceb4a8f0a204c5ca7f391e7ffd9b7808f ;
