 reg  ['hff:0] [$clog2('h7000+1)-1:0] Ib63bfb495d94b2b5cc4c9a90f4ac9fec84b80dd3e7527c86056af3ff3922a765 ;
