reg [fgallag_WDTH -1:0] I84ab01f2ac31304c9525b8983d34300d, I72dd1fc26b57d741390612b9bcffab1d;
reg [fgallag_WDTH -1:0] Iaf7ae8cb478fce9deaf537c13fa083cb, I98c43e93e5f943a7b07ef09985f97014;
reg [fgallag_WDTH -1:0] Idce9e18b46f498af68bbb108da7441bc, I434c16361fa147e26f4d2c4cc6d69150;
reg [fgallag_WDTH -1:0] Ie3954c25e29ea2d7e1340a59d3d7165f, I9e87743bade1ee6fbfdd119cbdb0a3cb;
reg [fgallag_WDTH -1:0] Iaa12f10c6588df5d8d8444c61b422c7c, I1e6255cf954cd5a58c52ff8e6a55bdbc;
reg [fgallag_WDTH -1:0] I9851178cd4e84140f2c244f19c285e4a, I77a73f3832687dababc30666ac62d1af;
reg [fgallag_WDTH -1:0] I463cc1b85874882aadc9fa0ed9eb7816, Iacdfa68e9ab161a0e6c7e559b9954640;
reg [fgallag_WDTH -1:0] I5249c4136a601a94d06d4955be304799, Iedc0dfa42eaada48be02e65be4b39615;
reg [fgallag_WDTH -1:0] I9ce88b0e18af39ed6dc46db59a2bb78b, Ib4fb78755c536a284004e41f584d99fb;
reg [fgallag_WDTH -1:0] I3695c8773a6d76c02a9f8849ada96902, I5156cd5e3f0fe53ad559b342c818f41a;
reg [fgallag_WDTH -1:0] I4783f15f954421f7538cf39210bb44d5, I3cf816bf7fd922df289b13766e931e17;
reg [fgallag_WDTH -1:0] Ia82244e3d80e219740368bab411242be, Ibf2a30f91bd9050391913c02be7c8cad;
reg [fgallag_WDTH -1:0] Ib42df9a31ffd2cfc4a63cf95cf89c4d7, Iea12e263d5883f93023d784884645969;
reg [fgallag_WDTH -1:0] I752d56e6caa726064dc20d4eeda763a9, I550762460d0217d3c91c5112546b7929;
reg [fgallag_WDTH -1:0] Ie339fd09fbad7893452b9a2f92d45932, I0d8eaf22a03a0102d8bf7a53a7737943;
reg [fgallag_WDTH -1:0] Ifd15d58d88de80f2cfc98c7f66f8f88d, I8017a4f092179605074076e8b5690842;
reg [fgallag_WDTH -1:0] I994cd956aabc31d730d77d9b67bbc1db, I57160990c295512e2d98c301632c5120;
reg [fgallag_WDTH -1:0] Ie7086ba45d27b8fd48ad4dbbc1a6466b, Id9f3f35bc6917416d6826d471f8ea441;
reg [fgallag_WDTH -1:0] I8539ebc561f7f4d823623b1f11255213, I6c9a443b704a7871ac13f164c1cdc88b;
reg [fgallag_WDTH -1:0] Iedbd35fd7ebaf3787a08b0551ffb324e, I76498f1e58ff35dc6153f76999f9f7a5;
reg [fgallag_WDTH -1:0] I23df575a91b34e0a642bf679a74a747c, I200025a860f318f6ff9aaf89b146d16f;
reg [fgallag_WDTH -1:0] Icce0e60e3e31993ef47683a80567b1c4, I107ae84d631e3a9574b62f4fdfe56140;
reg [fgallag_WDTH -1:0] I172b401633d8844fcabdd4b980f46c73, Ief394bcabeb27c95f3dabe3d5c0bd643;
reg [fgallag_WDTH -1:0] I71ed80b7d77c2a35edcefe9ce7db28af, Ibc52ae3742f657ac6abefd988494c8a1;
reg [fgallag_WDTH -1:0] Ib1873b0070c00bfe5ed6fda941cfe95e, I969ac5f2b8a9d6778300e3a91968ae4b;
reg [fgallag_WDTH -1:0] I6db83f8bbff7cde9c9db248c02fd9358, I3172be9cafebc7121994917ff35b25fb;
reg [fgallag_WDTH -1:0] If65d96ffe364426e1b90303ad323e7fb, I388e0d1c3f421d7522d6c0521538693e;
reg [fgallag_WDTH -1:0] I8e6c7979ddefa5e27581107ca2495e3e, I0fa0bdc864c6173b380c763cf3e794ba;
reg [fgallag_WDTH -1:0] I161c2f4e7657ff863ec2a319ee8d21d5, I9d6dc129ad747412224b487c4973db3a;
reg [fgallag_WDTH -1:0] Ic18bc04d9a02bccce383f311102a8b45, Ic1c5ee07ecd5c9fc9c2c1f9c33cdca08;
reg [fgallag_WDTH -1:0] I8a118ced20140ec0f90f1f82161bd2c1, I1b2ba3544e2d26b40edbfaedf137812b;
reg [fgallag_WDTH -1:0] I2b73e4b6134a9ca11b301452734741a1, Ieb654d27e0306c60cd9eff05f4be76ca;
reg [fgallag_WDTH -1:0] Ie432836bf5a95e8dbb6de2c29d9ab058, I462601141783fc299a3b081023233a56;
reg [fgallag_WDTH -1:0] I8a777efecfec25782e29fd4e8f270490, I4e4e1489c822058cf54782c75c8d6996;
reg [fgallag_WDTH -1:0] I3ad4e40b398385b2c3a94cabd4736926, I361a262df08182fcb917b7aa7aa73465;
reg [fgallag_WDTH -1:0] Ifcd756c806de58265e16199e27f64e22, Ic8092176d020f45ae84ae72da9ea20a8;
reg [fgallag_WDTH -1:0] Icac3b989b3d04d9c7a80d5eebcbb2027, I361a7201d61113929f346f8b22ac01ef;
reg [fgallag_WDTH -1:0] I806f4137adef04fa14f4c159fd47bb46, I616e26bab7d9ada350f152cce0ac3569;
reg [fgallag_WDTH -1:0] I6f6db1dfb50f19379683f16c549624b3, I7cb33be246a06045ff19436b47ccfdca;
reg [fgallag_WDTH -1:0] Ib26efe2924ee3c384a8f8b0f7f63e0f4, Ic5aad088ddcc97dd7a3c8244a27a288e;
reg [fgallag_WDTH -1:0] I0a45d8f9e12c5234855b972d39246589, I79c0e02b51ed3b20ca6de475189b6a48;
reg [fgallag_WDTH -1:0] I7a9fe30fbe486c1fd6d92b334f04a97b, I059966174241b59374640dc43018c49c;
reg [fgallag_WDTH -1:0] Ia5bc1b93ee0908ca26a967bc4720e5c3, I1b43d5eb392150245e2a303582b9226f;
reg [fgallag_WDTH -1:0] I6cd39d0d0d14283cd00870fa8697cbe2, Icc5e7d899df8ec350f804c1f32b9fe72;
reg [fgallag_WDTH -1:0] Id33e3cde2a62f32d114a78300c2fdc1b, I2f8fbab2b60878195ae8b2e1c0ff1208;
reg [fgallag_WDTH -1:0] I22f6c61d2512a383ecc57e2dac6e346a, I30e9a6bb0816599ede1e93a3091a572c;
reg [fgallag_WDTH -1:0] I00b3081cd7dd077a53bdd7781b98fe6c, I815a192d304aedca5f772d6bd401ad3f;
reg [fgallag_WDTH -1:0] Ibdf94fc4ee66c4af146968bf34ae4c0c, Id7c921ad25499d1e0bcf7dc1359e6b5d;
reg [fgallag_WDTH -1:0] Idadb48591ec328a331bdcf45e9156485, I83ce7e2b4c276008c33a5703eba16572;
reg [fgallag_WDTH -1:0] I6315c142854dc3c1893bcb08b46bc739, I96daacb3d66626af1c7b54c8be02a79b;
reg [fgallag_WDTH -1:0] I362b966433fe2df6176a09951d0d88db, I984e48eb72dcef91797c57289ba1322e;
reg [fgallag_WDTH -1:0] If210d0b145e2fd9cb2e1229c2c9c7a36, I8a0f063aab90c7f50f8eff7e3626483d;
reg [fgallag_WDTH -1:0] Ia133b750fb093f377556735adb4e3097, Ia49e2201160f9da0d475b16d22efcac1;
reg [fgallag_WDTH -1:0] I6d2fcf19c79a538ec57aff56b8579def, I59718bd7f0e7a0c9d63a038f2cb9d3eb;
reg [fgallag_WDTH -1:0] If507c9ebcb1bc24a59ab4a00fc902d88, I7e703dc56c5c5604eb8e7ed32fd6ce78;
reg [fgallag_WDTH -1:0] I70be43895e7446395ee6f209431a4b0e, I1475899d2bf7a51aeae5168d5af0d548;
reg [fgallag_WDTH -1:0] Iec863324907434f27365ce30e0a3a636, If3582b232dccd45a4f3c07514062003c;
reg [fgallag_WDTH -1:0] Ifdd6e035d37dc6a726502ea875e19bf2, I79a9448f1efc66a407e2dcc243638e6f;
reg [fgallag_WDTH -1:0] I0bac49aa5c179287d028c0bbe2f26646, I57fb6daf7238618d7ce10989a7f41025;
reg [fgallag_WDTH -1:0] I676f1d8111d39181de6fb867fcc8aad9, Ia677f2eaa008b296dc5eefdf680a2783;
reg [fgallag_WDTH -1:0] Ib6003647304cdf7e04f112ea1434d0c2, I629cd82c8226c17eb439cd2ad664a3b7;
reg [fgallag_WDTH -1:0] I32f1ca64465d5ffd4c0abef6a0713795, I181b85fc5fda9b5b99763bd8fa4a20b7;
reg [fgallag_WDTH -1:0] Iab2dbd174b3566d2eb0c32118a1d6ffc, Ida422d40a8abb52f4c78b63807f0ef16;
reg [fgallag_WDTH -1:0] I119a639a5c5243e5bbf6224fea9e0542, Ic91b7435580f54bb1e3ffa6ea1b21f69;
reg [fgallag_WDTH -1:0] I51a744f6026f58a3ff9d47f7ad8441c7, Id1651e9d3e909ddb1f3779b4129713fd;
reg [fgallag_WDTH -1:0] Ied88a6d77466adfacecc91792e092022, I470b1c602adb0b16c6b3a19133a97641;
reg [fgallag_WDTH -1:0] I531565b08841415ba9f98966030529f2, I81c0a5fad7512ba9d8537018d6df2c23;
reg [fgallag_WDTH -1:0] I35641e3719c76fbc8621771af415d10f, I0ea14616a599bd3f1c59dd57652ce967;
reg [fgallag_WDTH -1:0] I56baf72a394546e751edf096f5a87970, Ia6503d131655b73ae90b5553d116e92b;
reg [fgallag_WDTH -1:0] I07ab92c9ad141c03101d587f00202c81, I2548ee3c3bf2a2eaa2ed541546e58c04;
reg [fgallag_WDTH -1:0] I0143dfa3c201c85bdcce5739dee11814, I2c197653e4a8776ad3539f95aff27df5;
reg [fgallag_WDTH -1:0] Ie9a0ea695884198a9fd7e5de0a9f73d0, I0d6cfa3166445e1396871afad62fba40;
reg [fgallag_WDTH -1:0] I0a066ff1810c068d1807dd5999880170, Ie597ab8c4dd174055b4bda8dbdec0dd3;
reg [fgallag_WDTH -1:0] I3d390c1d2a5df6decbc45bd682760b84, I46ee4c21a9801d95f803c4408dba7ea0;
reg [fgallag_WDTH -1:0] I0b1c32f0732334693986eea6aaee2b12, I9426c6803cf8c7c6dbc422989eef5380;
reg [fgallag_WDTH -1:0] Ifb9c5b70184594cb9f7961cb99c0d62e, I299fbb7b05d282681f0e9704b7818b0d;
reg [fgallag_WDTH -1:0] I105a0656b51423653fd7428001efa81f, I947d66b22e42c68930e8bf7d1439a376;
reg [fgallag_WDTH -1:0] Id9515c02ee595dc6ce4353decfbd2928, I4e1752e19a8ec547211ca30f0e85c2d5;
reg [fgallag_WDTH -1:0] Ib1d40c92e79f6562475204ba330c15e3, I22715ee56f34e2c7cfdae2dd409ac653;
reg [fgallag_WDTH -1:0] Ief1a527fee16c6cb996ca3363d4713d8, I85be91ab3b8a799d6681b90e6f56ad5e;
reg [fgallag_WDTH -1:0] I5c7ed7d4a522cf1e94035b3475d07240, Id2e3d5dfe5c8ec9128f5a719175c0f35;
reg [fgallag_WDTH -1:0] Ie59496301d7ef6565b69072f4530ceee, I16d052ce0d66bc9f49489a124ccf6c69;
reg [fgallag_WDTH -1:0] I2d2b69150858f521850b9d71ee17acbf, I0f1ace68f720dfcca74605ec277d0067;
reg [fgallag_WDTH -1:0] I0556476f50843423945a3783fd5c9612, I02f31af05294d3f39fe7c2f3a71a300a;
reg [fgallag_WDTH -1:0] I34f9b6d4f00ab598a94274629c08e99c, Ia10e05a72a5d3c1e16b99510e94f6121;
reg [fgallag_WDTH -1:0] I2f16d9a27f31109e57160fbc03a98853, I8b94c6d56df2d4a9a2adc2c7ccb8a0a9;
reg [fgallag_WDTH -1:0] Ib19a79508dff3510b087cb2c1df176f9, I8b6f4ea7a19f4b359aa01867c4502ccf;
reg [fgallag_WDTH -1:0] I48ac3afb4f8b31f9aadc59aaf1a28a44, Id2add03142e6a3e5f4625082fbcc46ed;
reg [fgallag_WDTH -1:0] Ia3bbc4519f9cd9651e10efaace317875, I323124e6fcbab5bdda4bd24c7b2a99c1;
reg [fgallag_WDTH -1:0] I51118baae7de42e5f69f1a78d1ceccad, Ib943a483749ffc791a5965ed0840bb0f;
reg If379a89ad17fd061bf987e29aa713945 ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I72dd1fc26b57d741390612b9bcffab1d <= 'h0;
 I98c43e93e5f943a7b07ef09985f97014 <= 'h0;
 I434c16361fa147e26f4d2c4cc6d69150 <= 'h0;
 I9e87743bade1ee6fbfdd119cbdb0a3cb <= 'h0;
 I1e6255cf954cd5a58c52ff8e6a55bdbc <= 'h0;
 I77a73f3832687dababc30666ac62d1af <= 'h0;
 Iacdfa68e9ab161a0e6c7e559b9954640 <= 'h0;
 Iedc0dfa42eaada48be02e65be4b39615 <= 'h0;
 Ib4fb78755c536a284004e41f584d99fb <= 'h0;
 I5156cd5e3f0fe53ad559b342c818f41a <= 'h0;
 I3cf816bf7fd922df289b13766e931e17 <= 'h0;
 Ibf2a30f91bd9050391913c02be7c8cad <= 'h0;
 Iea12e263d5883f93023d784884645969 <= 'h0;
 I550762460d0217d3c91c5112546b7929 <= 'h0;
 I0d8eaf22a03a0102d8bf7a53a7737943 <= 'h0;
 I8017a4f092179605074076e8b5690842 <= 'h0;
 I57160990c295512e2d98c301632c5120 <= 'h0;
 Id9f3f35bc6917416d6826d471f8ea441 <= 'h0;
 I6c9a443b704a7871ac13f164c1cdc88b <= 'h0;
 I76498f1e58ff35dc6153f76999f9f7a5 <= 'h0;
 I200025a860f318f6ff9aaf89b146d16f <= 'h0;
 I107ae84d631e3a9574b62f4fdfe56140 <= 'h0;
 Ief394bcabeb27c95f3dabe3d5c0bd643 <= 'h0;
 Ibc52ae3742f657ac6abefd988494c8a1 <= 'h0;
 I969ac5f2b8a9d6778300e3a91968ae4b <= 'h0;
 I3172be9cafebc7121994917ff35b25fb <= 'h0;
 I388e0d1c3f421d7522d6c0521538693e <= 'h0;
 I0fa0bdc864c6173b380c763cf3e794ba <= 'h0;
 I9d6dc129ad747412224b487c4973db3a <= 'h0;
 Ic1c5ee07ecd5c9fc9c2c1f9c33cdca08 <= 'h0;
 I1b2ba3544e2d26b40edbfaedf137812b <= 'h0;
 Ieb654d27e0306c60cd9eff05f4be76ca <= 'h0;
 I462601141783fc299a3b081023233a56 <= 'h0;
 I4e4e1489c822058cf54782c75c8d6996 <= 'h0;
 I361a262df08182fcb917b7aa7aa73465 <= 'h0;
 Ic8092176d020f45ae84ae72da9ea20a8 <= 'h0;
 I361a7201d61113929f346f8b22ac01ef <= 'h0;
 I616e26bab7d9ada350f152cce0ac3569 <= 'h0;
 I7cb33be246a06045ff19436b47ccfdca <= 'h0;
 Ic5aad088ddcc97dd7a3c8244a27a288e <= 'h0;
 I79c0e02b51ed3b20ca6de475189b6a48 <= 'h0;
 I059966174241b59374640dc43018c49c <= 'h0;
 I1b43d5eb392150245e2a303582b9226f <= 'h0;
 Icc5e7d899df8ec350f804c1f32b9fe72 <= 'h0;
 I2f8fbab2b60878195ae8b2e1c0ff1208 <= 'h0;
 I30e9a6bb0816599ede1e93a3091a572c <= 'h0;
 I815a192d304aedca5f772d6bd401ad3f <= 'h0;
 Id7c921ad25499d1e0bcf7dc1359e6b5d <= 'h0;
 I83ce7e2b4c276008c33a5703eba16572 <= 'h0;
 I96daacb3d66626af1c7b54c8be02a79b <= 'h0;
 I984e48eb72dcef91797c57289ba1322e <= 'h0;
 I8a0f063aab90c7f50f8eff7e3626483d <= 'h0;
 Ia49e2201160f9da0d475b16d22efcac1 <= 'h0;
 I59718bd7f0e7a0c9d63a038f2cb9d3eb <= 'h0;
 I7e703dc56c5c5604eb8e7ed32fd6ce78 <= 'h0;
 I1475899d2bf7a51aeae5168d5af0d548 <= 'h0;
 If3582b232dccd45a4f3c07514062003c <= 'h0;
 I79a9448f1efc66a407e2dcc243638e6f <= 'h0;
 I57fb6daf7238618d7ce10989a7f41025 <= 'h0;
 Ia677f2eaa008b296dc5eefdf680a2783 <= 'h0;
 I629cd82c8226c17eb439cd2ad664a3b7 <= 'h0;
 I181b85fc5fda9b5b99763bd8fa4a20b7 <= 'h0;
 Ida422d40a8abb52f4c78b63807f0ef16 <= 'h0;
 Ic91b7435580f54bb1e3ffa6ea1b21f69 <= 'h0;
 Id1651e9d3e909ddb1f3779b4129713fd <= 'h0;
 I470b1c602adb0b16c6b3a19133a97641 <= 'h0;
 I81c0a5fad7512ba9d8537018d6df2c23 <= 'h0;
 I0ea14616a599bd3f1c59dd57652ce967 <= 'h0;
 Ia6503d131655b73ae90b5553d116e92b <= 'h0;
 I2548ee3c3bf2a2eaa2ed541546e58c04 <= 'h0;
 I2c197653e4a8776ad3539f95aff27df5 <= 'h0;
 I0d6cfa3166445e1396871afad62fba40 <= 'h0;
 Ie597ab8c4dd174055b4bda8dbdec0dd3 <= 'h0;
 I46ee4c21a9801d95f803c4408dba7ea0 <= 'h0;
 I9426c6803cf8c7c6dbc422989eef5380 <= 'h0;
 I299fbb7b05d282681f0e9704b7818b0d <= 'h0;
 I947d66b22e42c68930e8bf7d1439a376 <= 'h0;
 I4e1752e19a8ec547211ca30f0e85c2d5 <= 'h0;
 I22715ee56f34e2c7cfdae2dd409ac653 <= 'h0;
 I85be91ab3b8a799d6681b90e6f56ad5e <= 'h0;
 Id2e3d5dfe5c8ec9128f5a719175c0f35 <= 'h0;
 I16d052ce0d66bc9f49489a124ccf6c69 <= 'h0;
 I0f1ace68f720dfcca74605ec277d0067 <= 'h0;
 I02f31af05294d3f39fe7c2f3a71a300a <= 'h0;
 Ia10e05a72a5d3c1e16b99510e94f6121 <= 'h0;
 I8b94c6d56df2d4a9a2adc2c7ccb8a0a9 <= 'h0;
 I8b6f4ea7a19f4b359aa01867c4502ccf <= 'h0;
 Id2add03142e6a3e5f4625082fbcc46ed <= 'h0;
 I323124e6fcbab5bdda4bd24c7b2a99c1 <= 'h0;
 Ib943a483749ffc791a5965ed0840bb0f <= 'h0;
 If379a89ad17fd061bf987e29aa713945 <= 'h0;
end
else
begin
 I72dd1fc26b57d741390612b9bcffab1d <=  I84ab01f2ac31304c9525b8983d34300d;
 I98c43e93e5f943a7b07ef09985f97014 <=  Iaf7ae8cb478fce9deaf537c13fa083cb;
 I434c16361fa147e26f4d2c4cc6d69150 <=  Idce9e18b46f498af68bbb108da7441bc;
 I9e87743bade1ee6fbfdd119cbdb0a3cb <=  Ie3954c25e29ea2d7e1340a59d3d7165f;
 I1e6255cf954cd5a58c52ff8e6a55bdbc <=  Iaa12f10c6588df5d8d8444c61b422c7c;
 I77a73f3832687dababc30666ac62d1af <=  I9851178cd4e84140f2c244f19c285e4a;
 Iacdfa68e9ab161a0e6c7e559b9954640 <=  I463cc1b85874882aadc9fa0ed9eb7816;
 Iedc0dfa42eaada48be02e65be4b39615 <=  I5249c4136a601a94d06d4955be304799;
 Ib4fb78755c536a284004e41f584d99fb <=  I9ce88b0e18af39ed6dc46db59a2bb78b;
 I5156cd5e3f0fe53ad559b342c818f41a <=  I3695c8773a6d76c02a9f8849ada96902;
 I3cf816bf7fd922df289b13766e931e17 <=  I4783f15f954421f7538cf39210bb44d5;
 Ibf2a30f91bd9050391913c02be7c8cad <=  Ia82244e3d80e219740368bab411242be;
 Iea12e263d5883f93023d784884645969 <=  Ib42df9a31ffd2cfc4a63cf95cf89c4d7;
 I550762460d0217d3c91c5112546b7929 <=  I752d56e6caa726064dc20d4eeda763a9;
 I0d8eaf22a03a0102d8bf7a53a7737943 <=  Ie339fd09fbad7893452b9a2f92d45932;
 I8017a4f092179605074076e8b5690842 <=  Ifd15d58d88de80f2cfc98c7f66f8f88d;
 I57160990c295512e2d98c301632c5120 <=  I994cd956aabc31d730d77d9b67bbc1db;
 Id9f3f35bc6917416d6826d471f8ea441 <=  Ie7086ba45d27b8fd48ad4dbbc1a6466b;
 I6c9a443b704a7871ac13f164c1cdc88b <=  I8539ebc561f7f4d823623b1f11255213;
 I76498f1e58ff35dc6153f76999f9f7a5 <=  Iedbd35fd7ebaf3787a08b0551ffb324e;
 I200025a860f318f6ff9aaf89b146d16f <=  I23df575a91b34e0a642bf679a74a747c;
 I107ae84d631e3a9574b62f4fdfe56140 <=  Icce0e60e3e31993ef47683a80567b1c4;
 Ief394bcabeb27c95f3dabe3d5c0bd643 <=  I172b401633d8844fcabdd4b980f46c73;
 Ibc52ae3742f657ac6abefd988494c8a1 <=  I71ed80b7d77c2a35edcefe9ce7db28af;
 I969ac5f2b8a9d6778300e3a91968ae4b <=  Ib1873b0070c00bfe5ed6fda941cfe95e;
 I3172be9cafebc7121994917ff35b25fb <=  I6db83f8bbff7cde9c9db248c02fd9358;
 I388e0d1c3f421d7522d6c0521538693e <=  If65d96ffe364426e1b90303ad323e7fb;
 I0fa0bdc864c6173b380c763cf3e794ba <=  I8e6c7979ddefa5e27581107ca2495e3e;
 I9d6dc129ad747412224b487c4973db3a <=  I161c2f4e7657ff863ec2a319ee8d21d5;
 Ic1c5ee07ecd5c9fc9c2c1f9c33cdca08 <=  Ic18bc04d9a02bccce383f311102a8b45;
 I1b2ba3544e2d26b40edbfaedf137812b <=  I8a118ced20140ec0f90f1f82161bd2c1;
 Ieb654d27e0306c60cd9eff05f4be76ca <=  I2b73e4b6134a9ca11b301452734741a1;
 I462601141783fc299a3b081023233a56 <=  Ie432836bf5a95e8dbb6de2c29d9ab058;
 I4e4e1489c822058cf54782c75c8d6996 <=  I8a777efecfec25782e29fd4e8f270490;
 I361a262df08182fcb917b7aa7aa73465 <=  I3ad4e40b398385b2c3a94cabd4736926;
 Ic8092176d020f45ae84ae72da9ea20a8 <=  Ifcd756c806de58265e16199e27f64e22;
 I361a7201d61113929f346f8b22ac01ef <=  Icac3b989b3d04d9c7a80d5eebcbb2027;
 I616e26bab7d9ada350f152cce0ac3569 <=  I806f4137adef04fa14f4c159fd47bb46;
 I7cb33be246a06045ff19436b47ccfdca <=  I6f6db1dfb50f19379683f16c549624b3;
 Ic5aad088ddcc97dd7a3c8244a27a288e <=  Ib26efe2924ee3c384a8f8b0f7f63e0f4;
 I79c0e02b51ed3b20ca6de475189b6a48 <=  I0a45d8f9e12c5234855b972d39246589;
 I059966174241b59374640dc43018c49c <=  I7a9fe30fbe486c1fd6d92b334f04a97b;
 I1b43d5eb392150245e2a303582b9226f <=  Ia5bc1b93ee0908ca26a967bc4720e5c3;
 Icc5e7d899df8ec350f804c1f32b9fe72 <=  I6cd39d0d0d14283cd00870fa8697cbe2;
 I2f8fbab2b60878195ae8b2e1c0ff1208 <=  Id33e3cde2a62f32d114a78300c2fdc1b;
 I30e9a6bb0816599ede1e93a3091a572c <=  I22f6c61d2512a383ecc57e2dac6e346a;
 I815a192d304aedca5f772d6bd401ad3f <=  I00b3081cd7dd077a53bdd7781b98fe6c;
 Id7c921ad25499d1e0bcf7dc1359e6b5d <=  Ibdf94fc4ee66c4af146968bf34ae4c0c;
 I83ce7e2b4c276008c33a5703eba16572 <=  Idadb48591ec328a331bdcf45e9156485;
 I96daacb3d66626af1c7b54c8be02a79b <=  I6315c142854dc3c1893bcb08b46bc739;
 I984e48eb72dcef91797c57289ba1322e <=  I362b966433fe2df6176a09951d0d88db;
 I8a0f063aab90c7f50f8eff7e3626483d <=  If210d0b145e2fd9cb2e1229c2c9c7a36;
 Ia49e2201160f9da0d475b16d22efcac1 <=  Ia133b750fb093f377556735adb4e3097;
 I59718bd7f0e7a0c9d63a038f2cb9d3eb <=  I6d2fcf19c79a538ec57aff56b8579def;
 I7e703dc56c5c5604eb8e7ed32fd6ce78 <=  If507c9ebcb1bc24a59ab4a00fc902d88;
 I1475899d2bf7a51aeae5168d5af0d548 <=  I70be43895e7446395ee6f209431a4b0e;
 If3582b232dccd45a4f3c07514062003c <=  Iec863324907434f27365ce30e0a3a636;
 I79a9448f1efc66a407e2dcc243638e6f <=  Ifdd6e035d37dc6a726502ea875e19bf2;
 I57fb6daf7238618d7ce10989a7f41025 <=  I0bac49aa5c179287d028c0bbe2f26646;
 Ia677f2eaa008b296dc5eefdf680a2783 <=  I676f1d8111d39181de6fb867fcc8aad9;
 I629cd82c8226c17eb439cd2ad664a3b7 <=  Ib6003647304cdf7e04f112ea1434d0c2;
 I181b85fc5fda9b5b99763bd8fa4a20b7 <=  I32f1ca64465d5ffd4c0abef6a0713795;
 Ida422d40a8abb52f4c78b63807f0ef16 <=  Iab2dbd174b3566d2eb0c32118a1d6ffc;
 Ic91b7435580f54bb1e3ffa6ea1b21f69 <=  I119a639a5c5243e5bbf6224fea9e0542;
 Id1651e9d3e909ddb1f3779b4129713fd <=  I51a744f6026f58a3ff9d47f7ad8441c7;
 I470b1c602adb0b16c6b3a19133a97641 <=  Ied88a6d77466adfacecc91792e092022;
 I81c0a5fad7512ba9d8537018d6df2c23 <=  I531565b08841415ba9f98966030529f2;
 I0ea14616a599bd3f1c59dd57652ce967 <=  I35641e3719c76fbc8621771af415d10f;
 Ia6503d131655b73ae90b5553d116e92b <=  I56baf72a394546e751edf096f5a87970;
 I2548ee3c3bf2a2eaa2ed541546e58c04 <=  I07ab92c9ad141c03101d587f00202c81;
 I2c197653e4a8776ad3539f95aff27df5 <=  I0143dfa3c201c85bdcce5739dee11814;
 I0d6cfa3166445e1396871afad62fba40 <=  Ie9a0ea695884198a9fd7e5de0a9f73d0;
 Ie597ab8c4dd174055b4bda8dbdec0dd3 <=  I0a066ff1810c068d1807dd5999880170;
 I46ee4c21a9801d95f803c4408dba7ea0 <=  I3d390c1d2a5df6decbc45bd682760b84;
 I9426c6803cf8c7c6dbc422989eef5380 <=  I0b1c32f0732334693986eea6aaee2b12;
 I299fbb7b05d282681f0e9704b7818b0d <=  Ifb9c5b70184594cb9f7961cb99c0d62e;
 I947d66b22e42c68930e8bf7d1439a376 <=  I105a0656b51423653fd7428001efa81f;
 I4e1752e19a8ec547211ca30f0e85c2d5 <=  Id9515c02ee595dc6ce4353decfbd2928;
 I22715ee56f34e2c7cfdae2dd409ac653 <=  Ib1d40c92e79f6562475204ba330c15e3;
 I85be91ab3b8a799d6681b90e6f56ad5e <=  Ief1a527fee16c6cb996ca3363d4713d8;
 Id2e3d5dfe5c8ec9128f5a719175c0f35 <=  I5c7ed7d4a522cf1e94035b3475d07240;
 I16d052ce0d66bc9f49489a124ccf6c69 <=  Ie59496301d7ef6565b69072f4530ceee;
 I0f1ace68f720dfcca74605ec277d0067 <=  I2d2b69150858f521850b9d71ee17acbf;
 I02f31af05294d3f39fe7c2f3a71a300a <=  I0556476f50843423945a3783fd5c9612;
 Ia10e05a72a5d3c1e16b99510e94f6121 <=  I34f9b6d4f00ab598a94274629c08e99c;
 I8b94c6d56df2d4a9a2adc2c7ccb8a0a9 <=  I2f16d9a27f31109e57160fbc03a98853;
 I8b6f4ea7a19f4b359aa01867c4502ccf <=  Ib19a79508dff3510b087cb2c1df176f9;
 Id2add03142e6a3e5f4625082fbcc46ed <=  I48ac3afb4f8b31f9aadc59aaf1a28a44;
 I323124e6fcbab5bdda4bd24c7b2a99c1 <=  Ia3bbc4519f9cd9651e10efaace317875;
 Ib943a483749ffc791a5965ed0840bb0f <=  I51118baae7de42e5f69f1a78d1ceccad;
 If379a89ad17fd061bf987e29aa713945 <=  I7aa491e6301b27435c2dadebe447b43a;
end
