//`include "GF2_LDPC_flogtanh_0x0000b_assign_inc.sv"
//always_comb begin
              I111cd97f7c5c13e18b528ffe1d1a871f['h00000] = 
          (!flogtanh_sel['h0000b]) ? 
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00000] : //%
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00001] ;
//end
//always_comb begin
              I111cd97f7c5c13e18b528ffe1d1a871f['h00001] = 
          (!flogtanh_sel['h0000b]) ? 
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00002] : //%
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00003] ;
//end
//always_comb begin
              I111cd97f7c5c13e18b528ffe1d1a871f['h00002] = 
          (!flogtanh_sel['h0000b]) ? 
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00004] : //%
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00005] ;
//end
//always_comb begin
              I111cd97f7c5c13e18b528ffe1d1a871f['h00003] = 
          (!flogtanh_sel['h0000b]) ? 
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00006] : //%
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00007] ;
//end
//always_comb begin
              I111cd97f7c5c13e18b528ffe1d1a871f['h00004] = 
          (!flogtanh_sel['h0000b]) ? 
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00008] : //%
                       I1a62004aa5608ddf7a551106f9a8a7ac['h00009] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00005] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0000a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00006] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0000c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00007] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0000e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00008] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00010] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00009] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00012] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0000a] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00014] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0000b] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00016] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0000c] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00018] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0000d] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0001a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0000e] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0001c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0000f] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0001e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00010] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00020] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00011] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00022] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00012] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00024] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00013] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00026] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00014] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00028] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00015] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0002a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00016] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0002c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00017] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0002e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00018] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00030] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00019] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00032] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0001a] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00034] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0001b] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00036] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0001c] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00038] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0001d] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0003a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0001e] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0003c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0001f] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0003e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00020] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00040] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00021] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00042] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00022] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00044] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00023] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00046] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00024] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00048] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00025] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0004a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00026] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0004c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00027] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0004e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00028] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00050] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00029] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00052] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0002a] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00054] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0002b] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00056] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0002c] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00058] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0002d] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0005a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0002e] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0005c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0002f] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0005e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00030] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00060] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00031] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00062] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00032] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00064] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00033] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00066] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00034] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00068] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00035] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0006a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00036] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0006c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00037] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0006e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00038] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00070] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00039] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00072] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0003a] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00074] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0003b] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00076] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0003c] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00078] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0003d] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0007a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0003e] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0007c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0003f] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0007e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00040] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00080] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00041] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00082] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00042] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00084] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00043] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00086] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00044] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00088] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00045] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0008a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00046] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0008c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00047] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0008e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00048] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00090] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00049] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00092] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0004a] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00094] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0004b] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00096] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0004c] =  I1a62004aa5608ddf7a551106f9a8a7ac['h00098] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0004d] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0009a] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0004e] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0009c] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0004f] =  I1a62004aa5608ddf7a551106f9a8a7ac['h0009e] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00050] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000a0] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00051] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000a2] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00052] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000a4] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00053] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000a6] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00054] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000a8] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00055] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000aa] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00056] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000ac] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00057] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000ae] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00058] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000b0] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00059] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000b2] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0005a] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000b4] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0005b] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000b6] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0005c] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000b8] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0005d] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000ba] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0005e] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000bc] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0005f] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000be] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00060] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000c0] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00061] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000c2] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00062] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000c4] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00063] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000c6] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00064] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000c8] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00065] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000ca] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00066] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000cc] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00067] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000ce] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00068] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000d0] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00069] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000d2] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0006a] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000d4] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0006b] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000d6] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0006c] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000d8] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0006d] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000da] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0006e] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000dc] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0006f] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000de] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00070] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000e0] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00071] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000e2] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00072] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000e4] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00073] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000e6] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00074] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000e8] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00075] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000ea] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00076] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000ec] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00077] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000ee] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00078] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000f0] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h00079] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000f2] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0007a] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000f4] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0007b] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000f6] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0007c] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000f8] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0007d] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000fa] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0007e] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000fc] ;
//end
//always_comb begin // 
               I111cd97f7c5c13e18b528ffe1d1a871f['h0007f] =  I1a62004aa5608ddf7a551106f9a8a7ac['h000fe] ;
//end
