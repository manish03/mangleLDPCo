parameter n_minus_m = 'd40;
parameter n_int = 'd208;
parameter m_int = 'd168;



parameter z_int = 'd4;



wire I994cbc6885873064963da8c47d5c2e70;
assign I994cbc6885873064963da8c47d5c2e70 = 
        y_nr_enc[1] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[8] ^ 
0; ///1



wire I2fac502186f123c8c0e1f8ba47db2460;
assign I2fac502186f123c8c0e1f8ba47db2460 = 
        y_nr_enc[14] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[37] ^ 
0; ///1



wire I70c11219ebff2b8a0392cc86b520018e;
assign I70c11219ebff2b8a0392cc86b520018e = 
        y_nr_enc[3] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[17] ^ 
0; ///1



wire I992e58b451deb7696487ddc59ef08da0;
assign I992e58b451deb7696487ddc59ef08da0 = 
        y_nr_enc[21] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire I395529ff583f9095755408ca5d85baff;
assign I395529ff583f9095755408ca5d85baff = 
        y_nr_enc[32] ^ 
        y_nr_enc[36] ^ 
        y_nr_enc[1] ^ 
0; ///1



wire I876a69bffa44696d92588ad80044cf95;
assign I876a69bffa44696d92588ad80044cf95 = 
        y_nr_enc[6] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[16] ^ 
0; ///1



wire I9592052279ccb8c52a1a8caac63a7c62;
assign I9592052279ccb8c52a1a8caac63a7c62 = 
        y_nr_enc[32] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[10] ^ 
0; ///1



wire Iefe1af67dd8717d051bffbc6f661d75d;
assign Iefe1af67dd8717d051bffbc6f661d75d = 
        y_nr_enc[18] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[25] ^ 
0; ///1



wire I2057df68f1ce06d8239dd8d9e7701a8b;
assign I2057df68f1ce06d8239dd8d9e7701a8b = 
        y_nr_enc[30] ^ 
        y_nr_enc[34] ^ 
        y_nr_enc[36] ^ 
0; ///1



    assign y_nr_p40 = 
I994cbc6885873064963da8c47d5c2e70 ^ 
I2fac502186f123c8c0e1f8ba47db2460 ^ 
I70c11219ebff2b8a0392cc86b520018e ^ 
I992e58b451deb7696487ddc59ef08da0 ^ 
I395529ff583f9095755408ca5d85baff ^ 
I876a69bffa44696d92588ad80044cf95 ^ 
I9592052279ccb8c52a1a8caac63a7c62 ^ 
Iefe1af67dd8717d051bffbc6f661d75d ^ 
I2057df68f1ce06d8239dd8d9e7701a8b ^ 
0; ///3



wire I3e129bded9d18251ce586cd98add20e7;
assign I3e129bded9d18251ce586cd98add20e7 = 
        y_nr_enc[2] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[9] ^ 
0; ///1



wire I1fd4089605a638510a157fd18eb32a5a;
assign I1fd4089605a638510a157fd18eb32a5a = 
        y_nr_enc[15] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[38] ^ 
0; ///1



wire I850eea9bb2cf06a59e25c6522c05c0c7;
assign I850eea9bb2cf06a59e25c6522c05c0c7 = 
        y_nr_enc[0] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[18] ^ 
0; ///1



wire Ia971e5d00ab87c820cd7f5ad1382fc23;
assign Ia971e5d00ab87c820cd7f5ad1382fc23 = 
        y_nr_enc[22] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire Id60c1aa86b3b01ae907eaa263261a3aa;
assign Id60c1aa86b3b01ae907eaa263261a3aa = 
        y_nr_enc[33] ^ 
        y_nr_enc[37] ^ 
        y_nr_enc[2] ^ 
0; ///1



wire I36f5910c0eb68590c91f46a77a76230d;
assign I36f5910c0eb68590c91f46a77a76230d = 
        y_nr_enc[7] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[17] ^ 
0; ///1



wire I2391cbda2dcefab98d2abc32bf35793c;
assign I2391cbda2dcefab98d2abc32bf35793c = 
        y_nr_enc[33] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[11] ^ 
0; ///1



wire Ic712fa03817f6be676254d76ef09e52d;
assign Ic712fa03817f6be676254d76ef09e52d = 
        y_nr_enc[19] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[26] ^ 
0; ///1



wire I39670247d92107aefaa13a4c66180c32;
assign I39670247d92107aefaa13a4c66180c32 = 
        y_nr_enc[31] ^ 
        y_nr_enc[35] ^ 
        y_nr_enc[37] ^ 
0; ///1



    assign y_nr_p41 = 
I3e129bded9d18251ce586cd98add20e7 ^ 
I1fd4089605a638510a157fd18eb32a5a ^ 
I850eea9bb2cf06a59e25c6522c05c0c7 ^ 
Ia971e5d00ab87c820cd7f5ad1382fc23 ^ 
Id60c1aa86b3b01ae907eaa263261a3aa ^ 
I36f5910c0eb68590c91f46a77a76230d ^ 
I2391cbda2dcefab98d2abc32bf35793c ^ 
Ic712fa03817f6be676254d76ef09e52d ^ 
I39670247d92107aefaa13a4c66180c32 ^ 
0; ///3



wire Iba029c82f31be025f157a5023c20d5cf;
assign Iba029c82f31be025f157a5023c20d5cf = 
        y_nr_enc[3] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[10] ^ 
0; ///1



wire If0913b8102a7eac0a62f9347b5048f10;
assign If0913b8102a7eac0a62f9347b5048f10 = 
        y_nr_enc[12] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[39] ^ 
0; ///1



wire I53525c14fee1e385ab3c926ca48c1128;
assign I53525c14fee1e385ab3c926ca48c1128 = 
        y_nr_enc[1] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[19] ^ 
0; ///1



wire I2fc248f9e649ef07db39d4d748995395;
assign I2fc248f9e649ef07db39d4d748995395 = 
        y_nr_enc[23] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire I2acf14e7b7a3008a3d20d0a98535015e;
assign I2acf14e7b7a3008a3d20d0a98535015e = 
        y_nr_enc[34] ^ 
        y_nr_enc[38] ^ 
        y_nr_enc[3] ^ 
0; ///1



wire I04057e7513ede3b836482c26caae4ede;
assign I04057e7513ede3b836482c26caae4ede = 
        y_nr_enc[4] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[18] ^ 
0; ///1



wire I8ec8397a7d3923824774a6212f8a387f;
assign I8ec8397a7d3923824774a6212f8a387f = 
        y_nr_enc[34] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[8] ^ 
0; ///1



wire I8f959f9964c8199a48f2bd1ccd5da3d2;
assign I8f959f9964c8199a48f2bd1ccd5da3d2 = 
        y_nr_enc[16] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[27] ^ 
0; ///1



wire I2ba0e30e00f77b16d8114e7a0b5d96a3;
assign I2ba0e30e00f77b16d8114e7a0b5d96a3 = 
        y_nr_enc[28] ^ 
        y_nr_enc[32] ^ 
        y_nr_enc[38] ^ 
0; ///1



    assign y_nr_p42 = 
Iba029c82f31be025f157a5023c20d5cf ^ 
If0913b8102a7eac0a62f9347b5048f10 ^ 
I53525c14fee1e385ab3c926ca48c1128 ^ 
I2fc248f9e649ef07db39d4d748995395 ^ 
I2acf14e7b7a3008a3d20d0a98535015e ^ 
I04057e7513ede3b836482c26caae4ede ^ 
I8ec8397a7d3923824774a6212f8a387f ^ 
I8f959f9964c8199a48f2bd1ccd5da3d2 ^ 
I2ba0e30e00f77b16d8114e7a0b5d96a3 ^ 
0; ///3



wire Idcf41bb2c1479baa76f8b3a2e8330df6;
assign Idcf41bb2c1479baa76f8b3a2e8330df6 = 
        y_nr_enc[0] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[11] ^ 
0; ///1



wire If3b5dfac0756d58b6da5978614646801;
assign If3b5dfac0756d58b6da5978614646801 = 
        y_nr_enc[13] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[36] ^ 
0; ///1



wire I2c39a9b52d070b51dd228f1a1c2747bb;
assign I2c39a9b52d070b51dd228f1a1c2747bb = 
        y_nr_enc[2] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[16] ^ 
0; ///1



wire I0be5ec80851ad6a5046700ca53b52337;
assign I0be5ec80851ad6a5046700ca53b52337 = 
        y_nr_enc[20] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire I16e3486a0bc5ba4a8dbfda3450be8316;
assign I16e3486a0bc5ba4a8dbfda3450be8316 = 
        y_nr_enc[35] ^ 
        y_nr_enc[39] ^ 
        y_nr_enc[0] ^ 
0; ///1



wire If42dba2a723efec3d8bc4700dc67933d;
assign If42dba2a723efec3d8bc4700dc67933d = 
        y_nr_enc[5] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[19] ^ 
0; ///1



wire I2cea417f39b000297083a01babf87045;
assign I2cea417f39b000297083a01babf87045 = 
        y_nr_enc[35] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[9] ^ 
0; ///1



wire I44fa537a6f8066c2ea9d4744a3b61969;
assign I44fa537a6f8066c2ea9d4744a3b61969 = 
        y_nr_enc[17] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[24] ^ 
0; ///1



wire I511872d7f5cd394da368a73796ceca4f;
assign I511872d7f5cd394da368a73796ceca4f = 
        y_nr_enc[29] ^ 
        y_nr_enc[33] ^ 
        y_nr_enc[39] ^ 
0; ///1



    assign y_nr_p43 = 
Idcf41bb2c1479baa76f8b3a2e8330df6 ^ 
If3b5dfac0756d58b6da5978614646801 ^ 
I2c39a9b52d070b51dd228f1a1c2747bb ^ 
I0be5ec80851ad6a5046700ca53b52337 ^ 
I16e3486a0bc5ba4a8dbfda3450be8316 ^ 
If42dba2a723efec3d8bc4700dc67933d ^ 
I2cea417f39b000297083a01babf87045 ^ 
I44fa537a6f8066c2ea9d4744a3b61969 ^ 
I511872d7f5cd394da368a73796ceca4f ^ 
0; ///3



wire I6e45115565a9662cc84c6067388f05aa;
assign I6e45115565a9662cc84c6067388f05aa = 
        y_nr_enc[1] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[8] ^ 
0; ///1



wire I68ca461b3d0eb4b6b6f41afa634d027b;
assign I68ca461b3d0eb4b6b6f41afa634d027b = 
        y_nr_enc[14] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[37] ^ 
0; ///1



wire I5b948982eec619889dee0777579ce449;
assign I5b948982eec619889dee0777579ce449 = 
        y_nr_enc[40] ^ 
0; ///1



    assign y_nr_p44 = 
I6e45115565a9662cc84c6067388f05aa ^ 
I68ca461b3d0eb4b6b6f41afa634d027b ^ 
I5b948982eec619889dee0777579ce449 ^ 
0; ///3



wire Ifa54e7ee30596fa80775c572c9217080;
assign Ifa54e7ee30596fa80775c572c9217080 = 
        y_nr_enc[2] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[9] ^ 
0; ///1



wire I6cfbce3ab9fbdda39ce970082acb4634;
assign I6cfbce3ab9fbdda39ce970082acb4634 = 
        y_nr_enc[15] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[38] ^ 
0; ///1



wire Icb30b911650ff935b32f81840f36b633;
assign Icb30b911650ff935b32f81840f36b633 = 
        y_nr_enc[41] ^ 
0; ///1



    assign y_nr_p45 = 
Ifa54e7ee30596fa80775c572c9217080 ^ 
I6cfbce3ab9fbdda39ce970082acb4634 ^ 
Icb30b911650ff935b32f81840f36b633 ^ 
0; ///3



wire Iea1e8bbfc64310269762d2aa735179e9;
assign Iea1e8bbfc64310269762d2aa735179e9 = 
        y_nr_enc[3] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[10] ^ 
0; ///1



wire Ie22a51a7271befd7ac2ad2b17ed57214;
assign Ie22a51a7271befd7ac2ad2b17ed57214 = 
        y_nr_enc[12] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[39] ^ 
0; ///1



wire Ic82c6d3d6ddabd90a7be9e27b3011628;
assign Ic82c6d3d6ddabd90a7be9e27b3011628 = 
        y_nr_enc[42] ^ 
0; ///1



    assign y_nr_p46 = 
Iea1e8bbfc64310269762d2aa735179e9 ^ 
Ie22a51a7271befd7ac2ad2b17ed57214 ^ 
Ic82c6d3d6ddabd90a7be9e27b3011628 ^ 
0; ///3



wire I4fea0065c281d915eeecd036641e63f8;
assign I4fea0065c281d915eeecd036641e63f8 = 
        y_nr_enc[0] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[11] ^ 
0; ///1



wire Iaee5b7677b303773b51dbbf3d52fd039;
assign Iaee5b7677b303773b51dbbf3d52fd039 = 
        y_nr_enc[13] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[36] ^ 
0; ///1



wire Iae8d787fb6550fcef4c10281e0eec3fc;
assign Iae8d787fb6550fcef4c10281e0eec3fc = 
        y_nr_enc[43] ^ 
0; ///1



    assign y_nr_p47 = 
I4fea0065c281d915eeecd036641e63f8 ^ 
Iaee5b7677b303773b51dbbf3d52fd039 ^ 
Iae8d787fb6550fcef4c10281e0eec3fc ^ 
0; ///3



wire I783a68caa51856938e8b99562710db73;
assign I783a68caa51856938e8b99562710db73 = 
        y_nr_enc[3] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[17] ^ 
0; ///1



wire Ie96d544bae373d562e8d030ec4de03e0;
assign Ie96d544bae373d562e8d030ec4de03e0 = 
        y_nr_enc[21] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire I6f14e012b9713a94c4f9ca64e9bda3bd;
assign I6f14e012b9713a94c4f9ca64e9bda3bd = 
        y_nr_enc[32] ^ 
        y_nr_enc[36] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p48 = 
I783a68caa51856938e8b99562710db73 ^ 
Ie96d544bae373d562e8d030ec4de03e0 ^ 
I6f14e012b9713a94c4f9ca64e9bda3bd ^ 
0; ///3



wire Ic4b097d301d6f96ce1fc0b09de4d6a23;
assign Ic4b097d301d6f96ce1fc0b09de4d6a23 = 
        y_nr_enc[0] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[18] ^ 
0; ///1



wire I9e0acdfd1ac1f4738406d11d73fcc65e;
assign I9e0acdfd1ac1f4738406d11d73fcc65e = 
        y_nr_enc[22] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire Ic5862f796199b32ba23d7e7df2c6f0ef;
assign Ic5862f796199b32ba23d7e7df2c6f0ef = 
        y_nr_enc[33] ^ 
        y_nr_enc[37] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p49 = 
Ic4b097d301d6f96ce1fc0b09de4d6a23 ^ 
I9e0acdfd1ac1f4738406d11d73fcc65e ^ 
Ic5862f796199b32ba23d7e7df2c6f0ef ^ 
0; ///3



wire I7364471fdbe4340497e3bad148a75393;
assign I7364471fdbe4340497e3bad148a75393 = 
        y_nr_enc[1] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[19] ^ 
0; ///1



wire Ib80c4cfd1fbd24337d41f77cfd03d088;
assign Ib80c4cfd1fbd24337d41f77cfd03d088 = 
        y_nr_enc[23] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire I05f8af669321e7bf504a2f3fb985b699;
assign I05f8af669321e7bf504a2f3fb985b699 = 
        y_nr_enc[34] ^ 
        y_nr_enc[38] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p50 = 
I7364471fdbe4340497e3bad148a75393 ^ 
Ib80c4cfd1fbd24337d41f77cfd03d088 ^ 
I05f8af669321e7bf504a2f3fb985b699 ^ 
0; ///3



wire I721d410b39d5c2e8cd992b4efa5d9842;
assign I721d410b39d5c2e8cd992b4efa5d9842 = 
        y_nr_enc[2] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[16] ^ 
0; ///1



wire I8fc1ba6df46b56693ee595f261d34130;
assign I8fc1ba6df46b56693ee595f261d34130 = 
        y_nr_enc[20] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire I4d9e5e86d2ae5b97a5a4da28348671fb;
assign I4d9e5e86d2ae5b97a5a4da28348671fb = 
        y_nr_enc[35] ^ 
        y_nr_enc[39] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p51 = 
I721d410b39d5c2e8cd992b4efa5d9842 ^ 
I8fc1ba6df46b56693ee595f261d34130 ^ 
I4d9e5e86d2ae5b97a5a4da28348671fb ^ 
0; ///3



wire I83a26de04f7c0bd283c0d4369f2f14da;
assign I83a26de04f7c0bd283c0d4369f2f14da = 
        y_nr_enc[4] ^ 
        y_nr_enc[10] ^ 
        y_nr_enc[18] ^ 
0; ///1



wire If8b44981a5a4afdcf9855caee86c210d;
assign If8b44981a5a4afdcf9855caee86c210d = 
        y_nr_enc[20] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire Id325ac8e45e72a368d21ba1ce755ef78;
assign Id325ac8e45e72a368d21ba1ce755ef78 = 
        y_nr_enc[34] ^ 
        y_nr_enc[36] ^ 
        y_nr_enc[40] ^ 
0; ///1



    assign y_nr_p52 = 
I83a26de04f7c0bd283c0d4369f2f14da ^ 
If8b44981a5a4afdcf9855caee86c210d ^ 
Id325ac8e45e72a368d21ba1ce755ef78 ^ 
0; ///3



wire I015f8243b630b6fda1e43cbf33cfb52e;
assign I015f8243b630b6fda1e43cbf33cfb52e = 
        y_nr_enc[5] ^ 
        y_nr_enc[11] ^ 
        y_nr_enc[19] ^ 
0; ///1



wire Ic8301fd1bfdf13a0dab0e02f900a6c99;
assign Ic8301fd1bfdf13a0dab0e02f900a6c99 = 
        y_nr_enc[21] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire Iadec5b0c6360d1491167c643ffa04ff6;
assign Iadec5b0c6360d1491167c643ffa04ff6 = 
        y_nr_enc[35] ^ 
        y_nr_enc[37] ^ 
        y_nr_enc[41] ^ 
0; ///1



    assign y_nr_p53 = 
I015f8243b630b6fda1e43cbf33cfb52e ^ 
Ic8301fd1bfdf13a0dab0e02f900a6c99 ^ 
Iadec5b0c6360d1491167c643ffa04ff6 ^ 
0; ///3



wire I4f1e9e3ba200348eac8910a857023db6;
assign I4f1e9e3ba200348eac8910a857023db6 = 
        y_nr_enc[6] ^ 
        y_nr_enc[8] ^ 
        y_nr_enc[16] ^ 
0; ///1



wire I68d72ba42f0f378959f36d6fd778c1e5;
assign I68d72ba42f0f378959f36d6fd778c1e5 = 
        y_nr_enc[22] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire I25eac8a2740f0128da2ba5a991b963a7;
assign I25eac8a2740f0128da2ba5a991b963a7 = 
        y_nr_enc[32] ^ 
        y_nr_enc[38] ^ 
        y_nr_enc[42] ^ 
0; ///1



    assign y_nr_p54 = 
I4f1e9e3ba200348eac8910a857023db6 ^ 
I68d72ba42f0f378959f36d6fd778c1e5 ^ 
I25eac8a2740f0128da2ba5a991b963a7 ^ 
0; ///3



wire I34187ea08b581b943a939d14dc1bf6aa;
assign I34187ea08b581b943a939d14dc1bf6aa = 
        y_nr_enc[7] ^ 
        y_nr_enc[9] ^ 
        y_nr_enc[17] ^ 
0; ///1



wire I67b9b8fd0d299610d169475adc91eccc;
assign I67b9b8fd0d299610d169475adc91eccc = 
        y_nr_enc[23] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire I46c81c9dba9d9e5eba8f7c1e2e344ac3;
assign I46c81c9dba9d9e5eba8f7c1e2e344ac3 = 
        y_nr_enc[33] ^ 
        y_nr_enc[39] ^ 
        y_nr_enc[43] ^ 
0; ///1



    assign y_nr_p55 = 
I34187ea08b581b943a939d14dc1bf6aa ^ 
I67b9b8fd0d299610d169475adc91eccc ^ 
I46c81c9dba9d9e5eba8f7c1e2e344ac3 ^ 
0; ///3



wire Iddbb8cadea75fe72c022210c810b8549;
assign Iddbb8cadea75fe72c022210c810b8549 = 
        y_nr_enc[3] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p56 = 
Iddbb8cadea75fe72c022210c810b8549 ^ 
0; ///3



wire Ia795dd007852ac6fc345e2dcf7354dcc;
assign Ia795dd007852ac6fc345e2dcf7354dcc = 
        y_nr_enc[0] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p57 = 
Ia795dd007852ac6fc345e2dcf7354dcc ^ 
0; ///3



wire Id7e208b8a84d5e8c925216f1830ab1dc;
assign Id7e208b8a84d5e8c925216f1830ab1dc = 
        y_nr_enc[1] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p58 = 
Id7e208b8a84d5e8c925216f1830ab1dc ^ 
0; ///3



wire I1d0080fa51dcaa096857cf8417eed37c;
assign I1d0080fa51dcaa096857cf8417eed37c = 
        y_nr_enc[2] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p59 = 
I1d0080fa51dcaa096857cf8417eed37c ^ 
0; ///3



wire I42937c2e177bda0fa8593fa2137b951f;
assign I42937c2e177bda0fa8593fa2137b951f = 
        y_nr_enc[3] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[22] ^ 
0; ///1



wire I3325e1a3557babba88703d757720bd23;
assign I3325e1a3557babba88703d757720bd23 = 
        y_nr_enc[31] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p60 = 
I42937c2e177bda0fa8593fa2137b951f ^ 
I3325e1a3557babba88703d757720bd23 ^ 
0; ///3



wire I2bcf445c4aef9bbe71c0cf1981ae879a;
assign I2bcf445c4aef9bbe71c0cf1981ae879a = 
        y_nr_enc[0] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[23] ^ 
0; ///1



wire I2feab319c9148ad7396c9a1182ffc420;
assign I2feab319c9148ad7396c9a1182ffc420 = 
        y_nr_enc[28] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p61 = 
I2bcf445c4aef9bbe71c0cf1981ae879a ^ 
I2feab319c9148ad7396c9a1182ffc420 ^ 
0; ///3



wire I5b6b64ad1bbf222f0073e92672bb0d83;
assign I5b6b64ad1bbf222f0073e92672bb0d83 = 
        y_nr_enc[1] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[20] ^ 
0; ///1



wire Ie230d9d3bec7814111d91fb18fff10cd;
assign Ie230d9d3bec7814111d91fb18fff10cd = 
        y_nr_enc[29] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p62 = 
I5b6b64ad1bbf222f0073e92672bb0d83 ^ 
Ie230d9d3bec7814111d91fb18fff10cd ^ 
0; ///3



wire I65a97bb5e117e4ea3f0142af00d7e97a;
assign I65a97bb5e117e4ea3f0142af00d7e97a = 
        y_nr_enc[2] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[21] ^ 
0; ///1



wire I8538dce6f44ae60e8ff829df755b7a73;
assign I8538dce6f44ae60e8ff829df755b7a73 = 
        y_nr_enc[30] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p63 = 
I65a97bb5e117e4ea3f0142af00d7e97a ^ 
I8538dce6f44ae60e8ff829df755b7a73 ^ 
0; ///3



wire I8fa493fbc2a4148584e8dbce01bdbc23;
assign I8fa493fbc2a4148584e8dbce01bdbc23 = 
        y_nr_enc[3] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire Idc5979a60a0d1e0451a5884e59da4269;
assign Idc5979a60a0d1e0451a5884e59da4269 = 
        y_nr_enc[36] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p64 = 
I8fa493fbc2a4148584e8dbce01bdbc23 ^ 
Idc5979a60a0d1e0451a5884e59da4269 ^ 
0; ///3



wire I7a3fa7bff345043428f4f4e3b975e75b;
assign I7a3fa7bff345043428f4f4e3b975e75b = 
        y_nr_enc[0] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire I3f593974c59abaed9b8083fb7788f057;
assign I3f593974c59abaed9b8083fb7788f057 = 
        y_nr_enc[37] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p65 = 
I7a3fa7bff345043428f4f4e3b975e75b ^ 
I3f593974c59abaed9b8083fb7788f057 ^ 
0; ///3



wire Id9221cfb0e0b336fbae90e9476a2a971;
assign Id9221cfb0e0b336fbae90e9476a2a971 = 
        y_nr_enc[1] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire I0b30a1bc77f2c147ce8aa12fd8df5bc2;
assign I0b30a1bc77f2c147ce8aa12fd8df5bc2 = 
        y_nr_enc[38] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p66 = 
Id9221cfb0e0b336fbae90e9476a2a971 ^ 
I0b30a1bc77f2c147ce8aa12fd8df5bc2 ^ 
0; ///3



wire If98dc167dcd322f1719476c9348409f1;
assign If98dc167dcd322f1719476c9348409f1 = 
        y_nr_enc[2] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire I8d242fc1fc6878d57ddcfefc46627097;
assign I8d242fc1fc6878d57ddcfefc46627097 = 
        y_nr_enc[39] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p67 = 
If98dc167dcd322f1719476c9348409f1 ^ 
I8d242fc1fc6878d57ddcfefc46627097 ^ 
0; ///3



wire I8dd8cab57144188f6e0773e1e5df58ce;
assign I8dd8cab57144188f6e0773e1e5df58ce = 
        y_nr_enc[5] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire Ia83c776387f608c5c3754055e4e0d19b;
assign Ia83c776387f608c5c3754055e4e0d19b = 
        y_nr_enc[47] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p68 = 
I8dd8cab57144188f6e0773e1e5df58ce ^ 
Ia83c776387f608c5c3754055e4e0d19b ^ 
0; ///3



wire I27c2fd00ed8a7b7439d6635ec4d266d9;
assign I27c2fd00ed8a7b7439d6635ec4d266d9 = 
        y_nr_enc[6] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire I269ab391add589034012f87db4bdddb8;
assign I269ab391add589034012f87db4bdddb8 = 
        y_nr_enc[44] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p69 = 
I27c2fd00ed8a7b7439d6635ec4d266d9 ^ 
I269ab391add589034012f87db4bdddb8 ^ 
0; ///3



wire Iaaa888522d4ca76f598b6a0c1983422a;
assign Iaaa888522d4ca76f598b6a0c1983422a = 
        y_nr_enc[7] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire I47e96683bf88c6cb83376141a8a5ab2f;
assign I47e96683bf88c6cb83376141a8a5ab2f = 
        y_nr_enc[45] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p70 = 
Iaaa888522d4ca76f598b6a0c1983422a ^ 
I47e96683bf88c6cb83376141a8a5ab2f ^ 
0; ///3



wire Ie9e355ee8fd99037b7a0bbe4a5f1c3af;
assign Ie9e355ee8fd99037b7a0bbe4a5f1c3af = 
        y_nr_enc[4] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire I05bbe6e423302fee1e4804f2bab58f75;
assign I05bbe6e423302fee1e4804f2bab58f75 = 
        y_nr_enc[46] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p71 = 
Ie9e355ee8fd99037b7a0bbe4a5f1c3af ^ 
I05bbe6e423302fee1e4804f2bab58f75 ^ 
0; ///3



wire Ia1c91fb831460d1c6785c3f5d18ec360;
assign Ia1c91fb831460d1c6785c3f5d18ec360 = 
        y_nr_enc[2] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p72 = 
Ia1c91fb831460d1c6785c3f5d18ec360 ^ 
0; ///3



wire I180cf5469404ec0d3aaaeb84eea26499;
assign I180cf5469404ec0d3aaaeb84eea26499 = 
        y_nr_enc[3] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p73 = 
I180cf5469404ec0d3aaaeb84eea26499 ^ 
0; ///3



wire Icf7aaea497def88eefb9921c4fbb9e5a;
assign Icf7aaea497def88eefb9921c4fbb9e5a = 
        y_nr_enc[0] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p74 = 
Icf7aaea497def88eefb9921c4fbb9e5a ^ 
0; ///3



wire I5c14ef919b15439738bf99616f369fc1;
assign I5c14ef919b15439738bf99616f369fc1 = 
        y_nr_enc[1] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p75 = 
I5c14ef919b15439738bf99616f369fc1 ^ 
0; ///3



wire Idaa3875ecebb798e7e3717e10b4b919c;
assign Idaa3875ecebb798e7e3717e10b4b919c = 
        y_nr_enc[7] ^ 
        y_nr_enc[33] ^ 
        y_nr_enc[41] ^ 
0; ///1



wire I1d64b5f50567a40e47d39838a2430dce;
assign I1d64b5f50567a40e47d39838a2430dce = 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p76 = 
Idaa3875ecebb798e7e3717e10b4b919c ^ 
I1d64b5f50567a40e47d39838a2430dce ^ 
0; ///3



wire I40fa3f3efaa5c05636ed9b28ad9cb4cc;
assign I40fa3f3efaa5c05636ed9b28ad9cb4cc = 
        y_nr_enc[4] ^ 
        y_nr_enc[34] ^ 
        y_nr_enc[42] ^ 
0; ///1



wire Ie39a04c5eb2c12c931f24ffd07f0c823;
assign Ie39a04c5eb2c12c931f24ffd07f0c823 = 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p77 = 
I40fa3f3efaa5c05636ed9b28ad9cb4cc ^ 
Ie39a04c5eb2c12c931f24ffd07f0c823 ^ 
0; ///3



wire If7994f23a88ab7918249a57fe68d1aed;
assign If7994f23a88ab7918249a57fe68d1aed = 
        y_nr_enc[5] ^ 
        y_nr_enc[35] ^ 
        y_nr_enc[43] ^ 
0; ///1



wire Ic2bb363719728467288480c88c2de30c;
assign Ic2bb363719728467288480c88c2de30c = 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p78 = 
If7994f23a88ab7918249a57fe68d1aed ^ 
Ic2bb363719728467288480c88c2de30c ^ 
0; ///3



wire I54c9487b4bf6274a0c842c5f48b57372;
assign I54c9487b4bf6274a0c842c5f48b57372 = 
        y_nr_enc[6] ^ 
        y_nr_enc[32] ^ 
        y_nr_enc[40] ^ 
0; ///1



wire I4343d69a86de24a2b7e25877091063d6;
assign I4343d69a86de24a2b7e25877091063d6 = 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p79 = 
I54c9487b4bf6274a0c842c5f48b57372 ^ 
I4343d69a86de24a2b7e25877091063d6 ^ 
0; ///3



wire I83ca53ce3c644409c24657bf1066f02a;
assign I83ca53ce3c644409c24657bf1066f02a = 
        y_nr_enc[3] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[24] ^ 
0; ///1



wire I3548442479fd1aebbee36894c23cc31b;
assign I3548442479fd1aebbee36894c23cc31b = 
        y_nr_enc[29] ^ 
0; ///1



    assign y_nr_p80 = 
I83ca53ce3c644409c24657bf1066f02a ^ 
I3548442479fd1aebbee36894c23cc31b ^ 
0; ///3



wire I6c38f79e06a784725ecbf2e01292c560;
assign I6c38f79e06a784725ecbf2e01292c560 = 
        y_nr_enc[0] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[25] ^ 
0; ///1



wire I5241d7f0ea17b4ade53110df329dd92f;
assign I5241d7f0ea17b4ade53110df329dd92f = 
        y_nr_enc[30] ^ 
0; ///1



    assign y_nr_p81 = 
I6c38f79e06a784725ecbf2e01292c560 ^ 
I5241d7f0ea17b4ade53110df329dd92f ^ 
0; ///3



wire I04585d1de8c679303e3fc3c4f6e49bbc;
assign I04585d1de8c679303e3fc3c4f6e49bbc = 
        y_nr_enc[1] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[26] ^ 
0; ///1



wire I395f7942d6b5587de0c31bc5e62df80c;
assign I395f7942d6b5587de0c31bc5e62df80c = 
        y_nr_enc[31] ^ 
0; ///1



    assign y_nr_p82 = 
I04585d1de8c679303e3fc3c4f6e49bbc ^ 
I395f7942d6b5587de0c31bc5e62df80c ^ 
0; ///3



wire Ib9a7d8a25e8613b233fe53dca55977bf;
assign Ib9a7d8a25e8613b233fe53dca55977bf = 
        y_nr_enc[2] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[27] ^ 
0; ///1



wire Icb45fc8caa92278663516903a1ade14f;
assign Icb45fc8caa92278663516903a1ade14f = 
        y_nr_enc[28] ^ 
0; ///1



    assign y_nr_p83 = 
Ib9a7d8a25e8613b233fe53dca55977bf ^ 
Icb45fc8caa92278663516903a1ade14f ^ 
0; ///3



wire Ia5660fac5b20fc46462eb24a518b52ad;
assign Ia5660fac5b20fc46462eb24a518b52ad = 
        y_nr_enc[3] ^ 
        y_nr_enc[28] ^ 
        y_nr_enc[38] ^ 
0; ///1



wire I68afcdc9b62948b07795f410996cdd4d;
assign I68afcdc9b62948b07795f410996cdd4d = 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p84 = 
Ia5660fac5b20fc46462eb24a518b52ad ^ 
I68afcdc9b62948b07795f410996cdd4d ^ 
0; ///3



wire I3f6f56151563dfdc84a6dcf118abab23;
assign I3f6f56151563dfdc84a6dcf118abab23 = 
        y_nr_enc[0] ^ 
        y_nr_enc[29] ^ 
        y_nr_enc[39] ^ 
0; ///1



wire I4683b8c397e9bd439ce6c7ce51768505;
assign I4683b8c397e9bd439ce6c7ce51768505 = 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p85 = 
I3f6f56151563dfdc84a6dcf118abab23 ^ 
I4683b8c397e9bd439ce6c7ce51768505 ^ 
0; ///3



wire Ifeab5e8f7acc3d83133f2ef19a8d8b63;
assign Ifeab5e8f7acc3d83133f2ef19a8d8b63 = 
        y_nr_enc[1] ^ 
        y_nr_enc[30] ^ 
        y_nr_enc[36] ^ 
0; ///1



wire I32632d4774f4bcaf13d81f00307bce78;
assign I32632d4774f4bcaf13d81f00307bce78 = 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p86 = 
Ifeab5e8f7acc3d83133f2ef19a8d8b63 ^ 
I32632d4774f4bcaf13d81f00307bce78 ^ 
0; ///3



wire I34fb25767233c3cee89f5c9d5cfcb237;
assign I34fb25767233c3cee89f5c9d5cfcb237 = 
        y_nr_enc[2] ^ 
        y_nr_enc[31] ^ 
        y_nr_enc[37] ^ 
0; ///1



wire If0195fbe9ce27a3bfb6b4ba74f9e98a6;
assign If0195fbe9ce27a3bfb6b4ba74f9e98a6 = 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p87 = 
I34fb25767233c3cee89f5c9d5cfcb237 ^ 
If0195fbe9ce27a3bfb6b4ba74f9e98a6 ^ 
0; ///3



wire Ie8378de324d09bea1c7dca1da1701818;
assign Ie8378de324d09bea1c7dca1da1701818 = 
        y_nr_enc[7] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p88 = 
Ie8378de324d09bea1c7dca1da1701818 ^ 
0; ///3



wire I5e8ee16f6a233f4fab248f41dca824f3;
assign I5e8ee16f6a233f4fab248f41dca824f3 = 
        y_nr_enc[4] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p89 = 
I5e8ee16f6a233f4fab248f41dca824f3 ^ 
0; ///3



wire I58b3695278fb37d733dacaba4d6dab8a;
assign I58b3695278fb37d733dacaba4d6dab8a = 
        y_nr_enc[5] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p90 = 
I58b3695278fb37d733dacaba4d6dab8a ^ 
0; ///3



wire Ied7345615b2c2a6da1191f107b5fc32d;
assign Ied7345615b2c2a6da1191f107b5fc32d = 
        y_nr_enc[6] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p91 = 
Ied7345615b2c2a6da1191f107b5fc32d ^ 
0; ///3



wire I783d115d823f18e427226c1a9c584629;
assign I783d115d823f18e427226c1a9c584629 = 
        y_nr_enc[3] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[34] ^ 
0; ///1



wire I759c20bf453b6b3267bf41dfa78f1b1b;
assign I759c20bf453b6b3267bf41dfa78f1b1b = 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p92 = 
I783d115d823f18e427226c1a9c584629 ^ 
I759c20bf453b6b3267bf41dfa78f1b1b ^ 
0; ///3



wire I14fed241f9bc3ea436ae883e5cecd350;
assign I14fed241f9bc3ea436ae883e5cecd350 = 
        y_nr_enc[0] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[35] ^ 
0; ///1



wire I7422232ccf20f912e0558bea4bed94c8;
assign I7422232ccf20f912e0558bea4bed94c8 = 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p93 = 
I14fed241f9bc3ea436ae883e5cecd350 ^ 
I7422232ccf20f912e0558bea4bed94c8 ^ 
0; ///3



wire I0242ed7821e573dccc9d95126d60f133;
assign I0242ed7821e573dccc9d95126d60f133 = 
        y_nr_enc[1] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[32] ^ 
0; ///1



wire I6e2d7831ed3a3c700fae32f4ce3b412a;
assign I6e2d7831ed3a3c700fae32f4ce3b412a = 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p94 = 
I0242ed7821e573dccc9d95126d60f133 ^ 
I6e2d7831ed3a3c700fae32f4ce3b412a ^ 
0; ///3



wire I97b5ba323cee8fdf6d26fd1aaf10c27d;
assign I97b5ba323cee8fdf6d26fd1aaf10c27d = 
        y_nr_enc[2] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[33] ^ 
0; ///1



wire I71ac6ddc03116ab4927dcb9d700b5ab7;
assign I71ac6ddc03116ab4927dcb9d700b5ab7 = 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p95 = 
I97b5ba323cee8fdf6d26fd1aaf10c27d ^ 
I71ac6ddc03116ab4927dcb9d700b5ab7 ^ 
0; ///3



wire If0ef4fd7e78e5c3ad88ecfc2819afdb7;
assign If0ef4fd7e78e5c3ad88ecfc2819afdb7 = 
        y_nr_enc[7] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[47] ^ 
0; ///1



wire I07052325724e5d7f3d18ee4a8932cc0b;
assign I07052325724e5d7f3d18ee4a8932cc0b = 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p96 = 
If0ef4fd7e78e5c3ad88ecfc2819afdb7 ^ 
I07052325724e5d7f3d18ee4a8932cc0b ^ 
0; ///3



wire I09c9635cb4f673f2bcbd56af308132ca;
assign I09c9635cb4f673f2bcbd56af308132ca = 
        y_nr_enc[4] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[44] ^ 
0; ///1



wire I62af0b0e7d6525bd6db456fdb3b8cd4b;
assign I62af0b0e7d6525bd6db456fdb3b8cd4b = 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p97 = 
I09c9635cb4f673f2bcbd56af308132ca ^ 
I62af0b0e7d6525bd6db456fdb3b8cd4b ^ 
0; ///3



wire I0846e43334feacce27262b2ae88f3652;
assign I0846e43334feacce27262b2ae88f3652 = 
        y_nr_enc[5] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[45] ^ 
0; ///1



wire I63e1595655b1012c655b72db7c18b99e;
assign I63e1595655b1012c655b72db7c18b99e = 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p98 = 
I0846e43334feacce27262b2ae88f3652 ^ 
I63e1595655b1012c655b72db7c18b99e ^ 
0; ///3



wire I69b387db12c0ba8c2ae044140263028a;
assign I69b387db12c0ba8c2ae044140263028a = 
        y_nr_enc[6] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[46] ^ 
0; ///1



wire Idecc6a323c06698f6acafcb9f185dbd6;
assign Idecc6a323c06698f6acafcb9f185dbd6 = 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p99 = 
I69b387db12c0ba8c2ae044140263028a ^ 
Idecc6a323c06698f6acafcb9f185dbd6 ^ 
0; ///3



wire I5348e033231c53f23e50ed0f3fd57387;
assign I5348e033231c53f23e50ed0f3fd57387 = 
        y_nr_enc[3] ^ 
        y_nr_enc[43] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p100 = 
I5348e033231c53f23e50ed0f3fd57387 ^ 
0; ///3



wire I7bf173000593c479ce07cd9718e2499b;
assign I7bf173000593c479ce07cd9718e2499b = 
        y_nr_enc[0] ^ 
        y_nr_enc[40] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p101 = 
I7bf173000593c479ce07cd9718e2499b ^ 
0; ///3



wire If042a8611c6b39451edd853e10593424;
assign If042a8611c6b39451edd853e10593424 = 
        y_nr_enc[1] ^ 
        y_nr_enc[41] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p102 = 
If042a8611c6b39451edd853e10593424 ^ 
0; ///3



wire I2ec30e3fb9e44de4dafff4be6dcb2435;
assign I2ec30e3fb9e44de4dafff4be6dcb2435 = 
        y_nr_enc[2] ^ 
        y_nr_enc[42] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p103 = 
I2ec30e3fb9e44de4dafff4be6dcb2435 ^ 
0; ///3



wire I552a0614d0064d7e9c0e67fe3d462598;
assign I552a0614d0064d7e9c0e67fe3d462598 = 
        y_nr_enc[7] ^ 
        y_nr_enc[38] ^ 
        y_nr_enc[44] ^ 
0; ///1



wire Ie31a3ac377fb81711e0d9d6a623e3bfa;
assign Ie31a3ac377fb81711e0d9d6a623e3bfa = 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p104 = 
I552a0614d0064d7e9c0e67fe3d462598 ^ 
Ie31a3ac377fb81711e0d9d6a623e3bfa ^ 
0; ///3



wire Ia0a3bb16f16bcb97403e7d4f1da97faf;
assign Ia0a3bb16f16bcb97403e7d4f1da97faf = 
        y_nr_enc[4] ^ 
        y_nr_enc[39] ^ 
        y_nr_enc[45] ^ 
0; ///1



wire Ia8c740bc63a78ce7385160458f4941bb;
assign Ia8c740bc63a78ce7385160458f4941bb = 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p105 = 
Ia0a3bb16f16bcb97403e7d4f1da97faf ^ 
Ia8c740bc63a78ce7385160458f4941bb ^ 
0; ///3



wire I3f3f24964631ff86486cb8ebe7ae804a;
assign I3f3f24964631ff86486cb8ebe7ae804a = 
        y_nr_enc[5] ^ 
        y_nr_enc[36] ^ 
        y_nr_enc[46] ^ 
0; ///1



wire I201cba1ca805deedd862b55b92ad33cc;
assign I201cba1ca805deedd862b55b92ad33cc = 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p106 = 
I3f3f24964631ff86486cb8ebe7ae804a ^ 
I201cba1ca805deedd862b55b92ad33cc ^ 
0; ///3



wire Ic02d10eb77626ab9989376b39126d8be;
assign Ic02d10eb77626ab9989376b39126d8be = 
        y_nr_enc[6] ^ 
        y_nr_enc[37] ^ 
        y_nr_enc[47] ^ 
0; ///1



wire Iaef7d50806bdd9e5821c10e9d7572566;
assign Iaef7d50806bdd9e5821c10e9d7572566 = 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p107 = 
Ic02d10eb77626ab9989376b39126d8be ^ 
Iaef7d50806bdd9e5821c10e9d7572566 ^ 
0; ///3



wire Id4b6cb8c33b1d59036203adfcc5672ed;
assign Id4b6cb8c33b1d59036203adfcc5672ed = 
        y_nr_enc[6] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[46] ^ 
0; ///1



wire I194f2f2342bfb13e6a9992c9e7995265;
assign I194f2f2342bfb13e6a9992c9e7995265 = 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p108 = 
Id4b6cb8c33b1d59036203adfcc5672ed ^ 
I194f2f2342bfb13e6a9992c9e7995265 ^ 
0; ///3



wire I3b6e24592cc80719b4dececa7a4e28cc;
assign I3b6e24592cc80719b4dececa7a4e28cc = 
        y_nr_enc[7] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[47] ^ 
0; ///1



wire I662239e5c4c519a9c31619149eaa7dfd;
assign I662239e5c4c519a9c31619149eaa7dfd = 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p109 = 
I3b6e24592cc80719b4dececa7a4e28cc ^ 
I662239e5c4c519a9c31619149eaa7dfd ^ 
0; ///3



wire I46ae162746bd979bb70a15b956cd2595;
assign I46ae162746bd979bb70a15b956cd2595 = 
        y_nr_enc[4] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[44] ^ 
0; ///1



wire I526a4856aa16e65b542805ae971e9be1;
assign I526a4856aa16e65b542805ae971e9be1 = 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p110 = 
I46ae162746bd979bb70a15b956cd2595 ^ 
I526a4856aa16e65b542805ae971e9be1 ^ 
0; ///3



wire I1732221ae74bdc2c54ec4c74a317a6ed;
assign I1732221ae74bdc2c54ec4c74a317a6ed = 
        y_nr_enc[5] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[45] ^ 
0; ///1



wire I74746a67d9f0f45605c46b9a8a5fe263;
assign I74746a67d9f0f45605c46b9a8a5fe263 = 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p111 = 
I1732221ae74bdc2c54ec4c74a317a6ed ^ 
I74746a67d9f0f45605c46b9a8a5fe263 ^ 
0; ///3



wire I8442ac3ae3b4a2c38ddf78d7a0990340;
assign I8442ac3ae3b4a2c38ddf78d7a0990340 = 
        y_nr_enc[0] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[30] ^ 
0; ///1



    assign y_nr_p112 = 
I8442ac3ae3b4a2c38ddf78d7a0990340 ^ 
0; ///3



wire I656a28386ecd524cdcd921b4b1115d12;
assign I656a28386ecd524cdcd921b4b1115d12 = 
        y_nr_enc[1] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[31] ^ 
0; ///1



    assign y_nr_p113 = 
I656a28386ecd524cdcd921b4b1115d12 ^ 
0; ///3



wire I3775e96b17d62750fa79474da0fab91d;
assign I3775e96b17d62750fa79474da0fab91d = 
        y_nr_enc[2] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[28] ^ 
0; ///1



    assign y_nr_p114 = 
I3775e96b17d62750fa79474da0fab91d ^ 
0; ///3



wire Ic44583baecc0ac0300afb12843594730;
assign Ic44583baecc0ac0300afb12843594730 = 
        y_nr_enc[3] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[29] ^ 
0; ///1



    assign y_nr_p115 = 
Ic44583baecc0ac0300afb12843594730 ^ 
0; ///3



wire I48f76466c82efdcdc7f8dce15170a938;
assign I48f76466c82efdcdc7f8dce15170a938 = 
        y_nr_enc[3] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[41] ^ 
0; ///1



    assign y_nr_p116 = 
I48f76466c82efdcdc7f8dce15170a938 ^ 
0; ///3



wire Id7a31089a62f31a38a03f60c7260f1c5;
assign Id7a31089a62f31a38a03f60c7260f1c5 = 
        y_nr_enc[0] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[42] ^ 
0; ///1



    assign y_nr_p117 = 
Id7a31089a62f31a38a03f60c7260f1c5 ^ 
0; ///3



wire Ia4289b88706434b24126468c6cc90a38;
assign Ia4289b88706434b24126468c6cc90a38 = 
        y_nr_enc[1] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[43] ^ 
0; ///1



    assign y_nr_p118 = 
Ia4289b88706434b24126468c6cc90a38 ^ 
0; ///3



wire I026e9e010674c4700dc146d51abf17c5;
assign I026e9e010674c4700dc146d51abf17c5 = 
        y_nr_enc[2] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[40] ^ 
0; ///1



    assign y_nr_p119 = 
I026e9e010674c4700dc146d51abf17c5 ^ 
0; ///3



wire If96ce0db664a443c59b3f5e77c92b0b4;
assign If96ce0db664a443c59b3f5e77c92b0b4 = 
        y_nr_enc[6] ^ 
        y_nr_enc[17] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p120 = 
If96ce0db664a443c59b3f5e77c92b0b4 ^ 
0; ///3



wire I4e1bcb771808ba3e7083e18a1c9fa44b;
assign I4e1bcb771808ba3e7083e18a1c9fa44b = 
        y_nr_enc[7] ^ 
        y_nr_enc[18] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p121 = 
I4e1bcb771808ba3e7083e18a1c9fa44b ^ 
0; ///3



wire I3ae53688f1ae7b6d991ff05e68177e84;
assign I3ae53688f1ae7b6d991ff05e68177e84 = 
        y_nr_enc[4] ^ 
        y_nr_enc[19] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p122 = 
I3ae53688f1ae7b6d991ff05e68177e84 ^ 
0; ///3



wire I9fa812ada94c4d9767e76b1b251e3f9c;
assign I9fa812ada94c4d9767e76b1b251e3f9c = 
        y_nr_enc[5] ^ 
        y_nr_enc[16] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p123 = 
I9fa812ada94c4d9767e76b1b251e3f9c ^ 
0; ///3



wire I9c8aa77496ca074b95ee44ca7e5b47c5;
assign I9c8aa77496ca074b95ee44ca7e5b47c5 = 
        y_nr_enc[0] ^ 
        y_nr_enc[34] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p124 = 
I9c8aa77496ca074b95ee44ca7e5b47c5 ^ 
0; ///3



wire Ic1ea390cb9f208be2940da3c25ac58e3;
assign Ic1ea390cb9f208be2940da3c25ac58e3 = 
        y_nr_enc[1] ^ 
        y_nr_enc[35] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p125 = 
Ic1ea390cb9f208be2940da3c25ac58e3 ^ 
0; ///3



wire I3e0b9e1e8b4ed8d6035305815d177106;
assign I3e0b9e1e8b4ed8d6035305815d177106 = 
        y_nr_enc[2] ^ 
        y_nr_enc[32] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p126 = 
I3e0b9e1e8b4ed8d6035305815d177106 ^ 
0; ///3



wire Id91f6d2f61111b53fd7a206db4a42623;
assign Id91f6d2f61111b53fd7a206db4a42623 = 
        y_nr_enc[3] ^ 
        y_nr_enc[33] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p127 = 
Id91f6d2f61111b53fd7a206db4a42623 ^ 
0; ///3



wire Id7c15cd8b9bd1567ba18287ca1f3c47d;
assign Id7c15cd8b9bd1567ba18287ca1f3c47d = 
        y_nr_enc[6] ^ 
        y_nr_enc[11] ^ 
0; ///1



    assign y_nr_p128 = 
Id7c15cd8b9bd1567ba18287ca1f3c47d ^ 
0; ///3



wire I1feeaebe0bae09f1e3cc862844af4118;
assign I1feeaebe0bae09f1e3cc862844af4118 = 
        y_nr_enc[7] ^ 
        y_nr_enc[8] ^ 
0; ///1



    assign y_nr_p129 = 
I1feeaebe0bae09f1e3cc862844af4118 ^ 
0; ///3



wire I464d94a17c1e2d73e5a78d5b93ff65bb;
assign I464d94a17c1e2d73e5a78d5b93ff65bb = 
        y_nr_enc[4] ^ 
        y_nr_enc[9] ^ 
0; ///1



    assign y_nr_p130 = 
I464d94a17c1e2d73e5a78d5b93ff65bb ^ 
0; ///3



wire I5d27f5a5a9f1c9b37abec760849f684d;
assign I5d27f5a5a9f1c9b37abec760849f684d = 
        y_nr_enc[5] ^ 
        y_nr_enc[10] ^ 
0; ///1



    assign y_nr_p131 = 
I5d27f5a5a9f1c9b37abec760849f684d ^ 
0; ///3



wire Ifd00fbc5ee7d9ede693f547cbfcf0783;
assign Ifd00fbc5ee7d9ede693f547cbfcf0783 = 
        y_nr_enc[3] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[22] ^ 
0; ///1



    assign y_nr_p132 = 
Ifd00fbc5ee7d9ede693f547cbfcf0783 ^ 
0; ///3



wire Ifdf5b6ae37f51d978e052dea4d3b1042;
assign Ifdf5b6ae37f51d978e052dea4d3b1042 = 
        y_nr_enc[0] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[23] ^ 
0; ///1



    assign y_nr_p133 = 
Ifdf5b6ae37f51d978e052dea4d3b1042 ^ 
0; ///3



wire I5aaaa1bd0f8f9a8e8f110f9af1019778;
assign I5aaaa1bd0f8f9a8e8f110f9af1019778 = 
        y_nr_enc[1] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[20] ^ 
0; ///1



    assign y_nr_p134 = 
I5aaaa1bd0f8f9a8e8f110f9af1019778 ^ 
0; ///3



wire I65d3fa7565b7736c71b79f801a9160ae;
assign I65d3fa7565b7736c71b79f801a9160ae = 
        y_nr_enc[2] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[21] ^ 
0; ///1



    assign y_nr_p135 = 
I65d3fa7565b7736c71b79f801a9160ae ^ 
0; ///3



wire Iacb7b499942da0f999c4db02b0f000d1;
assign Iacb7b499942da0f999c4db02b0f000d1 = 
        y_nr_enc[6] ^ 
        y_nr_enc[11] ^ 
        y_nr_enc[36] ^ 
0; ///1



    assign y_nr_p136 = 
Iacb7b499942da0f999c4db02b0f000d1 ^ 
0; ///3



wire Ie4b25c598547ad2754e5e37c4f6f270e;
assign Ie4b25c598547ad2754e5e37c4f6f270e = 
        y_nr_enc[7] ^ 
        y_nr_enc[8] ^ 
        y_nr_enc[37] ^ 
0; ///1



    assign y_nr_p137 = 
Ie4b25c598547ad2754e5e37c4f6f270e ^ 
0; ///3



wire I94b1799c5d2b8c6a303c1b1f233318f7;
assign I94b1799c5d2b8c6a303c1b1f233318f7 = 
        y_nr_enc[4] ^ 
        y_nr_enc[9] ^ 
        y_nr_enc[38] ^ 
0; ///1



    assign y_nr_p138 = 
I94b1799c5d2b8c6a303c1b1f233318f7 ^ 
0; ///3



wire Iff94a0966ab1d59373ec663f95b3b404;
assign Iff94a0966ab1d59373ec663f95b3b404 = 
        y_nr_enc[5] ^ 
        y_nr_enc[10] ^ 
        y_nr_enc[39] ^ 
0; ///1



    assign y_nr_p139 = 
Iff94a0966ab1d59373ec663f95b3b404 ^ 
0; ///3



wire I736e461f587ce87b578557c14a90ad27;
assign I736e461f587ce87b578557c14a90ad27 = 
        y_nr_enc[0] ^ 
        y_nr_enc[20] ^ 
0; ///1



    assign y_nr_p140 = 
I736e461f587ce87b578557c14a90ad27 ^ 
0; ///3



wire I9f7fc1ad1d5682b21bf08687b898d2dc;
assign I9f7fc1ad1d5682b21bf08687b898d2dc = 
        y_nr_enc[1] ^ 
        y_nr_enc[21] ^ 
0; ///1



    assign y_nr_p141 = 
I9f7fc1ad1d5682b21bf08687b898d2dc ^ 
0; ///3



wire I060921c8d21c334264eca4a5055c607e;
assign I060921c8d21c334264eca4a5055c607e = 
        y_nr_enc[2] ^ 
        y_nr_enc[22] ^ 
0; ///1



    assign y_nr_p142 = 
I060921c8d21c334264eca4a5055c607e ^ 
0; ///3



wire Ia7f663e3e88aa14c60e73f1151d58c77;
assign Ia7f663e3e88aa14c60e73f1151d58c77 = 
        y_nr_enc[3] ^ 
        y_nr_enc[23] ^ 
0; ///1



    assign y_nr_p143 = 
Ia7f663e3e88aa14c60e73f1151d58c77 ^ 
0; ///3



wire Id304ae830be08dfa5907350ed057f747;
assign Id304ae830be08dfa5907350ed057f747 = 
        y_nr_enc[9] ^ 
        y_nr_enc[31] ^ 
        y_nr_enc[48] ^ 
0; ///1



wire I4dba19d3dd5f39e88448eb13d38a7aa7;
assign I4dba19d3dd5f39e88448eb13d38a7aa7 = 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p144 = 
Id304ae830be08dfa5907350ed057f747 ^ 
I4dba19d3dd5f39e88448eb13d38a7aa7 ^ 
0; ///3



wire If25082bb5be2d557b83d46d899889cd3;
assign If25082bb5be2d557b83d46d899889cd3 = 
        y_nr_enc[10] ^ 
        y_nr_enc[28] ^ 
        y_nr_enc[49] ^ 
0; ///1



wire I77d94e0b0b74acc2095b1fc234cf2e80;
assign I77d94e0b0b74acc2095b1fc234cf2e80 = 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p145 = 
If25082bb5be2d557b83d46d899889cd3 ^ 
I77d94e0b0b74acc2095b1fc234cf2e80 ^ 
0; ///3



wire I6d697a13151c7d2980d3e0491e0a765a;
assign I6d697a13151c7d2980d3e0491e0a765a = 
        y_nr_enc[11] ^ 
        y_nr_enc[29] ^ 
        y_nr_enc[50] ^ 
0; ///1



wire Id8e54e9611355553f486a0e81e94936d;
assign Id8e54e9611355553f486a0e81e94936d = 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p146 = 
I6d697a13151c7d2980d3e0491e0a765a ^ 
Id8e54e9611355553f486a0e81e94936d ^ 
0; ///3



wire I8646f5f0671f46772414ad5876d2dec3;
assign I8646f5f0671f46772414ad5876d2dec3 = 
        y_nr_enc[8] ^ 
        y_nr_enc[30] ^ 
        y_nr_enc[51] ^ 
0; ///1



wire Icec96b5572185a51ff7503be19c93aca;
assign Icec96b5572185a51ff7503be19c93aca = 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p147 = 
I8646f5f0671f46772414ad5876d2dec3 ^ 
Icec96b5572185a51ff7503be19c93aca ^ 
0; ///3



wire I132094289f37c45eb195cc1f9018ec2f;
assign I132094289f37c45eb195cc1f9018ec2f = 
        y_nr_enc[0] ^ 
        y_nr_enc[27] ^ 
0; ///1



    assign y_nr_p148 = 
I132094289f37c45eb195cc1f9018ec2f ^ 
0; ///3



wire I957fb739fc10dada866bb153a7172c8b;
assign I957fb739fc10dada866bb153a7172c8b = 
        y_nr_enc[1] ^ 
        y_nr_enc[24] ^ 
0; ///1



    assign y_nr_p149 = 
I957fb739fc10dada866bb153a7172c8b ^ 
0; ///3



wire I73d2d279b02f97616af81893206308c5;
assign I73d2d279b02f97616af81893206308c5 = 
        y_nr_enc[2] ^ 
        y_nr_enc[25] ^ 
0; ///1



    assign y_nr_p150 = 
I73d2d279b02f97616af81893206308c5 ^ 
0; ///3



wire Ibc77ea6f27dd8b748f438f63b9687dc8;
assign Ibc77ea6f27dd8b748f438f63b9687dc8 = 
        y_nr_enc[3] ^ 
        y_nr_enc[26] ^ 
0; ///1



    assign y_nr_p151 = 
Ibc77ea6f27dd8b748f438f63b9687dc8 ^ 
0; ///3



wire I3431a1e2c7bb8260298394d9c76259bc;
assign I3431a1e2c7bb8260298394d9c76259bc = 
        y_nr_enc[6] ^ 
        y_nr_enc[9] ^ 
        y_nr_enc[23] ^ 
0; ///1



    assign y_nr_p152 = 
I3431a1e2c7bb8260298394d9c76259bc ^ 
0; ///3



wire Ib1f0a14b550ef15e5b8dc693357f66cc;
assign Ib1f0a14b550ef15e5b8dc693357f66cc = 
        y_nr_enc[7] ^ 
        y_nr_enc[10] ^ 
        y_nr_enc[20] ^ 
0; ///1



    assign y_nr_p153 = 
Ib1f0a14b550ef15e5b8dc693357f66cc ^ 
0; ///3



wire I1d61c6295cdba37ea84b8aea65eef2f2;
assign I1d61c6295cdba37ea84b8aea65eef2f2 = 
        y_nr_enc[4] ^ 
        y_nr_enc[11] ^ 
        y_nr_enc[21] ^ 
0; ///1



    assign y_nr_p154 = 
I1d61c6295cdba37ea84b8aea65eef2f2 ^ 
0; ///3



wire I21f88f49ed27f1cdf8dbef0d20922d39;
assign I21f88f49ed27f1cdf8dbef0d20922d39 = 
        y_nr_enc[5] ^ 
        y_nr_enc[8] ^ 
        y_nr_enc[22] ^ 
0; ///1



    assign y_nr_p155 = 
I21f88f49ed27f1cdf8dbef0d20922d39 ^ 
0; ///3



wire I8ad69370aae0f8055229dfbf0a64dfba;
assign I8ad69370aae0f8055229dfbf0a64dfba = 
        y_nr_enc[2] ^ 
        y_nr_enc[16] ^ 
0; ///1



    assign y_nr_p156 = 
I8ad69370aae0f8055229dfbf0a64dfba ^ 
0; ///3



wire Id1c589c3a43d58652a0db23fb9f88a0f;
assign Id1c589c3a43d58652a0db23fb9f88a0f = 
        y_nr_enc[3] ^ 
        y_nr_enc[17] ^ 
0; ///1



    assign y_nr_p157 = 
Id1c589c3a43d58652a0db23fb9f88a0f ^ 
0; ///3



wire I0a55590d50cb08a17a2a1af2aca93627;
assign I0a55590d50cb08a17a2a1af2aca93627 = 
        y_nr_enc[0] ^ 
        y_nr_enc[18] ^ 
0; ///1



    assign y_nr_p158 = 
I0a55590d50cb08a17a2a1af2aca93627 ^ 
0; ///3



wire I5d0c660ce8de5d8020cc65fcbb8b7eaa;
assign I5d0c660ce8de5d8020cc65fcbb8b7eaa = 
        y_nr_enc[1] ^ 
        y_nr_enc[19] ^ 
0; ///1



    assign y_nr_p159 = 
I5d0c660ce8de5d8020cc65fcbb8b7eaa ^ 
0; ///3



wire Iaaf46a284a83c2d3536e9c488bdd422b;
assign Iaaf46a284a83c2d3536e9c488bdd422b = 
        y_nr_enc[11] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire I622215b8d6537e1c8401acc8adeecd72;
assign I622215b8d6537e1c8401acc8adeecd72 = 
        y_nr_enc[36] ^ 
0; ///1



    assign y_nr_p160 = 
Iaaf46a284a83c2d3536e9c488bdd422b ^ 
I622215b8d6537e1c8401acc8adeecd72 ^ 
0; ///3



wire Iedb1d669307cb8c6f388817d981bd2b3;
assign Iedb1d669307cb8c6f388817d981bd2b3 = 
        y_nr_enc[8] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire I4009422c3627f7d7c61ae8920ce244a2;
assign I4009422c3627f7d7c61ae8920ce244a2 = 
        y_nr_enc[37] ^ 
0; ///1



    assign y_nr_p161 = 
Iedb1d669307cb8c6f388817d981bd2b3 ^ 
I4009422c3627f7d7c61ae8920ce244a2 ^ 
0; ///3



wire I20af0bd615898f2d09f249e8fad8744d;
assign I20af0bd615898f2d09f249e8fad8744d = 
        y_nr_enc[9] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire I91dc73be3f02f86c52aa7ed127aeaef7;
assign I91dc73be3f02f86c52aa7ed127aeaef7 = 
        y_nr_enc[38] ^ 
0; ///1



    assign y_nr_p162 = 
I20af0bd615898f2d09f249e8fad8744d ^ 
I91dc73be3f02f86c52aa7ed127aeaef7 ^ 
0; ///3



wire I2e1882ff44183a235dbc9458f5cc12d5;
assign I2e1882ff44183a235dbc9458f5cc12d5 = 
        y_nr_enc[10] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire I34df82ee57ca08021ad8d82cb7c51a39;
assign I34df82ee57ca08021ad8d82cb7c51a39 = 
        y_nr_enc[39] ^ 
0; ///1



    assign y_nr_p163 = 
I2e1882ff44183a235dbc9458f5cc12d5 ^ 
I34df82ee57ca08021ad8d82cb7c51a39 ^ 
0; ///3



wire I2cc04871cf7db5c113f63d9c1532ada4;
assign I2cc04871cf7db5c113f63d9c1532ada4 = 
        y_nr_enc[6] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p164 = 
I2cc04871cf7db5c113f63d9c1532ada4 ^ 
0; ///3



wire I5b21f49ef448970447352bcbb313b12e;
assign I5b21f49ef448970447352bcbb313b12e = 
        y_nr_enc[7] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p165 = 
I5b21f49ef448970447352bcbb313b12e ^ 
0; ///3



wire I39a0f30431bb80f07ad12103678d3491;
assign I39a0f30431bb80f07ad12103678d3491 = 
        y_nr_enc[4] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p166 = 
I39a0f30431bb80f07ad12103678d3491 ^ 
0; ///3



wire I493cb21c246bde0f5efd8aff89a1a1df;
assign I493cb21c246bde0f5efd8aff89a1a1df = 
        y_nr_enc[5] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p167 = 
I493cb21c246bde0f5efd8aff89a1a1df ^ 
0; ///3



wire I3bf088d9a090a28b32b7254bf6493fd0;
assign I3bf088d9a090a28b32b7254bf6493fd0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p168 = 
I3bf088d9a090a28b32b7254bf6493fd0 ^ 
0; ///3



wire Ib4996da5c27e98c3c70fb53153bf75c0;
assign Ib4996da5c27e98c3c70fb53153bf75c0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p169 = 
Ib4996da5c27e98c3c70fb53153bf75c0 ^ 
0; ///3



wire I5d7e01b038448c2c9c9aa34166eda5f0;
assign I5d7e01b038448c2c9c9aa34166eda5f0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p170 = 
I5d7e01b038448c2c9c9aa34166eda5f0 ^ 
0; ///3



wire Iebc5ba3282701ab0ab1349389109b4a0;
assign Iebc5ba3282701ab0ab1349389109b4a0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p171 = 
Iebc5ba3282701ab0ab1349389109b4a0 ^ 
0; ///3



wire Iaa24ca8ed0a2d257fc697e5ff95e028a;
assign Iaa24ca8ed0a2d257fc697e5ff95e028a = 
        y_nr_enc[8] ^ 
        y_nr_enc[28] ^ 
        y_nr_enc[43] ^ 
0; ///1



    assign y_nr_p172 = 
Iaa24ca8ed0a2d257fc697e5ff95e028a ^ 
0; ///3



wire I08b68c9f4ae1975a8644d215bdb27fbf;
assign I08b68c9f4ae1975a8644d215bdb27fbf = 
        y_nr_enc[9] ^ 
        y_nr_enc[29] ^ 
        y_nr_enc[40] ^ 
0; ///1



    assign y_nr_p173 = 
I08b68c9f4ae1975a8644d215bdb27fbf ^ 
0; ///3



wire I037045883ea9fdc4f01f5366ac14a79c;
assign I037045883ea9fdc4f01f5366ac14a79c = 
        y_nr_enc[10] ^ 
        y_nr_enc[30] ^ 
        y_nr_enc[41] ^ 
0; ///1



    assign y_nr_p174 = 
I037045883ea9fdc4f01f5366ac14a79c ^ 
0; ///3



wire Iaacd417ffb9927da6d2d261f79e332f3;
assign Iaacd417ffb9927da6d2d261f79e332f3 = 
        y_nr_enc[11] ^ 
        y_nr_enc[31] ^ 
        y_nr_enc[42] ^ 
0; ///1



    assign y_nr_p175 = 
Iaacd417ffb9927da6d2d261f79e332f3 ^ 
0; ///3



wire I2a8ea7b7aa9c2d83921c19d79068bb41;
assign I2a8ea7b7aa9c2d83921c19d79068bb41 = 
        y_nr_enc[3] ^ 
        y_nr_enc[49] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p176 = 
I2a8ea7b7aa9c2d83921c19d79068bb41 ^ 
0; ///3



wire I0115b1811fe5f13c3b531f2125427c5a;
assign I0115b1811fe5f13c3b531f2125427c5a = 
        y_nr_enc[0] ^ 
        y_nr_enc[50] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p177 = 
I0115b1811fe5f13c3b531f2125427c5a ^ 
0; ///3



wire Ia75912167f884f97790ca7891f0c8a24;
assign Ia75912167f884f97790ca7891f0c8a24 = 
        y_nr_enc[1] ^ 
        y_nr_enc[51] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p178 = 
Ia75912167f884f97790ca7891f0c8a24 ^ 
0; ///3



wire Ifb16c5b88ecd639e3b9378cb25e20b8a;
assign Ifb16c5b88ecd639e3b9378cb25e20b8a = 
        y_nr_enc[2] ^ 
        y_nr_enc[48] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p179 = 
Ifb16c5b88ecd639e3b9378cb25e20b8a ^ 
0; ///3



wire Ia84c83fdf902c5d802c27e6648b910cb;
assign Ia84c83fdf902c5d802c27e6648b910cb = 
        y_nr_enc[5] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p180 = 
Ia84c83fdf902c5d802c27e6648b910cb ^ 
0; ///3



wire I9adb83fe9a66bdfb27d45c3b6e973bd1;
assign I9adb83fe9a66bdfb27d45c3b6e973bd1 = 
        y_nr_enc[6] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p181 = 
I9adb83fe9a66bdfb27d45c3b6e973bd1 ^ 
0; ///3



wire If89e677c2f7e810bb36bb93276186928;
assign If89e677c2f7e810bb36bb93276186928 = 
        y_nr_enc[7] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p182 = 
If89e677c2f7e810bb36bb93276186928 ^ 
0; ///3



wire Ie2570a4283d5fc1e46aba92d5ab4dca6;
assign Ie2570a4283d5fc1e46aba92d5ab4dca6 = 
        y_nr_enc[4] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p183 = 
Ie2570a4283d5fc1e46aba92d5ab4dca6 ^ 
0; ///3



wire I23a380ce0596fbc938eef5a78c9b89ba;
assign I23a380ce0596fbc938eef5a78c9b89ba = 
        y_nr_enc[0] ^ 
        y_nr_enc[10] ^ 
        y_nr_enc[30] ^ 
0; ///1



    assign y_nr_p184 = 
I23a380ce0596fbc938eef5a78c9b89ba ^ 
0; ///3



wire Id393725bab01e3f363f5038ba5f70e1a;
assign Id393725bab01e3f363f5038ba5f70e1a = 
        y_nr_enc[1] ^ 
        y_nr_enc[11] ^ 
        y_nr_enc[31] ^ 
0; ///1



    assign y_nr_p185 = 
Id393725bab01e3f363f5038ba5f70e1a ^ 
0; ///3



wire I3c1797b1c25c91fd41cf42dc2d220a71;
assign I3c1797b1c25c91fd41cf42dc2d220a71 = 
        y_nr_enc[2] ^ 
        y_nr_enc[8] ^ 
        y_nr_enc[28] ^ 
0; ///1



    assign y_nr_p186 = 
I3c1797b1c25c91fd41cf42dc2d220a71 ^ 
0; ///3



wire I9c917b1f6dfada02da562816e2d7631a;
assign I9c917b1f6dfada02da562816e2d7631a = 
        y_nr_enc[3] ^ 
        y_nr_enc[9] ^ 
        y_nr_enc[29] ^ 
0; ///1



    assign y_nr_p187 = 
I9c917b1f6dfada02da562816e2d7631a ^ 
0; ///3



wire I0bcbe782440e3c5b310a9f50a0dee451;
assign I0bcbe782440e3c5b310a9f50a0dee451 = 
        y_nr_enc[43] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p188 = 
I0bcbe782440e3c5b310a9f50a0dee451 ^ 
0; ///3



wire Iadd3239fa89efd2de8387c69b78c8a3a;
assign Iadd3239fa89efd2de8387c69b78c8a3a = 
        y_nr_enc[40] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p189 = 
Iadd3239fa89efd2de8387c69b78c8a3a ^ 
0; ///3



wire Ic39ac97e1121894b3efbba7ddd49e96f;
assign Ic39ac97e1121894b3efbba7ddd49e96f = 
        y_nr_enc[41] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p190 = 
Ic39ac97e1121894b3efbba7ddd49e96f ^ 
0; ///3



wire Ieeba56b21b21de0a3e58a479e445d91b;
assign Ieeba56b21b21de0a3e58a479e445d91b = 
        y_nr_enc[42] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p191 = 
Ieeba56b21b21de0a3e58a479e445d91b ^ 
0; ///3



wire Ifcc90797b4315701c136c4412f3f73f9;
assign Ifcc90797b4315701c136c4412f3f73f9 = 
        y_nr_enc[7] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p192 = 
Ifcc90797b4315701c136c4412f3f73f9 ^ 
0; ///3



wire Idc50751db38b20a4c10007bd9865490c;
assign Idc50751db38b20a4c10007bd9865490c = 
        y_nr_enc[4] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p193 = 
Idc50751db38b20a4c10007bd9865490c ^ 
0; ///3



wire I638ab1171b5e44484f0d2fff3fdb341c;
assign I638ab1171b5e44484f0d2fff3fdb341c = 
        y_nr_enc[5] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p194 = 
I638ab1171b5e44484f0d2fff3fdb341c ^ 
0; ///3



wire I5ec13d81e5e97dabed31d7fdde0ea208;
assign I5ec13d81e5e97dabed31d7fdde0ea208 = 
        y_nr_enc[6] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p195 = 
I5ec13d81e5e97dabed31d7fdde0ea208 ^ 
0; ///3



wire I79526ec250471ae5a81fab270e4d0ca3;
assign I79526ec250471ae5a81fab270e4d0ca3 = 
        y_nr_enc[3] ^ 
        y_nr_enc[28] ^ 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p196 = 
I79526ec250471ae5a81fab270e4d0ca3 ^ 
0; ///3



wire Iad9a6dc642b78393d4c6280fbb4dc8e6;
assign Iad9a6dc642b78393d4c6280fbb4dc8e6 = 
        y_nr_enc[0] ^ 
        y_nr_enc[29] ^ 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p197 = 
Iad9a6dc642b78393d4c6280fbb4dc8e6 ^ 
0; ///3



wire I641b2ccb0c26416d32a01168d530779e;
assign I641b2ccb0c26416d32a01168d530779e = 
        y_nr_enc[1] ^ 
        y_nr_enc[30] ^ 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p198 = 
I641b2ccb0c26416d32a01168d530779e ^ 
0; ///3



wire I4a11d7b58150d41429bb67f79e7c9db6;
assign I4a11d7b58150d41429bb67f79e7c9db6 = 
        y_nr_enc[2] ^ 
        y_nr_enc[31] ^ 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p199 = 
I4a11d7b58150d41429bb67f79e7c9db6 ^ 
0; ///3



wire I8adbebd85e789eeb0cac394c9e0a8e40;
assign I8adbebd85e789eeb0cac394c9e0a8e40 = 
        y_nr_enc[8] ^ 
        y_nr_enc[43] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p200 = 
I8adbebd85e789eeb0cac394c9e0a8e40 ^ 
0; ///3



wire I8eb469c3d856a33f1e16e6805abe19c9;
assign I8eb469c3d856a33f1e16e6805abe19c9 = 
        y_nr_enc[9] ^ 
        y_nr_enc[40] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p201 = 
I8eb469c3d856a33f1e16e6805abe19c9 ^ 
0; ///3



wire I5087bded2ded6668f1b2f9358a630698;
assign I5087bded2ded6668f1b2f9358a630698 = 
        y_nr_enc[10] ^ 
        y_nr_enc[41] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p202 = 
I5087bded2ded6668f1b2f9358a630698 ^ 
0; ///3



wire I3142c3d0ebdb884727dd18e17e71fde9;
assign I3142c3d0ebdb884727dd18e17e71fde9 = 
        y_nr_enc[11] ^ 
        y_nr_enc[42] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p203 = 
I3142c3d0ebdb884727dd18e17e71fde9 ^ 
0; ///3



wire I3f109fecebd9633b72dd5b58451f5969;
assign I3f109fecebd9633b72dd5b58451f5969 = 
        y_nr_enc[5] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p204 = 
I3f109fecebd9633b72dd5b58451f5969 ^ 
0; ///3



wire I311e0804831415fc0a4f108f6d5d9945;
assign I311e0804831415fc0a4f108f6d5d9945 = 
        y_nr_enc[6] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p205 = 
I311e0804831415fc0a4f108f6d5d9945 ^ 
0; ///3



wire Ic28767fb71b682f873988cfe9485c7d6;
assign Ic28767fb71b682f873988cfe9485c7d6 = 
        y_nr_enc[7] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p206 = 
Ic28767fb71b682f873988cfe9485c7d6 ^ 
0; ///3



wire I01b0a5d63b2b0cc2a17be22f9b7d2cc5;
assign I01b0a5d63b2b0cc2a17be22f9b7d2cc5 = 
        y_nr_enc[4] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p207 = 
I01b0a5d63b2b0cc2a17be22f9b7d2cc5 ^ 
0; ///3



