 reg  ['h7:0] [$clog2('h7000+1)-1:0] I00c7f323bbe2c226738efd26b205128d ;
