 reg  ['h7fff:0] [$clog2('h7000+1)-1:0] I2442159d7608347d1912b360378cc98d4372944f49dd911ce914ea8de1d3caa1 ;
