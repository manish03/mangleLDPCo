//`include "GF2_LDPC_flogtanh_0x0000d_assign_inc.sv"
//always_comb begin
              Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00000] = 
          (!flogtanh_sel['h0000d]) ? 
                       I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00000] : //%
                       I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00001] ;
//end
//always_comb begin
              Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00001] = 
          (!flogtanh_sel['h0000d]) ? 
                       I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00002] : //%
                       I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00003] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00002] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00004] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00003] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00006] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00004] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00008] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00005] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000a] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00006] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000c] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00007] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0000e] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00008] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00010] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00009] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00012] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000a] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00014] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000b] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00016] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000c] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00018] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000d] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001a] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000e] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001c] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0000f] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0001e] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00010] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00020] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00011] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00022] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00012] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00024] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00013] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00026] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00014] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00028] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00015] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002a] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00016] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002c] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00017] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0002e] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00018] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00030] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h00019] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00032] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001a] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00034] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001b] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00036] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001c] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h00038] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001d] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003a] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001e] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003c] ;
//end
//always_comb begin // 
               Id7629d0b91e01521c86c4e2f042518a92cbeefb68f14a9e332526a1425568478['h0001f] =  I3906fe88c24736f0823c1771293c3ca8ae92021844f3dc040deee9504a7f24ef['h0003e] ;
//end
