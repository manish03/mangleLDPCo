 reg  ['hf:0] [$clog2('h7000+1)-1:0] Iaf491f5f8d1574e1cb610cbd3edeca68 ;
