//`include "GF2_LDPC_flogtanh_0x00008_assign_inc.sv"
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00000] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00000] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00001] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00001] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00002] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00003] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00002] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00004] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00005] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00003] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00006] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00007] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00004] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00008] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00009] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00005] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000a] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000b] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00006] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000c] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000d] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00007] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000e] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0000f] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00008] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00010] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00011] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00009] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00012] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00013] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000a] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00014] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00015] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000b] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00016] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00017] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000c] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00018] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00019] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000d] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001a] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001b] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000e] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001c] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001d] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000f] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001e] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0001f] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00010] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00020] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00021] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00011] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00022] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00023] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00012] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00024] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00025] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00013] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00026] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00027] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00014] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00028] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00029] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00015] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002a] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002b] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00016] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002c] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002d] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00017] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002e] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0002f] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00018] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00030] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00031] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00019] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00032] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00033] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001a] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00034] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00035] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001b] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00036] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00037] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001c] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00038] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00039] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001d] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003a] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003b] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003c] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001f] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003e] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0003f] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00020] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00040] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00021] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00042] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00022] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00044] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00023] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00046] ;
//end
//always_comb begin
              Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00024] = 
          (!flogtanh_sel['h00008]) ? 
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00048] : //%
                       Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00049] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00025] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00026] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00027] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0004e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00028] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00050] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00029] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00052] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00054] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00056] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00058] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0005e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00030] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00060] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00031] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00062] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00032] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00064] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00033] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00066] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00034] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00068] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00035] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00036] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00037] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0006e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00038] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00070] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00039] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00072] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00074] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00076] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00078] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0007e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00040] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00080] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00041] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00082] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00042] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00084] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00043] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00086] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00044] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00088] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00045] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00046] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00047] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0008e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00048] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00090] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00049] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00092] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00094] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00096] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00098] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0009e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00050] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00051] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00052] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00053] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00054] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000a8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00055] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000aa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00056] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ac] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00057] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ae] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00058] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00059] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000b8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ba] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000bc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000be] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00060] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00061] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00062] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00063] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00064] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000c8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00065] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ca] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00066] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000cc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00067] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ce] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00068] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00069] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000d8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000da] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000dc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000de] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00070] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00071] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00072] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00073] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00074] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000e8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00075] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ea] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00076] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ec] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00077] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000ee] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00078] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00079] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000f8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000fa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000fc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h000fe] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00080] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00100] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00081] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00102] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00082] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00104] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00083] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00106] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00084] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00108] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00085] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00086] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00087] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0010e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00088] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00110] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00089] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00112] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00114] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00116] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00118] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0011e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00090] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00120] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00091] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00122] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00092] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00124] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00093] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00126] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00094] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00128] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00095] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00096] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00097] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0012e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00098] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00130] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00099] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00132] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00134] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00136] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00138] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0013e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00140] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00142] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00144] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00146] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00148] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0014e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00150] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00152] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000aa] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00154] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ab] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00156] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ac] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00158] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ad] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ae] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000af] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0015e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00160] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00162] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00164] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00166] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00168] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0016e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00170] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00172] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ba] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00174] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000bb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00176] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000bc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00178] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000bd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000be] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000bf] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0017e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00180] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00182] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00184] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00186] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00188] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0018e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00190] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00192] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ca] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00194] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000cb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00196] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000cc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00198] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000cd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ce] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000cf] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0019e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001a8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001aa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ac] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ae] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000da] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000db] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000dc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001b8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000dd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ba] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000de] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001bc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000df] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001be] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001c8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ca] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001cc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ce] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ea] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000eb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ec] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001d8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ed] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001da] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ee] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001dc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ef] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001de] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001e8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ea] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ec] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001ee] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000fa] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000fb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000fc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001f8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000fd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001fa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000fe] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001fc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ff] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h001fe] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00100] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00200] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00101] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00202] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00102] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00204] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00103] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00206] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00104] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00208] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00105] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00106] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00107] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0020e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00108] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00210] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00109] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00212] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00214] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00216] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00218] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0021e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00110] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00220] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00111] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00222] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00112] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00224] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00113] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00226] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00114] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00228] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00115] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00116] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00117] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0022e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00118] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00230] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00119] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00232] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00234] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00236] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00238] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0023e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00120] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00240] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00121] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00242] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00122] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00244] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00123] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00246] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00124] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00248] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00125] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00126] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00127] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0024e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00128] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00250] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00129] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00252] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00254] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00256] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00258] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0025e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00130] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00260] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00131] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00262] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00132] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00264] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00133] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00266] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00134] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00268] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00135] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00136] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00137] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0026e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00138] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00270] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00139] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00272] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00274] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00276] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00278] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0027e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00140] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00280] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00141] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00282] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00142] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00284] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00143] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00286] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00144] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00288] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00145] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00146] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00147] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0028e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00148] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00290] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00149] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00292] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00294] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00296] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00298] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0029e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00150] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00151] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00152] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00153] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00154] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002a8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00155] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002aa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00156] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ac] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00157] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ae] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00158] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00159] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002b8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ba] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002bc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002be] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00160] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00161] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00162] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00163] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00164] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002c8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00165] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ca] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00166] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002cc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00167] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ce] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00168] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00169] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002d8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002da] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002dc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002de] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00170] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00171] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00172] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00173] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00174] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002e8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00175] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ea] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00176] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ec] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00177] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002ee] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00178] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00179] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002f8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002fa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002fc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h002fe] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00180] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00300] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00181] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00302] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00182] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00304] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00183] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00306] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00184] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00308] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00185] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00186] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00187] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0030e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00188] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00310] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00189] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00312] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00314] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00316] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00318] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0031e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00190] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00320] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00191] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00322] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00192] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00324] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00193] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00326] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00194] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00328] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00195] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00196] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00197] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0032e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00198] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00330] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00199] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00332] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00334] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00336] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00338] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0033e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00340] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00342] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00344] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00346] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00348] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0034e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00350] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00352] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001aa] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00354] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ab] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00356] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ac] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00358] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ad] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ae] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001af] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0035e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00360] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00362] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00364] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00366] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00368] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0036e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00370] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00372] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ba] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00374] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001bb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00376] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001bc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00378] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001bd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001be] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001bf] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0037e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00380] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00382] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00384] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00386] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00388] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0038e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00390] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00392] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ca] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00394] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001cb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00396] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001cc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00398] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001cd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ce] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001cf] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0039e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003a8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003aa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ac] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ae] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001da] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001db] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001dc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003b8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001dd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ba] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001de] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003bc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001df] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003be] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003c8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ca] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003cc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ce] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ea] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001eb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ec] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003d8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ed] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003da] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ee] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003dc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ef] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003de] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003e8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ea] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ec] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003ee] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001fa] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001fb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001fc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003f8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001fd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003fa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001fe] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003fc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ff] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h003fe] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00200] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00400] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00201] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00402] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00202] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00404] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00203] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00406] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00204] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00408] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00205] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00206] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00207] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0040e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00208] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00410] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00209] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00412] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00414] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00416] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00418] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0041e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00210] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00420] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00211] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00422] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00212] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00424] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00213] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00426] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00214] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00428] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00215] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00216] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00217] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0042e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00218] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00430] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00219] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00432] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00434] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00436] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00438] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0043e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00220] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00440] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00221] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00442] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00222] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00444] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00223] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00446] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00224] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00448] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00225] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00226] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00227] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0044e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00228] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00450] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00229] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00452] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00454] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00456] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00458] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0045e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00230] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00460] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00231] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00462] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00232] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00464] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00233] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00466] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00234] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00468] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00235] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00236] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00237] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0046e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00238] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00470] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00239] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00472] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00474] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00476] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00478] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0047e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00240] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00480] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00241] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00482] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00242] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00484] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00243] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00486] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00244] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00488] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00245] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00246] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00247] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0048e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00248] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00490] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00249] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00492] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00494] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00496] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00498] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0049e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00250] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00251] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00252] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00253] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00254] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004a8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00255] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004aa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00256] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ac] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00257] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ae] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00258] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00259] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004b8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ba] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004bc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004be] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00260] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00261] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00262] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00263] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00264] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004c8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00265] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ca] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00266] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004cc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00267] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ce] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00268] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00269] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004d8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004da] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004dc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004de] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00270] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00271] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00272] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00273] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00274] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004e8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00275] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ea] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00276] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ec] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00277] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004ee] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00278] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00279] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004f8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004fa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004fc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h004fe] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00280] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00500] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00281] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00502] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00282] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00504] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00283] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00506] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00284] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00508] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00285] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00286] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00287] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0050e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00288] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00510] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00289] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00512] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00514] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00516] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00518] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0051e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00290] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00520] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00291] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00522] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00292] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00524] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00293] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00526] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00294] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00528] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00295] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00296] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00297] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0052e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00298] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00530] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00299] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00532] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00534] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00536] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00538] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0053e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00540] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00542] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00544] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00546] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00548] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0054e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00550] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00552] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002aa] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00554] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ab] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00556] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ac] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00558] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ad] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ae] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002af] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0055e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00560] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00562] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00564] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00566] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00568] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0056e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00570] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00572] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ba] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00574] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002bb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00576] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002bc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00578] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002bd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002be] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002bf] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0057e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00580] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00582] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00584] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00586] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00588] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0058e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00590] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00592] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ca] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00594] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002cb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00596] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002cc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00598] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002cd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ce] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002cf] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0059e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005a8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005aa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ac] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ae] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002da] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002db] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002dc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005b8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002dd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ba] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002de] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005bc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002df] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005be] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005c8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ca] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005cc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ce] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ea] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002eb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ec] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005d8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ed] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005da] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ee] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005dc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ef] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005de] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005e8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ea] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ec] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005ee] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002fa] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002fb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002fc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005f8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002fd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005fa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002fe] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005fc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ff] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h005fe] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00300] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00600] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00301] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00602] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00302] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00604] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00303] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00606] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00304] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00608] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00305] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00306] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00307] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0060e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00308] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00610] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00309] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00612] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00614] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00616] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00618] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0061e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00310] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00620] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00311] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00622] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00312] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00624] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00313] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00626] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00314] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00628] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00315] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00316] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00317] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0062e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00318] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00630] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00319] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00632] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00634] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00636] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00638] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0063e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00320] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00640] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00321] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00642] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00322] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00644] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00323] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00646] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00324] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00648] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00325] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00326] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00327] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0064e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00328] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00650] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00329] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00652] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00654] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00656] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00658] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0065e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00330] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00660] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00331] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00662] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00332] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00664] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00333] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00666] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00334] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00668] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00335] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00336] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00337] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0066e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00338] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00670] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00339] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00672] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00674] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00676] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00678] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0067e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00340] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00680] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00341] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00682] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00342] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00684] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00343] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00686] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00344] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00688] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00345] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00346] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00347] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0068e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00348] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00690] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00349] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00692] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00694] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00696] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00698] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0069e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00350] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00351] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00352] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00353] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00354] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006a8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00355] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006aa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00356] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ac] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00357] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ae] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00358] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00359] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006b8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ba] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006bc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006be] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00360] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00361] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00362] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00363] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00364] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006c8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00365] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ca] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00366] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006cc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00367] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ce] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00368] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00369] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006d8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006da] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006dc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006de] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00370] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00371] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00372] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00373] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00374] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006e8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00375] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ea] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00376] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ec] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00377] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006ee] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00378] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00379] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006f8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006fa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006fc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h006fe] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00380] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00700] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00381] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00702] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00382] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00704] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00383] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00706] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00384] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00708] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00385] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00386] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00387] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0070e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00388] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00710] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00389] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00712] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00714] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00716] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00718] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0071e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00390] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00720] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00391] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00722] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00392] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00724] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00393] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00726] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00394] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00728] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00395] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00396] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00397] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0072e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00398] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00730] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00399] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00732] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039a] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00734] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039b] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00736] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039c] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00738] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039d] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039e] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039f] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0073e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00740] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00742] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00744] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00746] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00748] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0074e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00750] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00752] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003aa] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00754] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ab] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00756] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ac] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00758] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ad] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ae] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003af] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0075e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00760] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00762] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00764] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00766] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00768] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0076e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00770] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00772] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ba] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00774] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003bb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00776] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003bc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00778] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003bd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003be] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003bf] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0077e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00780] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00782] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00784] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00786] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00788] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0078e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00790] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00792] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ca] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00794] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003cb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00796] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003cc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h00798] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003cd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079a] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ce] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079c] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003cf] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h0079e] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007a8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007aa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ac] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ae] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003da] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003db] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003dc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007b8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003dd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ba] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003de] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007bc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003df] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007be] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007c8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ca] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007cc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ce] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ea] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003eb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ec] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007d8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ed] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007da] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ee] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007dc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ef] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007de] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f0] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f1] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f2] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f3] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f4] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007e8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f5] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ea] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f6] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ec] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f7] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007ee] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f8] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f0] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f9] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f2] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003fa] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f4] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003fb] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f6] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003fc] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007f8] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003fd] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007fa] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003fe] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007fc] ;
//end
//always_comb begin // 
               Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ff] =  Id31f95377162c3f3bbc6cc895cc8ec54c7d906654125ec25295e3e5ac86f8756['h007fe] ;
//end
