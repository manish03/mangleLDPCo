              Ic4683a9b9f7e9b353f08f15f15d0cf43 = 
          (!flogtanh_sel[8]) ? 
                       If04be38ec93a9a9feffc2f86ea41a93e: 
                       I1732286809e19edc6b76b52139553c35;
               Ieec3fac0fc7bb3625400a15f74b1a15e =  0;
