              I51db5b688feb51ec24e6127d4c3dfdae = 
          (!flogtanh_sel[3]) ? 
                       I12635a66e3fe4dd930e858a0a7580cea: 
                       I71130fa5b933e0e26dbab66f37fb8925;
              Ibc891c78cf9dbf2365d9c88acc400657 = 
          (!flogtanh_sel[3]) ? 
                       I9371a6ffdba2a5bd6c4ac3fb38010117: 
                       I4001f1ca6d56d63aca19160a999b23de;
              I690dfdbfc7e73591927914aeb8cb121a = 
          (!flogtanh_sel[3]) ? 
                       Icf4458bcd36b49edb3c99d94980b2fcf: 
                       Ia336a15ef64f48975747202ff0586f96;
              I531efe3d41d7bc16091c3c247cebaaf0 = 
          (!flogtanh_sel[3]) ? 
                       I0ab4d4499b838b988c31c5d2162b0aa2: 
                       I8cc0695ebf79a9943050729478d73c9c;
              Icf7b3d66021580efed4e68c38d44ac48 = 
          (!flogtanh_sel[3]) ? 
                       I1207b10797bccdad5ee7e32abbfc9531: 
                       Ie37f7a4132d9db8e6589e4818da8f71e;
              I93d13a86c9d185bf2c3cf5c34eeeb016 = 
          (!flogtanh_sel[3]) ? 
                       Ief67dacff61c30f4f07a8b9426499320: 
                       I64c9510573d0b631cd08f41a30b4bf94;
              I3ded617611b49004853f17e60013d498 = 
          (!flogtanh_sel[3]) ? 
                       I496d08bbbe57943dde0a060794dd44f2: 
                       I6ea770088be3718bb9cbbf4015d7a698;
              Ia2414bf52998b14337d78da6aeaec255 = 
          (!flogtanh_sel[3]) ? 
                       I96e8e53f5e2fe546281cb33632075218: 
                       Iad67f635fc879ccccb83e4e8090e851f;
              Ieac60a94c2a709b738af1f3465a59240 = 
          (!flogtanh_sel[3]) ? 
                       Ic4eeb8715a3ab8d9da059d43c2f73e31: 
                       I06d19f878da9b67396ff63c2b0ac8a1e;
              I88349c865dbc4ddba373b69215a50400 = 
          (!flogtanh_sel[3]) ? 
                       Ied5797945822a58d6850b3d5472b6657: 
                       I79706d7caf960d3eee136724e1474c14;
              I72adcb5f4bd99318abd40c3b63287f93 = 
          (!flogtanh_sel[3]) ? 
                       Ic43fc3a05372e660dd974dd41d61966d: 
                       Id05004336c93a8f315406a56d1ea9401;
              I6cda0f5db099dbb900cd3d0a8f6dc245 = 
          (!flogtanh_sel[3]) ? 
                       I4257f21c0512ab632f6d8e3e49b6bc86: 
                       I38e64d8c0bfe85f483b46ad9d510bbf1;
              I4b7867a55677b1a9264c6d1c3eac25e4 = 
          (!flogtanh_sel[3]) ? 
                       If9f0572284b7c7b6fe299fb8f45c57d5: 
                       I248384903432b0ea141bdb0ba98bd3a3;
              I09a6bc8c6f42aa92f4b08511d5cd98b8 = 
          (!flogtanh_sel[3]) ? 
                       I81f42775b2a3e4badcc3910838808691: 
                       Iec5241a1c42d080412dff5e9494851e9;
              Ia64c991ab9c3fc3488a835de4fdb60b1 = 
          (!flogtanh_sel[3]) ? 
                       I1f10ad5fe2f55ebdb372cc672d8dd978: 
                       I1ca0505131c6887eaf1e7e80473e3add;
              I94cfcd3eeef047bb244a722337080b4d = 
          (!flogtanh_sel[3]) ? 
                       Ib49ad95d66dc9b1f5b9b225aa8124010: 
                       I1d942dd2be55359b99052dc72e795590;
               Ibebed3263875106ae630c0656211ee39 =  Id414b502a923f77f986b3c2f223798c4 ;
              I0439fd68942b4d70cdad2d56ee4b954c = 
          (!flogtanh_sel[3]) ? 
                       I1178b66ba1832d0acdf2683631bcebcc: 
                       I361d0be38e55d517342ea4b081c0fc23;
               If4c337b9bbfc2530377ac6db8f13014c =  I11ea42222da256fa229e3f7f74a29fd1 ;
               I9b705704a3308d69156c7343fa4eb777 =  I7714bd5031cea3a279cf989b22b30579 ;
               I5849744db9fdcad905885f296a170c02 =  Ic1ffa3d6c9037998cdf86b17c269216b ;
               I7cdf69d491d37935cef6eca36eb3fe81 =  I7780a0f25847a4e699619e564751c9a2 ;
              Idde15d5b821d09d8a406e09d1e4bda88 = 
          (!flogtanh_sel[3]) ? 
                       I64e434f7354d5b36a40f23792bed6616: 
                       Iae66d17c285d26bc13a560a3c46768ca;
               I944a0b47e85dab69de22e950ba042e2a =  0;
