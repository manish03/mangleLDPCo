              I48b438f1cbf654dacb5ca6bd28e924d6 = 
          (!flogtanh_sel[6]) ? 
                       I0ebde8b0a0a9c3a82d4f39df14847380: 
                       I2ae51e715df3b82f8423e1ff250759f8;
              I5e1d2582c82a255ad5580f16c60761e1 = 
          (!flogtanh_sel[6]) ? 
                       I07f0737fd7f5850a2cdb598766659236: 
                       Ie16c5883507cd5b149f7a43cd008f5ef;
              I32198fda41835969465ac7244753c104 = 
          (!flogtanh_sel[6]) ? 
                       I3c21bd722bd9c579d4bc131cce931bcf: 
                       I2c5fbe64fd51b745d0db44e5464155b0;
               I059f3ca58475484c4ed68b5ab609dbdf =  0;
