 parameter flogtanh_WDTH =  20 ;
 reg  [flogtanh_WDTH -1 :0] flogtanh_sel ;
 reg  ['h7ffff:0] [$clog2('h7000+1)-1:0] Ica91d9bac0dd49c3d4a33cbeec278026d5f4b3f1e4fdf2d3d75f4d666e11a0b2 ;
