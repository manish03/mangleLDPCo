//`include "GF2_LDPC_fgallag_0x00007_assign_inc.sv"
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00000] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00000] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00001] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00001] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00002] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00003] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00002] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00004] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00005] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00003] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00006] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00007] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00004] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00008] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00009] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00005] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000a] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000b] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00006] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000c] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000d] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00007] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000e] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0000f] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00008] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00010] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00011] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00009] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00012] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00013] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000a] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00014] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00015] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000b] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00016] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00017] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000c] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00018] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00019] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000d] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001a] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001b] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000e] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001c] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001d] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0000f] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001e] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0001f] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00010] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00020] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00021] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00011] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00022] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00023] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00012] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00024] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00025] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00013] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00026] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00027] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00014] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00028] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00029] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00015] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002a] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002b] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00016] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002c] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002d] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00017] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002e] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0002f] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00018] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00030] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00031] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00019] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00032] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00033] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001a] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00034] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00035] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001b] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00036] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00037] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001c] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00038] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00039] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001d] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003a] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003b] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001e] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003c] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003d] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0001f] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003e] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0003f] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00020] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00040] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00041] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00021] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00042] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00043] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00022] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00044] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00045] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00023] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00046] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00047] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00024] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00048] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00049] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00025] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004a] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004b] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00026] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004c] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004d] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00027] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004e] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0004f] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00028] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00050] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00051] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00029] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00052] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00053] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002a] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00054] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00055] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002b] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00056] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00057] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002c] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00058] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00059] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002d] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005a] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005b] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002e] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005c] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005d] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0002f] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005e] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0005f] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00030] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00060] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00061] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00031] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00062] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00063] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00032] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00064] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00065] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00033] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00066] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00067] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00034] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00068] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00069] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00035] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006a] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00036] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006c] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006d] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00037] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0006e] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00038] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00070] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00071] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00039] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00072] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00074] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003b] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00076] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00077] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00078] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007c] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0003f] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007e] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0007f] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00040] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00080] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00041] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00082] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00042] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00084] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00043] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00086] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00044] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00088] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00045] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00046] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00047] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0008e] ;
//end
//always_comb begin
              I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00048] = 
          (!fgallag_sel['h00007]) ? 
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00090] : //%
                       I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00091] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00049] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00092] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00094] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00096] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00098] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0004f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0009e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00050] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00051] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00052] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00053] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00054] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00055] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00056] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00057] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00058] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00059] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0005f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00060] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00061] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00062] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00063] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00064] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00065] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00066] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00067] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00068] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00069] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0006f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00070] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00071] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00072] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00073] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00074] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00075] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00076] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00077] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00078] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00079] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0007f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h000fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00080] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00100] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00081] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00102] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00082] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00104] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00083] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00106] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00084] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00108] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00085] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00086] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00087] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0010e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00088] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00110] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00089] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00112] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00114] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00116] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00118] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0008f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0011e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00090] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00120] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00091] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00122] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00092] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00124] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00093] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00126] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00094] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00128] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00095] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00096] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00097] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0012e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00098] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00130] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00099] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00132] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00134] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00136] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00138] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0009f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0013e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00140] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00142] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00144] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00146] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00148] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0014e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00150] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000a9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00152] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000aa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00154] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ab] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00156] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ac] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00158] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ad] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ae] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000af] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0015e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00160] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00162] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00164] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00166] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00168] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0016e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00170] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000b9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00172] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ba] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00174] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000bb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00176] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000bc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00178] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000bd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000be] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000bf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0017e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00180] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00182] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00184] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00186] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00188] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0018e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00190] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000c9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00192] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ca] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00194] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000cb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00196] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000cc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00198] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000cd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ce] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000cf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0019e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000d9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000da] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000db] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000dc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000dd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000de] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000df] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000e9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ea] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000eb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ec] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ed] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ee] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ef] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000f9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000fa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000fb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000fc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000fd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000fe] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h000ff] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h001fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00100] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00200] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00101] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00202] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00102] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00204] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00103] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00206] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00104] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00208] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00105] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00106] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00107] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0020e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00108] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00210] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00109] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00212] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00214] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00216] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00218] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0010f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0021e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00110] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00220] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00111] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00222] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00112] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00224] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00113] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00226] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00114] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00228] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00115] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00116] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00117] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0022e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00118] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00230] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00119] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00232] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00234] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00236] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00238] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0011f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0023e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00120] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00240] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00121] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00242] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00122] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00244] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00123] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00246] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00124] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00248] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00125] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00126] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00127] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0024e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00128] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00250] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00129] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00252] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00254] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00256] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00258] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0012f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0025e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00130] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00260] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00131] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00262] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00132] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00264] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00133] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00266] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00134] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00268] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00135] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00136] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00137] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0026e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00138] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00270] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00139] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00272] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00274] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00276] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00278] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0013f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0027e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00140] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00280] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00141] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00282] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00142] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00284] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00143] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00286] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00144] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00288] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00145] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00146] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00147] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0028e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00148] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00290] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00149] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00292] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00294] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00296] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00298] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0014f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0029e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00150] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00151] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00152] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00153] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00154] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00155] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00156] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00157] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00158] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00159] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0015f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00160] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00161] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00162] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00163] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00164] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00165] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00166] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00167] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00168] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00169] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0016f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00170] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00171] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00172] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00173] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00174] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00175] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00176] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00177] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00178] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00179] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0017f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h002fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00180] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00300] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00181] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00302] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00182] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00304] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00183] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00306] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00184] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00308] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00185] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00186] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00187] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0030e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00188] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00310] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00189] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00312] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00314] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00316] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00318] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0018f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0031e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00190] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00320] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00191] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00322] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00192] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00324] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00193] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00326] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00194] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00328] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00195] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00196] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00197] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0032e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00198] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00330] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00199] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00332] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00334] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00336] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00338] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0019f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0033e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00340] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00342] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00344] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00346] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00348] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0034e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00350] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001a9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00352] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001aa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00354] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ab] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00356] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ac] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00358] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ad] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ae] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001af] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0035e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00360] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00362] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00364] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00366] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00368] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0036e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00370] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001b9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00372] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ba] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00374] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001bb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00376] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001bc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00378] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001bd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001be] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001bf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0037e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00380] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00382] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00384] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00386] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00388] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0038e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00390] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001c9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00392] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ca] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00394] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001cb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00396] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001cc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00398] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001cd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ce] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001cf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0039e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001d9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001da] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001db] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001dc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001dd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001de] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001df] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001e9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ea] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001eb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ec] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ed] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ee] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ef] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001f9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001fa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001fb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001fc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001fd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001fe] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h001ff] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h003fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00200] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00400] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00201] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00402] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00202] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00404] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00203] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00406] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00204] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00408] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00205] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00206] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00207] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0040e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00208] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00410] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00209] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00412] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00414] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00416] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00418] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0020f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0041e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00210] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00420] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00211] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00422] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00212] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00424] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00213] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00426] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00214] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00428] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00215] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00216] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00217] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0042e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00218] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00430] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00219] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00432] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00434] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00436] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00438] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0021f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0043e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00220] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00440] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00221] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00442] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00222] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00444] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00223] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00446] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00224] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00448] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00225] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00226] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00227] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0044e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00228] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00450] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00229] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00452] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00454] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00456] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00458] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0022f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0045e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00230] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00460] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00231] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00462] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00232] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00464] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00233] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00466] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00234] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00468] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00235] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00236] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00237] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0046e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00238] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00470] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00239] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00472] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00474] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00476] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00478] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0023f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0047e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00240] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00480] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00241] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00482] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00242] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00484] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00243] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00486] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00244] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00488] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00245] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00246] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00247] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0048e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00248] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00490] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00249] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00492] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00494] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00496] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00498] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0024f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0049e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00250] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00251] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00252] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00253] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00254] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00255] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00256] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00257] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00258] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00259] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0025f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00260] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00261] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00262] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00263] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00264] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00265] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00266] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00267] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00268] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00269] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0026f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00270] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00271] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00272] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00273] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00274] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00275] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00276] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00277] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00278] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00279] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0027f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h004fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00280] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00500] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00281] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00502] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00282] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00504] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00283] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00506] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00284] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00508] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00285] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00286] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00287] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0050e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00288] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00510] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00289] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00512] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00514] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00516] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00518] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0028f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0051e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00290] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00520] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00291] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00522] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00292] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00524] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00293] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00526] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00294] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00528] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00295] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00296] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00297] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0052e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00298] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00530] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00299] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00532] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00534] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00536] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00538] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0029f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0053e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00540] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00542] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00544] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00546] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00548] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0054e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00550] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002a9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00552] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002aa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00554] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ab] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00556] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ac] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00558] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ad] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ae] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002af] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0055e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00560] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00562] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00564] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00566] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00568] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0056e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00570] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002b9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00572] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ba] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00574] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002bb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00576] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002bc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00578] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002bd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002be] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002bf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0057e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00580] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00582] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00584] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00586] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00588] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0058e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00590] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002c9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00592] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ca] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00594] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002cb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00596] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002cc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00598] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002cd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ce] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002cf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0059e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002d9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002da] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002db] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002dc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002dd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002de] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002df] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002e9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ea] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002eb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ec] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ed] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ee] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ef] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002f9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002fa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002fb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002fc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002fd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002fe] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h002ff] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h005fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00300] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00600] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00301] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00602] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00302] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00604] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00303] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00606] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00304] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00608] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00305] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00306] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00307] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0060e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00308] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00610] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00309] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00612] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00614] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00616] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00618] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0030f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0061e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00310] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00620] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00311] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00622] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00312] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00624] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00313] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00626] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00314] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00628] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00315] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00316] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00317] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0062e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00318] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00630] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00319] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00632] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00634] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00636] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00638] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0031f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0063e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00320] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00640] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00321] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00642] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00322] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00644] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00323] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00646] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00324] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00648] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00325] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00326] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00327] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0064e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00328] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00650] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00329] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00652] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00654] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00656] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00658] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0032f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0065e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00330] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00660] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00331] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00662] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00332] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00664] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00333] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00666] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00334] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00668] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00335] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00336] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00337] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0066e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00338] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00670] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00339] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00672] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00674] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00676] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00678] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0033f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0067e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00340] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00680] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00341] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00682] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00342] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00684] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00343] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00686] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00344] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00688] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00345] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00346] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00347] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0068e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00348] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00690] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00349] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00692] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00694] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00696] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00698] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0034f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0069e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00350] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00351] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00352] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00353] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00354] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00355] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00356] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00357] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00358] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00359] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0035f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00360] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00361] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00362] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00363] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00364] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00365] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00366] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00367] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00368] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00369] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0036f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00370] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00371] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00372] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00373] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00374] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00375] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00376] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00377] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00378] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00379] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0037f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h006fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00380] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00700] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00381] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00702] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00382] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00704] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00383] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00706] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00384] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00708] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00385] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00386] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00387] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0070e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00388] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00710] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00389] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00712] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00714] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00716] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00718] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0038f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0071e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00390] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00720] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00391] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00722] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00392] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00724] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00393] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00726] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00394] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00728] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00395] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00396] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00397] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0072e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00398] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00730] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00399] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00732] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00734] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00736] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00738] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0039f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0073e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00740] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00742] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00744] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00746] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00748] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0074e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00750] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003a9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00752] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003aa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00754] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ab] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00756] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ac] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00758] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ad] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ae] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003af] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0075e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00760] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00762] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00764] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00766] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00768] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0076e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00770] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003b9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00772] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ba] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00774] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003bb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00776] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003bc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00778] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003bd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003be] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003bf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0077e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00780] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00782] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00784] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00786] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00788] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0078e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00790] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003c9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00792] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ca] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00794] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003cb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00796] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003cc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00798] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003cd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ce] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003cf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0079e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003d9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003da] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003db] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003dc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003dd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003de] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003df] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003e9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ea] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003eb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ec] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ed] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ee] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ef] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003f9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003fa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003fb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003fc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003fd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003fe] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h003ff] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h007fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00400] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00800] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00401] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00802] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00402] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00804] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00403] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00806] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00404] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00808] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00405] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00406] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00407] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0080e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00408] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00810] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00409] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00812] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00814] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00816] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00818] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0040f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0081e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00410] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00820] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00411] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00822] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00412] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00824] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00413] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00826] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00414] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00828] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00415] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00416] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00417] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0082e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00418] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00830] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00419] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00832] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00834] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00836] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00838] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0041f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0083e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00420] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00840] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00421] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00842] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00422] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00844] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00423] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00846] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00424] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00848] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00425] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00426] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00427] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0084e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00428] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00850] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00429] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00852] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00854] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00856] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00858] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0042f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0085e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00430] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00860] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00431] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00862] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00432] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00864] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00433] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00866] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00434] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00868] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00435] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00436] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00437] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0086e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00438] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00870] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00439] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00872] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00874] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00876] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00878] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0043f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0087e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00440] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00880] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00441] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00882] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00442] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00884] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00443] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00886] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00444] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00888] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00445] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00446] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00447] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0088e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00448] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00890] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00449] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00892] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00894] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00896] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00898] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0044f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0089e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00450] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00451] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00452] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00453] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00454] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00455] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00456] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00457] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00458] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00459] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0045f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00460] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00461] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00462] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00463] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00464] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00465] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00466] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00467] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00468] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00469] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0046f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00470] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00471] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00472] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00473] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00474] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00475] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00476] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00477] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00478] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00479] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0047f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h008fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00480] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00900] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00481] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00902] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00482] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00904] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00483] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00906] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00484] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00908] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00485] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00486] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00487] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0090e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00488] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00910] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00489] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00912] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00914] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00916] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00918] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0048f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0091e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00490] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00920] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00491] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00922] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00492] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00924] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00493] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00926] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00494] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00928] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00495] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00496] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00497] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0092e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00498] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00930] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00499] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00932] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00934] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00936] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00938] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0049f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0093e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00940] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00942] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00944] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00946] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00948] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0094e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00950] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004a9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00952] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004aa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00954] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ab] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00956] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ac] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00958] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ad] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ae] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004af] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0095e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00960] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00962] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00964] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00966] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00968] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0096e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00970] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004b9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00972] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ba] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00974] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004bb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00976] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004bc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00978] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004bd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004be] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004bf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0097e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00980] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00982] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00984] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00986] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00988] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0098e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00990] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004c9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00992] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ca] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00994] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004cb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00996] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004cc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00998] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004cd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ce] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004cf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h0099e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009a8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009aa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004d9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004da] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004db] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004dc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009b8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004dd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004de] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009bc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004df] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009be] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009c8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009cc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004e9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ea] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004eb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ec] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009d8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ed] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009da] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ee] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009dc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ef] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009de] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009e8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009ee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004f9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004fa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004fb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004fc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009f8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004fd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009fa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004fe] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009fc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h004ff] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h009fe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00500] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a00] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00501] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a02] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00502] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a04] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00503] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a06] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00504] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a08] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00505] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00506] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00507] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a0e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00508] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a10] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00509] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a12] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a14] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a16] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a18] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0050f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a1e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00510] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a20] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00511] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a22] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00512] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a24] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00513] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a26] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00514] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a28] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00515] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00516] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00517] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a2e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00518] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a30] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00519] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a32] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a34] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a36] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a38] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0051f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a3e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00520] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a40] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00521] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a42] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00522] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a44] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00523] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a46] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00524] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a48] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00525] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00526] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00527] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a4e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00528] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a50] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00529] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a52] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a54] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a56] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a58] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0052f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a5e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00530] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a60] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00531] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a62] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00532] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a64] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00533] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a66] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00534] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a68] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00535] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00536] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00537] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a6e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00538] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a70] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00539] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a72] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a74] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a76] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a78] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0053f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a7e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00540] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a80] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00541] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a82] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00542] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a84] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00543] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a86] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00544] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a88] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00545] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00546] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00547] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a8e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00548] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a90] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00549] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a92] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a94] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a96] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a98] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0054f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00a9e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00550] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00551] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00552] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00553] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00554] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aa8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00555] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aaa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00556] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00557] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00558] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00559] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ab8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00abc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0055f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00abe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00560] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00561] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00562] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00563] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00564] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ac8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00565] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00566] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00acc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00567] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ace] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00568] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00569] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ad8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ada] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00adc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0056f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ade] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00570] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00571] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00572] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00573] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00574] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ae8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00575] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00576] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00577] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00aee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00578] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00579] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00af8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00afa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00afc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0057f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00afe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00580] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b00] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00581] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b02] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00582] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b04] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00583] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b06] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00584] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b08] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00585] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00586] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00587] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b0e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00588] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b10] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00589] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b12] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b14] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b16] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b18] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0058f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b1e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00590] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b20] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00591] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b22] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00592] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b24] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00593] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b26] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00594] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b28] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00595] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00596] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00597] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b2e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00598] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b30] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00599] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b32] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b34] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b36] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b38] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0059f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b3e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b40] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b42] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b44] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b46] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b48] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b4e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b50] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005a9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b52] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005aa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b54] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ab] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b56] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ac] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b58] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ad] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ae] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005af] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b5e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b60] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b62] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b64] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b66] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b68] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b6e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b70] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005b9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b72] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ba] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b74] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005bb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b76] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005bc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b78] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005bd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005be] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005bf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b7e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b80] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b82] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b84] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b86] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b88] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b8e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b90] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005c9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b92] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ca] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b94] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005cb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b96] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005cc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b98] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005cd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ce] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005cf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00b9e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ba8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00baa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005d9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005da] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005db] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005dc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bb8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005dd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005de] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bbc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005df] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bbe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bc8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bcc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005e9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ea] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005eb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ec] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bd8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ed] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bda] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ee] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bdc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ef] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bde] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00be8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005f9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005fa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005fb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005fc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bf8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005fd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bfa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005fe] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bfc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h005ff] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00bfe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00600] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c00] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00601] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c02] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00602] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c04] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00603] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c06] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00604] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c08] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00605] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00606] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00607] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c0e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00608] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c10] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00609] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c12] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c14] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c16] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c18] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0060f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c1e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00610] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c20] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00611] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c22] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00612] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c24] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00613] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c26] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00614] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c28] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00615] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00616] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00617] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c2e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00618] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c30] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00619] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c32] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c34] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c36] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c38] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0061f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c3e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00620] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c40] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00621] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c42] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00622] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c44] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00623] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c46] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00624] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c48] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00625] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00626] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00627] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c4e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00628] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c50] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00629] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c52] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c54] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c56] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c58] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0062f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c5e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00630] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c60] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00631] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c62] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00632] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c64] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00633] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c66] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00634] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c68] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00635] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00636] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00637] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c6e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00638] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c70] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00639] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c72] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c74] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c76] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c78] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0063f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c7e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00640] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c80] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00641] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c82] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00642] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c84] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00643] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c86] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00644] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c88] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00645] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00646] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00647] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c8e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00648] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c90] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00649] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c92] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c94] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c96] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c98] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0064f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00c9e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00650] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00651] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00652] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00653] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00654] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ca8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00655] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00caa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00656] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00657] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00658] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00659] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cb8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cbc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0065f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cbe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00660] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00661] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00662] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00663] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00664] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cc8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00665] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00666] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ccc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00667] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00668] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00669] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cd8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cda] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cdc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0066f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cde] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00670] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00671] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00672] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00673] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00674] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ce8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00675] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00676] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00677] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00678] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00679] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cf8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cfa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cfc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0067f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00cfe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00680] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d00] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00681] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d02] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00682] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d04] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00683] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d06] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00684] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d08] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00685] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00686] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00687] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d0e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00688] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d10] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00689] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d12] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d14] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d16] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d18] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0068f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d1e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00690] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d20] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00691] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d22] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00692] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d24] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00693] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d26] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00694] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d28] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00695] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00696] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00697] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d2e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00698] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d30] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00699] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d32] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d34] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d36] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d38] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0069f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d3e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d40] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d42] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d44] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d46] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d48] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d4e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d50] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006a9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d52] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006aa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d54] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ab] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d56] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ac] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d58] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ad] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ae] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006af] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d5e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d60] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d62] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d64] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d66] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d68] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d6e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d70] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006b9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d72] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ba] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d74] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006bb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d76] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006bc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d78] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006bd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006be] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006bf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d7e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d80] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d82] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d84] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d86] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d88] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d8e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d90] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006c9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d92] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ca] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d94] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006cb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d96] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006cc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d98] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006cd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ce] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006cf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00d9e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00da8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00daa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006d9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006da] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006db] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006dc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00db8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006dd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006de] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dbc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006df] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dbe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dc8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dcc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006e9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ea] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006eb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ec] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dd8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ed] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dda] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ee] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ddc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ef] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dde] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00de8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006f9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006fa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006fb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006fc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00df8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006fd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dfa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006fe] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dfc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h006ff] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00dfe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00700] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e00] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00701] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e02] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00702] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e04] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00703] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e06] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00704] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e08] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00705] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00706] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00707] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e0e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00708] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e10] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00709] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e12] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e14] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e16] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e18] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0070f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e1e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00710] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e20] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00711] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e22] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00712] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e24] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00713] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e26] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00714] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e28] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00715] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00716] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00717] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e2e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00718] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e30] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00719] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e32] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e34] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e36] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e38] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0071f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e3e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00720] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e40] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00721] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e42] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00722] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e44] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00723] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e46] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00724] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e48] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00725] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00726] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00727] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e4e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00728] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e50] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00729] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e52] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e54] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e56] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e58] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0072f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e5e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00730] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e60] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00731] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e62] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00732] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e64] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00733] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e66] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00734] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e68] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00735] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00736] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00737] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e6e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00738] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e70] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00739] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e72] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e74] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e76] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e78] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0073f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e7e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00740] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e80] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00741] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e82] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00742] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e84] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00743] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e86] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00744] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e88] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00745] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00746] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00747] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e8e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00748] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e90] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00749] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e92] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e94] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e96] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e98] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0074f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00e9e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00750] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00751] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00752] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00753] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00754] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ea8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00755] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eaa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00756] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00757] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00758] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00759] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eb8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ebc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0075f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ebe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00760] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00761] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00762] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00763] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00764] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ec8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00765] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00766] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ecc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00767] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ece] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00768] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00769] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ed8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eda] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00edc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0076f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ede] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00770] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00771] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00772] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00773] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00774] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ee8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00775] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00776] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00777] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00eee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00778] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00779] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ef8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00efa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00efc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0077f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00efe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00780] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f00] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00781] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f02] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00782] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f04] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00783] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f06] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00784] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f08] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00785] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00786] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00787] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f0e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00788] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f10] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00789] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f12] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f14] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f16] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f18] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0078f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f1e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00790] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f20] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00791] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f22] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00792] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f24] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00793] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f26] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00794] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f28] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00795] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00796] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00797] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f2e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00798] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f30] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h00799] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f32] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079a] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f34] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079b] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f36] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079c] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f38] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079d] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079e] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h0079f] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f3e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f40] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f42] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f44] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f46] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f48] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f4e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f50] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007a9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f52] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007aa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f54] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ab] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f56] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ac] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f58] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ad] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ae] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007af] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f5e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f60] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f62] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f64] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f66] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f68] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f6e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f70] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007b9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f72] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ba] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f74] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007bb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f76] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007bc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f78] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007bd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007be] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007bf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f7e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f80] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f82] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f84] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f86] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f88] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f8e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f90] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007c9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f92] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ca] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f94] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007cb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f96] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007cc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f98] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007cd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9a] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ce] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9c] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007cf] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00f9e] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fa8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00faa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fac] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fae] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007d9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007da] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007db] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007dc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fb8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007dd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fba] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007de] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fbc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007df] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fbe] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fc8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fca] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fcc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fce] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007e9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ea] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007eb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ec] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fd8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ed] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fda] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ee] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fdc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ef] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fde] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f0] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f1] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f2] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f3] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f4] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fe8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f5] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fea] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f6] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fec] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f7] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00fee] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f8] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff0] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007f9] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff2] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007fa] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff4] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007fb] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff6] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007fc] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ff8] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007fd] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ffa] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007fe] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ffc] ;
//end
//always_comb begin // 
               I0c57c163ee894fdcb1c6da15086e6ec08b964c5000d5982e713702657833a2ed['h007ff] =  I20046edea7caab9a45d6a51441f123cad6d25f9c59fe5a903c9a070b3e16dbb9['h00ffe] ;
//end
