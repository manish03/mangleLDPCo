              I67f92596363d7abd702880c8dd319453 = 
          (!fgallag_sel[3]) ? 
                       I2e449260cbba5283dbe9d183eaa3006b: 
                       Ie43af039b1e5b11fe91210b644a1a31e;
              I58dc37dd8f90b2815ebae43223ff2268 = 
          (!fgallag_sel[3]) ? 
                       Iebddca10e7f7c3688d5011f147ffcd4a: 
                       I93b9a635a3e05192ad53b6e264275aa9;
              Ic5c9b0ef750a107380673521819d09e5 = 
          (!fgallag_sel[3]) ? 
                       Ie3012c652b244e53fc44455982b5eefa: 
                       Ie287c2f7d9779d50be27d3d5a9de6a33;
              I6d82716e87b1ac554c6ff5e4169afe0b = 
          (!fgallag_sel[3]) ? 
                       Ia9327a6a37a1de7dbf3839eafb5d941e: 
                       I47705f99ef5cb6172811f4046484597c;
              I64fc488e4651b1cde21e870d2528613c = 
          (!fgallag_sel[3]) ? 
                       Ie1c96dc77190cd04130a400e869a5abd: 
                       Iafcc3b17af5dbd70300172c2e2742206;
              Ice7c81f4524a3e2a6ec0b6e7d76fe9b6 = 
          (!fgallag_sel[3]) ? 
                       I47731679e4d0f87f9d19934c25f2bdcb: 
                       I9608c445e266884a86508e3ea3a53853;
              If1b3191923af5d433e5d97adf41bd97f = 
          (!fgallag_sel[3]) ? 
                       I0fb3749641e7b5675524cd796ef4127c: 
                       Id5b6b690dc055c374a44fb1ecfd54198;
              If2cca0ade959a72defe62fb3eef484e4 = 
          (!fgallag_sel[3]) ? 
                       I6ae44809304b38046cc0afb4317a3f43: 
                       I3ef49ef515a84b68f7bff1fbc0f05be7;
              Ida8b253166cc056c54916e14755c6aa6 = 
          (!fgallag_sel[3]) ? 
                       I62939bc5509a6ca4278bedb7be3f4534: 
                       Ieaaab9e41c6a940e06ce877c3e6faebc;
              If1ac872a756deb15fa93f38bc63700c3 = 
          (!fgallag_sel[3]) ? 
                       Iadf3bdeaff4bc193443ef22aef0ad7b7: 
                       Ic65a2079483506c24674715cc402a81b;
              Ia8342322e4b86c946f8a133fc284bd4f = 
          (!fgallag_sel[3]) ? 
                       Ia7641d441a79bfea63ba407052928bc5: 
                       I299c542d09419d0998b59bf1f184a78a;
              I316bb23418efb56e676cc0a58e8f0e19 = 
          (!fgallag_sel[3]) ? 
                       I8aa5ad4f2f437be64a88554e6dfc3c6b: 
                       Iaf0980a21e4ee5e842a5b6db664264f6;
              Ib659aa347010e749163015d2457712b7 = 
          (!fgallag_sel[3]) ? 
                       I80df82d24c9507274353efb085b46fda: 
                       I1db5a382bb7c2317716c3137fd10d07c;
              Id87f3e882b2fb1c5af8b4134c83dff16 = 
          (!fgallag_sel[3]) ? 
                       Icb748243d2a5f8cc86c44566e1732232: 
                       I90a0c6bd80d2357d7b865f61a18ae13b;
              I0eda2f2f507535ab778d59c7ce193447 = 
          (!fgallag_sel[3]) ? 
                       I16af13e02ee36dbcdeab785596175a3c: 
                       Id0e47470fba20bc467a05d0dd09bf560;
              If36a4176048d1fec4e9646d016b5a33b = 
          (!fgallag_sel[3]) ? 
                       I944adac3cc097911cde333e806fa004c: 
                       I3292848fc7b015c9900b92b702ba7be9;
               Id3ffa72548f440a0e3a90db8b5ff1c39 =  Ie09561c5bcd6107bd956faddcdddc89c ;
              Ic36450e12061ae80189b6f16d1cab329 = 
          (!fgallag_sel[3]) ? 
                       I4274fedf54de3b2a34285844c7a34519: 
                       I4fae388e04252b896bd4e9c527a8c0af;
               Iec0fe238288bd4b3f41ddec347477271 =  Ia3c4f467d029cc1ea1c0993e0d314978 ;
               Iff515d269a292258ff61605083324963 =  I38fe32f3f6de6ff9c3fcb5644ac3eb66 ;
               I13b529dfc9f09f5208d2df5a91e4eabe =  If54d6a9d910097237f3e20059257bf57 ;
               If5686d7de8ada834d078111dd1557853 =  I16027735edf5e40e34bd73920ae40fb7 ;
              I4393932a40ca1c79aa95d652d504c5f6 = 
          (!fgallag_sel[3]) ? 
                       Ib819132b8eb007862e294bb775a7cd3b: 
                       Icfd0596c8f143d0536c06d827bc30018;
               Ia4abb71881c5f95a1a30badf83a0a567 =  0;
