reg [fgallag_WDTH -1:0] fgallag0x00005_0, fgallag0x00005_0_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_1, fgallag0x00005_1_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_2, fgallag0x00005_2_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_3, fgallag0x00005_3_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_4, fgallag0x00005_4_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_5, fgallag0x00005_5_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_6, fgallag0x00005_6_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_7, fgallag0x00005_7_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_8, fgallag0x00005_8_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_9, fgallag0x00005_9_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_10, fgallag0x00005_10_q;
reg [fgallag_WDTH -1:0] fgallag0x00005_11, fgallag0x00005_11_q;
reg start_d_fgallag0x00005_q ;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 fgallag0x00005_0_q <= 'h0;
 fgallag0x00005_1_q <= 'h0;
 fgallag0x00005_2_q <= 'h0;
 fgallag0x00005_3_q <= 'h0;
 fgallag0x00005_4_q <= 'h0;
 fgallag0x00005_5_q <= 'h0;
 fgallag0x00005_6_q <= 'h0;
 fgallag0x00005_7_q <= 'h0;
 fgallag0x00005_8_q <= 'h0;
 fgallag0x00005_9_q <= 'h0;
 fgallag0x00005_10_q <= 'h0;
 fgallag0x00005_11_q <= 'h0;
 start_d_fgallag0x00005_q <= 'h0;
end
else
begin
 fgallag0x00005_0_q <=  fgallag0x00005_0;
 fgallag0x00005_1_q <=  fgallag0x00005_1;
 fgallag0x00005_2_q <=  fgallag0x00005_2;
 fgallag0x00005_3_q <=  fgallag0x00005_3;
 fgallag0x00005_4_q <=  fgallag0x00005_4;
 fgallag0x00005_5_q <=  fgallag0x00005_5;
 fgallag0x00005_6_q <=  fgallag0x00005_6;
 fgallag0x00005_7_q <=  fgallag0x00005_7;
 fgallag0x00005_8_q <=  fgallag0x00005_8;
 fgallag0x00005_9_q <=  fgallag0x00005_9;
 fgallag0x00005_10_q <=  fgallag0x00005_10;
 fgallag0x00005_11_q <=  fgallag0x00005_11;
 start_d_fgallag0x00005_q <=  start_d_fgallag0x00004_q;
end
