//`include "GF2_LDPC_flogtanh_0x00010_assign_inc.sv"
//always_comb begin
              Ib43d6a3ec9a1741fe7beed3535eddb34['h00000] = 
          (!flogtanh_sel['h00010]) ? 
                       I00c7f323bbe2c226738efd26b205128d['h00000] : //%
                       I00c7f323bbe2c226738efd26b205128d['h00001] ;
//end
//always_comb begin // 
               Ib43d6a3ec9a1741fe7beed3535eddb34['h00001] =  I00c7f323bbe2c226738efd26b205128d['h00002] ;
//end
//always_comb begin // 
               Ib43d6a3ec9a1741fe7beed3535eddb34['h00002] =  I00c7f323bbe2c226738efd26b205128d['h00004] ;
//end
//always_comb begin // 
               Ib43d6a3ec9a1741fe7beed3535eddb34['h00003] =  I00c7f323bbe2c226738efd26b205128d['h00006] ;
//end
