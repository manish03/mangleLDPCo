 reg  ['h3:0] [$clog2('h7000+1)-1:0] Ib43d6a3ec9a1741fe7beed3535eddb34 ;
