 reg  ['h3:0] [$clog2('h7000+1)-1:0] I23c1c03fb2d7ef8b2dc0921ddaf652a0 ;
