 reg  ['h1ffff:0] [$clog2('h7000+1)-1:0] I76b88463fe716cf89c65112ab35e2f39 ;
