//`include "GF2_LDPC_flogtanh_0x0000c_assign_inc.sv"
//always_comb begin
              Ie4acdb20b1de9050267f708a13a337e0['h00000] = 
          (!flogtanh_sel['h0000c]) ? 
                       I111cd97f7c5c13e18b528ffe1d1a871f['h00000] : //%
                       I111cd97f7c5c13e18b528ffe1d1a871f['h00001] ;
//end
//always_comb begin
              Ie4acdb20b1de9050267f708a13a337e0['h00001] = 
          (!flogtanh_sel['h0000c]) ? 
                       I111cd97f7c5c13e18b528ffe1d1a871f['h00002] : //%
                       I111cd97f7c5c13e18b528ffe1d1a871f['h00003] ;
//end
//always_comb begin
              Ie4acdb20b1de9050267f708a13a337e0['h00002] = 
          (!flogtanh_sel['h0000c]) ? 
                       I111cd97f7c5c13e18b528ffe1d1a871f['h00004] : //%
                       I111cd97f7c5c13e18b528ffe1d1a871f['h00005] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00003] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00006] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00004] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00008] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00005] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0000a] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00006] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0000c] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00007] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0000e] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00008] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00010] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00009] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00012] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0000a] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00014] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0000b] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00016] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0000c] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00018] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0000d] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0001a] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0000e] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0001c] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0000f] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0001e] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00010] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00020] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00011] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00022] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00012] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00024] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00013] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00026] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00014] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00028] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00015] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0002a] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00016] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0002c] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00017] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0002e] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00018] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00030] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00019] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00032] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0001a] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00034] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0001b] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00036] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0001c] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00038] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0001d] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0003a] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0001e] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0003c] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0001f] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0003e] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00020] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00040] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00021] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00042] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00022] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00044] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00023] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00046] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00024] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00048] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00025] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0004a] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00026] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0004c] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00027] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0004e] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00028] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00050] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00029] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00052] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0002a] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00054] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0002b] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00056] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0002c] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00058] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0002d] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0005a] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0002e] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0005c] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0002f] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0005e] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00030] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00060] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00031] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00062] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00032] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00064] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00033] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00066] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00034] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00068] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00035] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0006a] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00036] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0006c] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00037] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0006e] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00038] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00070] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h00039] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00072] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0003a] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00074] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0003b] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00076] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0003c] =  I111cd97f7c5c13e18b528ffe1d1a871f['h00078] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0003d] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0007a] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0003e] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0007c] ;
//end
//always_comb begin // 
               Ie4acdb20b1de9050267f708a13a337e0['h0003f] =  I111cd97f7c5c13e18b528ffe1d1a871f['h0007e] ;
//end
