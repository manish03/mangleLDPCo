//`include "GF2_LDPC_fgallag_0x0000d_assign_inc.sv"
//always_comb begin
              Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00000] = 
          (!fgallag_sel['h0000d]) ? 
                       Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00000] : //%
                       Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00001] ;
//end
//always_comb begin
              Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00001] = 
          (!fgallag_sel['h0000d]) ? 
                       Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00002] : //%
                       Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00003] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00002] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00004] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00003] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00006] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00004] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00008] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00005] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0000a] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00006] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0000c] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00007] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0000e] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00008] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00010] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00009] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00012] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000a] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00014] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000b] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00016] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000c] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00018] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000d] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0001a] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000e] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0001c] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0000f] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0001e] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00010] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00020] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00011] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00022] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00012] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00024] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00013] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00026] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00014] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00028] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00015] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0002a] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00016] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0002c] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00017] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0002e] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00018] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00030] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h00019] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00032] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001a] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00034] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001b] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00036] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001c] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h00038] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001d] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0003a] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001e] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0003c] ;
//end
//always_comb begin // 
               Id18c9b63a7692cd190147c4a515a897a2801605bcfeba142ecaeb4a102f6187d['h0001f] =  Ibadc2e1716f3631bf6927ab6aa76689d577d209baf59b74521b39c268f0c78b6['h0003e] ;
//end
