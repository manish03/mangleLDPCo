 reg  ['h3fff:0] [$clog2('h7000+1)-1:0] Ib8f6031ee1aaf052d1ff517a16f81423d544c8722ad77f26af27e52332a8b50b ;
