 reg  ['hff:0] [$clog2('h7000+1)-1:0] I45c1a80dd59b47025bbf3f233589964b ;
