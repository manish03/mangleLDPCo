//`include "GF2_LDPC_flogtanh_0x00009_assign_inc.sv"
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00000] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00000] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00001] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00001] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00002] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00003] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00002] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00004] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00005] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00003] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00006] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00007] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00004] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00008] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00009] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00005] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000a] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000b] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00006] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000c] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000d] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00007] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000e] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0000f] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00008] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00010] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00011] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00009] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00012] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00013] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000a] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00014] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00015] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000b] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00016] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00017] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000c] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00018] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00019] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000d] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001a] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001b] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000e] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001c] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001d] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000f] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001e] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0001f] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00010] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00020] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00011] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00022] ;
//end
//always_comb begin
              I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00012] = 
          (!flogtanh_sel['h00009]) ? 
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00024] : //%
                       Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00025] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00013] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00026] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00014] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00028] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00015] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00016] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00017] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0002e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00018] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00030] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00019] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00032] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00034] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00036] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00038] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0003e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00020] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00040] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00021] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00042] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00022] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00044] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00023] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00046] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00024] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00048] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00025] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00026] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00027] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0004e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00028] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00050] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00029] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00052] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00054] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00056] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00058] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0005e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00030] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00060] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00031] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00062] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00032] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00064] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00033] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00066] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00034] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00068] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00035] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00036] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00037] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0006e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00038] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00070] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00039] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00072] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00074] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00076] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00078] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0007e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00040] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00080] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00041] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00082] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00042] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00084] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00043] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00086] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00044] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00088] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00045] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00046] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00047] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0008e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00048] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00090] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00049] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00092] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00094] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00096] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00098] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0009e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00050] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00051] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00052] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00053] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00054] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000a8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00055] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000aa] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00056] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ac] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00057] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ae] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00058] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00059] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000b8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ba] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000bc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000be] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00060] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00061] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00062] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00063] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00064] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000c8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00065] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ca] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00066] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000cc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00067] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ce] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00068] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00069] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000d8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000da] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000dc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000de] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00070] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00071] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00072] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00073] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00074] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000e8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00075] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ea] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00076] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ec] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00077] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000ee] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00078] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00079] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000f8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000fa] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000fc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h000fe] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00080] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00100] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00081] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00102] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00082] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00104] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00083] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00106] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00084] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00108] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00085] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00086] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00087] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0010e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00088] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00110] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00089] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00112] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00114] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00116] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00118] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0011e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00090] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00120] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00091] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00122] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00092] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00124] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00093] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00126] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00094] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00128] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00095] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00096] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00097] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0012e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00098] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00130] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00099] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00132] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00134] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00136] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00138] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0013e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00140] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00142] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00144] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00146] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00148] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0014e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00150] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00152] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000aa] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00154] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ab] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00156] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ac] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00158] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ad] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ae] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000af] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0015e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00160] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00162] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00164] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00166] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00168] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0016e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00170] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00172] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ba] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00174] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000bb] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00176] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000bc] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00178] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000bd] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000be] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000bf] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0017e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00180] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00182] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00184] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00186] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00188] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0018e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00190] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00192] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ca] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00194] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000cb] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00196] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000cc] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00198] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000cd] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ce] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000cf] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0019e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001a8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001aa] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ac] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ae] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000da] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000db] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000dc] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001b8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000dd] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ba] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000de] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001bc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000df] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001be] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001c8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ca] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001cc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ce] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ea] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000eb] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ec] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001d8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ed] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001da] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ee] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001dc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ef] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001de] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001e8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ea] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ec] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001ee] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000fa] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000fb] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000fc] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001f8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000fd] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001fa] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000fe] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001fc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ff] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h001fe] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00100] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00200] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00101] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00202] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00102] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00204] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00103] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00206] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00104] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00208] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00105] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00106] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00107] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0020e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00108] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00210] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00109] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00212] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00214] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00216] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00218] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0021e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00110] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00220] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00111] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00222] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00112] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00224] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00113] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00226] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00114] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00228] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00115] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00116] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00117] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0022e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00118] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00230] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00119] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00232] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00234] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00236] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00238] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0023e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00120] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00240] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00121] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00242] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00122] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00244] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00123] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00246] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00124] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00248] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00125] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00126] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00127] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0024e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00128] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00250] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00129] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00252] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00254] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00256] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00258] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0025e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00130] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00260] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00131] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00262] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00132] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00264] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00133] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00266] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00134] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00268] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00135] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00136] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00137] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0026e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00138] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00270] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00139] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00272] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00274] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00276] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00278] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0027e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00140] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00280] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00141] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00282] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00142] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00284] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00143] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00286] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00144] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00288] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00145] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00146] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00147] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0028e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00148] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00290] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00149] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00292] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00294] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00296] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00298] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0029e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00150] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00151] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00152] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00153] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00154] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002a8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00155] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002aa] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00156] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ac] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00157] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ae] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00158] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00159] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002b8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ba] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002bc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002be] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00160] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00161] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00162] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00163] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00164] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002c8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00165] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ca] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00166] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002cc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00167] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ce] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00168] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00169] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002d8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002da] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002dc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002de] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00170] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00171] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00172] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00173] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00174] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002e8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00175] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ea] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00176] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ec] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00177] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002ee] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00178] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00179] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002f8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002fa] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002fc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h002fe] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00180] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00300] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00181] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00302] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00182] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00304] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00183] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00306] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00184] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00308] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00185] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00186] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00187] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0030e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00188] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00310] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00189] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00312] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00314] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00316] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00318] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0031e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00190] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00320] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00191] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00322] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00192] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00324] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00193] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00326] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00194] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00328] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00195] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00196] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00197] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0032e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00198] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00330] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00199] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00332] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019a] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00334] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019b] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00336] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019c] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00338] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019d] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019e] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019f] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0033e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00340] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00342] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00344] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00346] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00348] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0034e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00350] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00352] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001aa] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00354] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ab] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00356] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ac] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00358] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ad] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ae] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001af] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0035e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00360] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00362] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00364] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00366] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00368] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0036e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00370] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00372] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ba] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00374] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001bb] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00376] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001bc] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00378] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001bd] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001be] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001bf] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0037e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00380] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00382] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00384] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00386] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00388] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0038e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00390] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00392] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ca] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00394] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001cb] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00396] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001cc] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h00398] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001cd] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039a] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ce] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039c] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001cf] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h0039e] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003a8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003aa] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ac] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ae] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001da] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001db] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001dc] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003b8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001dd] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ba] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001de] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003bc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001df] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003be] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003c8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ca] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003cc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ce] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ea] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001eb] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ec] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003d8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ed] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003da] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ee] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003dc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ef] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003de] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f0] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f1] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f2] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f3] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f4] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003e8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f5] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ea] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f6] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ec] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f7] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003ee] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f8] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f0] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f9] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f2] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001fa] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f4] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001fb] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f6] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001fc] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003f8] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001fd] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003fa] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001fe] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003fc] ;
//end
//always_comb begin // 
               I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ff] =  Ic1bf043b809d2d1ac03904940e7ca4b6dcd8582b75bb3593bbf904983c9b5441['h003fe] ;
//end
