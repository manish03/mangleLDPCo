 reg  ['h1fff:0] [$clog2('h7000+1)-1:0] If409768b648a33a7ed878a070d4f6251 ;
