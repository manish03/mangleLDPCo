reg [fgallag_WDTH -1:0] I0b93aca5ef7c84ffba0064eb4a53ec4f,  I53846946a877f30f72076ee6f633a0e5;
reg [fgallag_WDTH -1:0] Id37ee8cb85e5cd05bbe92dd90fd22777,  I5d219e3294f2763bc17209a55758ab54;
reg [fgallag_WDTH -1:0] I41450c30addcb3bb1d2c1c036dc26d2f,  I6273ee09aacad20f733530af1a987ff3;
reg [fgallag_WDTH -1:0] I078a7802a3340b0c207a002a4046a4e3,  Ie0f63a67c0a6ec07e7bcb943e7804f9a;
reg [fgallag_WDTH -1:0] I5a33c28f0bc44840136790663423bd48,  I7b83ef4e45fe20e023e08aa3e56bb21e;
reg [fgallag_WDTH -1:0] I777e21d17f74d2fe893977e1654e2c2d,  Ibc8f334cefc147e5c58e7542d26fbe2b;
reg [fgallag_WDTH -1:0] I0b457f5bce1ac08077d7c061655dd03f,  I662a566f576ee431bced6f852294713e;
reg [fgallag_WDTH -1:0] I8d508a837624b899a748b9152f4a787d,  I2a4bc966b71864a79f582727f122ab60;
reg [fgallag_WDTH -1:0] Ib226330c1225db758177402a9bcb4848,  I23d9f47edf51ff1c2a6275531a1f66be;
reg [fgallag_WDTH -1:0] Ic9d6b4cdd3bfef73660bcd8319a9a7be,  Id46ae2d16f43af3529d91eb4d6bd098e;
reg [fgallag_WDTH -1:0] I8e094e0c0b13b04dee8f4f70fdee87c4,  I51298122656d9b893c1dbb33a281f134;
reg [fgallag_WDTH -1:0] I5469abe94b035be8eb8713d061774eb5,  I22e0a22ed1768671dbe3caef8ac499cb;
reg [fgallag_WDTH -1:0] Ic6dd18ea6082a83222edb24cff9873da,  Ifb9327c663379f77471d460eced9c1b7;
reg [fgallag_WDTH -1:0] If46aa2c29de75a5a44a4d629204b0963,  Id6080749dda3cd29c1ce36ab39759709;
reg [fgallag_WDTH -1:0] I86f471de37f4d7f2599425d1f7ae60b9,  I532fd8f9065e524727e276a1a8408008;
reg [fgallag_WDTH -1:0] Id4063c01903ecbf60f39cc2a65c5b73e,  I1f0b23c673ff55115f55c80a970172fc;
reg [fgallag_WDTH -1:0] I1be4f732652b930e60cb6bf53fbb7132,  I9f99ad4587fb6907b3804c11125f738f;
reg [fgallag_WDTH -1:0] I64355c5e822a8d545c6fded925a984b6,  I719bd7e94d4289c6fd59bb91ee559980;
reg [fgallag_WDTH -1:0] I865085332575d46654188a23e78a5ab5,  I9103b57e3550cb68266ba8b102e50dfd;
reg [fgallag_WDTH -1:0] I5a3af3b67e01e19177daaa19b995b876,  I89fca1c1832813b84cafe145377d7b5e;
reg [fgallag_WDTH -1:0] Ic82f2a7d5019f0912c100d6336dfb3a8,  Ie17de6e388779502a143212813a50317;
reg [fgallag_WDTH -1:0] Icaa4f34ed9aaa9f1690a03ff7c374de4,  Ifcc046128364b8da7bc3d9ddab96a061;
reg [fgallag_WDTH -1:0] I7662e29bd142424284880f29b6d32038,  Iabe4b7a23f682ed62162dfde9e15d6cf;
reg [fgallag_WDTH -1:0] Ib9befe6fabe9ca87ddb96713b6c6e0d4,  I734eaef0b7d7f6ae5d668ac9b374ff51;
reg [fgallag_WDTH -1:0] I69bd49e2f242a3c2a32d182a32cf39f8,  I0e0e9fdfeb3e2115deb903b973217384;
reg [fgallag_WDTH -1:0] I820044a9516905bcd63a9e6d98ec961d,  Ibfd2fd7aa2426054706d0c4e4c0a7cba;
reg [fgallag_WDTH -1:0] I4b1cce4cb416fc1776b09254d2589bfe,  I0906247e3ba96971232bc42185c9a9b8;
reg [fgallag_WDTH -1:0] I9cae305381503e9d92a4a8240bb2aac0,  Ia3908fda391d7caf1b479d9655164c30;
reg [fgallag_WDTH -1:0] I5a1301cdc00c141cd57b0c4b90d7dd7a,  I820e95cdc583108195e8dd0e2d1f4b7f;
reg [fgallag_WDTH -1:0] I98abd404eafd5efdc2a990f2760fb0d9,  Ibdf5c2c57269da1b04748a59802c8e2a;
reg [fgallag_WDTH -1:0] I3e8a5169cec2e8120a2ba6b6dc0f5742,  Idd85c8c853438679d99bed4d0ba46af7;
reg [fgallag_WDTH -1:0] I8b50f6cf167c2ec62d739f294512c324,  I4d617d0b669b3ff1b08dcd4b7440af33;
reg [fgallag_WDTH -1:0] Ib0fffb83f9af51787fff93443dd10287,  I60d579b60b02f9fc14e98d7d0eb54c18;
reg [fgallag_WDTH -1:0] I3e4d4fb93b28d431849e2dd307f91197,  Ic1a37750fc3d7eb08ad649de157f45a9;
reg [fgallag_WDTH -1:0] I85b43efcd6de020aceb66ed5948fd901,  I0c13ec63e7208b35a1d4511e1da29fa3;
reg [fgallag_WDTH -1:0] Ibf4c9739576bfc4c8d79dcdbdb629a6d,  If10c9545a713996735934c5f15cf5365;
reg [fgallag_WDTH -1:0] Ib96063e5603755f2354a15d573374fe0,  Ic475963164a956dd24ede91e9d61003d;
reg [fgallag_WDTH -1:0] I5f07fe122c1bb26c6805a7f9d31218db,  I42001c4b6ab9fb03489ca25defb6c222;
reg [fgallag_WDTH -1:0] I0ed871a78ca4e2815ce45133571353a1,  Idcfb16adf2996c8cb51e402daafd1734;
reg [fgallag_WDTH -1:0] Ib0ba4dc6303dade812ab25816938899e,  I924108a2723afd07735574a6f4ebe671;
reg [fgallag_WDTH -1:0] Iea7ffe40a13deb5bfe2903c2965e4b63,  If9fd9ae380997e75ebed2ddd3f93e76f;
reg [fgallag_WDTH -1:0] Iad7d1d253ed65347182adf53486dc1de,  Ief876b7b2af1fbed4d3f457cdb46e0d9;
reg [fgallag_WDTH -1:0] Ie4cc734fa69e1b46577b5df885ba3592,  Id2bd196ca25e1a077fb2a9207f143c01;
reg [fgallag_WDTH -1:0] I75554ec87598151940cd118e6ee59741,  I926e2a038d48db29b5ce215cd6cf6a04;
reg [fgallag_WDTH -1:0] Ifec751297668f80d860a9d6cc176e5f8,  I4ba2cfd94590dee1723ce63afd0926ab;
reg [fgallag_WDTH -1:0] I8fcbbdfd901920672268b4d6ca269849,  I0d42326464ae4c3a55038e0343cebf5a;
reg [fgallag_WDTH -1:0] Id16656f72b76591b0bd03a3c2750684c,  If05fde321fd1456422550f5c3903b826;
reg [fgallag_WDTH -1:0] Iefa235bdb6e83afe1f793787d8dfca2f,  I41ec48a5a1d657a6266b8f845550d0c2;
reg [fgallag_WDTH -1:0] Id4fc19c089fa63c1b901fb64c9c0e064,  I76473b4885d423029324fe74ed13d6ed;
reg [fgallag_WDTH -1:0] Ib22f4bce6db16f279ad4085901174664,  I8ef2366947e3f1352f3874e4ac58d7b2;
reg [fgallag_WDTH -1:0] I432b06e788f0047c5e66cac253186eca,  I874c1e455f85e617a5032ec230fdfdc5;
reg [fgallag_WDTH -1:0] I51d270bbc6e26272e0d6998307c33272,  I16d6b6b19890a6bbdf15ddc27717aa30;
reg [fgallag_WDTH -1:0] I7f0c42c0c3c63ba11cdd3c26093bc3f5,  I6af6d04126eec9eb91e5653cc95c9ef3;
reg [fgallag_WDTH -1:0] Ibe2e871186cde032e6ce4de65c0fbf75,  If501a668f24fd62a69d0e3c253739c79;
reg [fgallag_WDTH -1:0] I9aaab4112c129c0563c8983c3cb372ba,  I9b70e215a2a1578811b40c669826d41a;
reg [fgallag_WDTH -1:0] I58b6cde8739d1e98ccbdd13b1a963c8f,  I26d82966efbe51e03edcd66a5a507ebb;
reg [fgallag_WDTH -1:0] I6d3d948976b4f578039a6dbaa8f08642,  I2e4afb94e4af76b4e3d859815bb338fb;
reg [fgallag_WDTH -1:0] I714b8ce615cf088e1ac52a7e22eb69df,  Ie19faf5d037b74974102c386a13f4946;
reg [fgallag_WDTH -1:0] I7672fb8749f7573c27144fffd1721ef7,  I2d56338af0755ae5c4ef71ddad3112b1;
reg [fgallag_WDTH -1:0] I5fa7ef4e8130409885342236b9f60fcd,  I99ab212db901b0e65eb33be27c46bd19;
reg [fgallag_WDTH -1:0] I2ab7e691bb0a2f89f9cdbfbad80d7120,  If8c09c14d78b1deaf76df6f4de910c64;
reg [fgallag_WDTH -1:0] Idc22eb4529d6e2f82fd6c23a113809da,  I1b0ccac0f5cc741403fd6e680899f96f;
reg [fgallag_WDTH -1:0] I449ee1a89494568e104c9e29f66d4262,  I38153cd88e8b2452977d7dc9b9f44a74;
reg [fgallag_WDTH -1:0] I5e8f226f92643e61ad527be4f148de00,  Ic32064fc62eb1cdcdf416a6fe78becfd;
reg [fgallag_WDTH -1:0] I56a2b51825ae20cd1d9b434aa976b4dd,  Ic10eb104fe38a176a51507e748406958;
reg [fgallag_WDTH -1:0] I580e0ae47b151812c4373cb1f268e4fe,  I979fd1b01c99b76a4ff2d0abfb0c2ae9;
reg [fgallag_WDTH -1:0] I69e6eeed488ce445421bf458f3d1baaf,  Ibe530a86c501fbc8dba64ed24806bdf4;
reg [fgallag_WDTH -1:0] Ie3781ac0023a6e8091d66990ee3983ff,  If03531315c68272f7de2b0e969770f48;
reg [fgallag_WDTH -1:0] Ia6a4c1e9dcb6ab1ad0114e2da7a396bc,  I20160f4e380b0920bcb30a0321b7bfa8;
reg [fgallag_WDTH -1:0] I91ed400a23a8aa771dbb930317b63466,  I2bbbe5d3a72af5f654976a7fde2d2d16;
reg [fgallag_WDTH -1:0] I15c7e1315b03dc87984424245b7e6dab,  I70f4396800d2cb065ad5fe655bacbfd0;
reg [fgallag_WDTH -1:0] I4ae2e6ccef3d457713203f83eb10d60d,  If27a0187d1188cf7a8aba100a90cb069;
reg [fgallag_WDTH -1:0] I08a273aa764a26045fd205007493d27a,  I8994866d080b1befe414fea347e7e74a;
reg [fgallag_WDTH -1:0] Ifae99596becf8c2c7b69fc3e508a362a,  Iab6971c846299eec0a5cc93ad10e569c;
reg [fgallag_WDTH -1:0] Ib080cdead060a391cb67c54d97c7fb0b,  I8730924fec54ffaa78a0ffea7e8386ba;
reg [fgallag_WDTH -1:0] Ie14db629163bf8c01b457b0df3bbb634,  I338fb9183219691c6b50e6a824fcb14c;
reg [fgallag_WDTH -1:0] Ib4c7a688661be990227b9902dcaa0721,  I1a3d82eaf2fc9235163c0a50765f4ef5;
reg [fgallag_WDTH -1:0] I4b33852fd89354d5eeaaf75dcb84e726,  I922539f8d9ffc119ed3a5c92a21f149e;
reg [fgallag_WDTH -1:0] I982d1672a39f86bf7da5bb7844bd57f9,  I3bc0f1eaad327d5990adb826e54c6d2f;
reg [fgallag_WDTH -1:0] I29949584d0bbd464970883cc5724f8a4,  I3009d4cc0371f83e6bec8fb38ae461bd;
reg [fgallag_WDTH -1:0] I03ec49385def83a3f577d847012976fc,  I2e0ae02d7a3cdfa36e8645cc7dd0bce6;
reg [fgallag_WDTH -1:0] I6bb12bbec43b6315c92ac22f43ef5a60,  If2c59f326f3658dee0fd3b048af14cb7;
reg [fgallag_WDTH -1:0] I5c49372712967408ed819ba89624dc98,  I04431bd4be4601d3cb700c0cd6d9fd24;
reg [fgallag_WDTH -1:0] I477fb86a2ad5f7ed4f225b0c85609bee,  I7a6fe8c804087a19e32e760f50e3edfa;
reg [fgallag_WDTH -1:0] I67099935c6636fc80d472f193753ba55,  I979817e250e46dcc05f8a6690c2380f9;
reg [fgallag_WDTH -1:0] Icf692082f362b6bb08f320e2b27853c7,  I3bbb836eee6b5e10fe55879f8620b888;
reg [fgallag_WDTH -1:0] Iae5385d0436fb1f5c949c0d1e8c3aa96,  I8bc5128382cbffa289caec56f9b4a3f3;
reg [fgallag_WDTH -1:0] I6951d4063e974375523406edae080570,  Iee4dafc9d42609fae74410897f29a78d;
reg [fgallag_WDTH -1:0] I54e637eae832d289eeba34eda853a657,  I4ea5b39ed827d8d4618bcfd9283dfa83;
reg [fgallag_WDTH -1:0] I89479946789730c4000d8166356cb964,  I19aa6440394778642eb50f3b94098ea3;
reg [fgallag_WDTH -1:0] Ide9c460b12322a14105bd0484d4b9135,  I0653a9ef861e5d8af22d120172c2dc03;
reg [fgallag_WDTH -1:0] Icb6633d32c69b880dea230dbae0896cd,  Ie0aafaeee1abf6d27a70535385ab88b5;
reg [fgallag_WDTH -1:0] Icc91b46df090bdc04306996433be6136,  I1583cdcd13120f953691a5a60ee72b11;
reg [fgallag_WDTH -1:0] I5ac7c7696f008ebbaf6019fa5ad57302,  I8080b45a37a3de79ccb338f353f19529;
reg [fgallag_WDTH -1:0] Iab7f04bf5075b64439bff52f4779ca67,  I9bd98a9d18ce7c07e85287f6b80bfd31;
reg [fgallag_WDTH -1:0] I9c3e9f415a26edb9fedf25288a8fa453,  Ife85d240c60084dce9b3d7cd87060727;
reg [fgallag_WDTH -1:0] If0e39a30beb041d9c6b3c168e965a1af,  I11f2e4eafc706b43c10a26edc8567052;
reg [fgallag_WDTH -1:0] Ibb59c086a89025918626f18799e73605,  Iad3a9febf269d9607eedf29912b04af9;
reg [fgallag_WDTH -1:0] Ic436ebe8aa48c3e6e935f6ce0b3f43d5,  I75705fa2cc0ac0577570501510e4e0fc;
reg [fgallag_WDTH -1:0] I05239dbfe2cd2ef57477ecb654880bf4,  I7674ab7538766e842366dd08ddbbcb28;
reg [fgallag_WDTH -1:0] I1765216a10c88b6081f34198e8a5d26f,  I8cefcac1f7fa2df45bb8a2f3d64f99c3;
reg [fgallag_WDTH -1:0] I37b9f75cb896a9e45a650b6dadd0b2ff,  I5fd378ba266fd930a839cad56e500ef4;
reg [fgallag_WDTH -1:0] Ib9eeab393231e41cca081394b036bde6,  I71a33ca1c7d18d5089d08a8476c8baf7;
reg [fgallag_WDTH -1:0] I499fb85792bd0c5a73022ac96ac27f13,  Ic85b012b9fa77becd419cac0f3692aed;
reg [fgallag_WDTH -1:0] I3da1d9759bbad87b216b2bc8afc19f8e,  I0ae9b4ca5ebb5f3d2e8b02884069e4e7;
reg [fgallag_WDTH -1:0] Ie220bafbf40ee68b7591948b607fcaa0,  Ief312304eec0415d1ab208ed6726dd12;
reg [fgallag_WDTH -1:0] I34b7451c43eee381ab7b3f1e2a816b99,  Icb9ebf1f5becaede273da59f466506ac;
reg [fgallag_WDTH -1:0] I5a3b2767a2c2b41984b6f2a7f05dfcbc,  I465b9607a8dad0f1c499318d04f42aea;
reg [fgallag_WDTH -1:0] I8ad73072ca340501c2b14404b9353b08,  I2523c109974807b3b1c0f4b34693e255;
reg [fgallag_WDTH -1:0] Id3987a88bcc92458973c9ee529f52a56,  Ib4e3121afd90b877b94c4c7cd29e9334;
reg [fgallag_WDTH -1:0] I49666607354671cb5d6ec9c3e6354f42,  Ibfb66b89c59008f3d4497ee16dad6712;
reg [fgallag_WDTH -1:0] I4da0ec3a6c662f7e76bd3f6c43b40722,  I2d042c4ef15b2f3bdebbc7cbd6c00a1f;
reg [fgallag_WDTH -1:0] I039f5eff8e87d37a9cf7d754a82df849,  I489d1b46970800e9684c68b439c15be1;
reg [fgallag_WDTH -1:0] Ia6fa92e40471f5741d59b8515c67c24b,  I835143e23243f3fd25cc1ab0ba5c123a;
reg [fgallag_WDTH -1:0] Ib4ce242cd8f88c4eb147129be5e6785c,  I028ef05ea84be3bc45c518f4f45653d2;
reg [fgallag_WDTH -1:0] Icc28fa9f2f20d09b439a9553b6e592fa,  Ia5a39eeda95dfdb2ab8b55ea9f8b62c5;
reg [fgallag_WDTH -1:0] I8b4b437c18f15ae386e0c12371151913,  If5a85945ad1f8d9bdc9213c5ae2c890f;
reg [fgallag_WDTH -1:0] I7c34ca74407090b532ec5f0f65e5dc74,  I6011a5fc7b168a28fc9a45f796629b59;
reg [fgallag_WDTH -1:0] I1f69904e43d7fb93f39873efcbbb558b,  Ie703b5f1eeedaaaddf56ded14b1765bc;
reg [fgallag_WDTH -1:0] Ie1f3985459b6de4b08d14263f5b1aa18,  I21f34fbc269f5424ea30334ff7ab54f5;
reg [fgallag_WDTH -1:0] I3640c422ee8389926afc8108564b593b,  I07b47fce56edeb30319038e3a093efd7;
reg [fgallag_WDTH -1:0] Ie11fa9bb26231d41be8646707525d022,  I24e7e5c391285f28c20f74820a05b552;
reg [fgallag_WDTH -1:0] Ibabb39952458fdb3127ed17f3909e043,  Iee1b23b99f7de56829706633297a0513;
reg [fgallag_WDTH -1:0] I8b1452ad1732c78b5397caddc0d43daa,  Ib4b61d3293900c38e8aa7df0a617b476;
reg [fgallag_WDTH -1:0] I5adc876cca35af9714a2cb9ca0eb3ae1,  Ifd5fcb1552fb372ae203fd0166d3df2c;
reg [fgallag_WDTH -1:0] Ia2848a15587c0e23eef1de69c2a238b1,  Ibb2fb63aef1d336dfa829cd5ab3675b7;
reg [fgallag_WDTH -1:0] Ic4119a74d5a813a98baede5515be91bc,  I1672371cf33b259cf87210cc49aa35c8;
reg [fgallag_WDTH -1:0] Id3b3231272ef7b602acb9b7dcd5033e8,  Ia34735ee7f7ca164c2ae71980060f56b;
reg [fgallag_WDTH -1:0] I05e604f9ffc573b44538d9d864dd4e92,  I2372d0a72998f0630e994aa3e1c20ff4;
reg [fgallag_WDTH -1:0] I116d21ad2753927dbf389f373bb1a344,  I8e363e0bd65cae9725cdd70e46778fee;
reg [fgallag_WDTH -1:0] I3805a70a8e257eeea2bdc179fba1d185,  Id6af962a16ff79ac6e9da3b4518b80b2;
reg [fgallag_WDTH -1:0] Ie2d31cc4673f92faf8545984e9b52031,  I7fc8c9245183d05370746c9b2fdabd0f;
reg [fgallag_WDTH -1:0] I5bbb1e57ed53613e06ba3fe1cc4fd266,  I693f2c9a5d4da90c3105876991c4f4ba;
reg [fgallag_WDTH -1:0] Ic4e117cdda2e62382412fb1dfb9c850d,  Id6c07cd1f9f428b0d971639939b9eb8e;
reg [fgallag_WDTH -1:0] Iab33d8521b7118693333cb5f624f3904,  Id6561e53aa8f9fd116159969afaa20ae;
reg [fgallag_WDTH -1:0] I4183bbdffed2418b9190d610ef9c85a5,  I8267af03225d6d1155142645ad7f53a8;
reg [fgallag_WDTH -1:0] Ibee805f0c9d18428759c5ce6c61f4dee,  I567872d8892064b62caeb3dcdc39e89c;
reg [fgallag_WDTH -1:0] Ic8255e62414174e60282be5b4d63c494,  I5072b405191b837596b5efe4ec159519;
reg [fgallag_WDTH -1:0] Ie76911ee442cfab80022b3a534438350,  Ia4e5d30bc160c1f72c8f39cdcd13e5a4;
reg [fgallag_WDTH -1:0] Ie9d09a2059dea91a80a00bdeb56940f2,  Ic46dd8ff5a79971f7c22f4be0f1f4b23;
reg [fgallag_WDTH -1:0] I86ecfe340941ed77c09fd4c69f5c272a,  Ifdd13523ba0ce3329e3aca49a0a36385;
reg [fgallag_WDTH -1:0] I511c8519304a31c10313838c1a053f85,  Ib449b5d80a7f5a1c5d0d3784d8f236b6;
reg [fgallag_WDTH -1:0] I8824abf0eb1a4d6b48a26abae23d0bff,  I134d223e71b68cc9c76379f1368fb0f1;
reg [fgallag_WDTH -1:0] I5d8953fa34cb14027d8375d02999f132,  Ifa82272c492ce1ed4b223c0cb2b135e1;
reg [fgallag_WDTH -1:0] I0d8e31fd51ec5b82c5206c307e0d53f7,  Ie501d0f392be1309df48c1616ace5a27;
reg [fgallag_WDTH -1:0] Ie1ea3318d114c790e9343e45555755ab,  I29468f8318cd5bebb5cea27e1ee57b7f;
reg [fgallag_WDTH -1:0] I495a91d95803df2b5cfca5053bf13a9b,  Ie3f06a529d5f22198b3b33d649b740e1;
reg [fgallag_WDTH -1:0] Ide9b85fb8d57bdfbf9b8de9c18e9c5cd,  I6740505fac3e83de4a6525ac9cf489d1;
reg [fgallag_WDTH -1:0] I9cd4f5d3b10c25759e7993f9292a7390,  I0456541b6e82ffeb05fc4052fafc41f7;
reg [fgallag_WDTH -1:0] I5ea9ea2fd34572dc6833ccf368e52ccb,  I6d5739cf589ed46b6f57075a3b2a974d;
reg [fgallag_WDTH -1:0] If3883c5646540cf78aee0589c3cd3022,  Iabe05603679da24a44565e756adc0881;
reg [fgallag_WDTH -1:0] I61df05bea32eda79ed88930bbc84a13f,  Icaed4c0a915898eea654ab6f93973ff3;
reg [fgallag_WDTH -1:0] I7f1a2ad313f7af4a0f9eb4311f35ac12,  I98805e117c2f4ba4a8f6c2755ebe1fee;
reg [fgallag_WDTH -1:0] I685601482e2bded73351f69f3f5c21b2,  I766076681dc49b817ec9302eae86d64b;
reg [fgallag_WDTH -1:0] I484b91ff2256c38308e18bc50afed4ef,  Ia82b6e01034a63c2a1a446029f58f1c6;
reg [fgallag_WDTH -1:0] Id86467d5f10985a00ab65a8b029a8c82,  I05de7fd67a0e226201b563fa6c50f362;
reg [fgallag_WDTH -1:0] I56110e27931a312345e239eaf42781a2,  I8df8f128712fe5445a97566f8f29ecd4;
reg [fgallag_WDTH -1:0] Iee57da8134718b73f0598a1884ecf424,  Iae9103582be213e81ea0a25e5d49004f;
reg [fgallag_WDTH -1:0] I7de0f163ab38efee6f9c2f362708f4a0,  Ibcab213dbb173403005b3d65f780fa2d;
reg [fgallag_WDTH -1:0] Id397e815fb86c38fbb509692ec4dab0b,  Ic59b57cadd4b8cbe63f996111e9211b1;
reg [fgallag_WDTH -1:0] I2c5e75d48e9ca1a198d70980900bdc41,  Ide1a993a1dfca37107fc81e985714d93;
reg [fgallag_WDTH -1:0] If728db81c67f83aab133c8ceaa3a5c7b,  I7004a1bc0ec2272163d33907d21616ea;
reg [fgallag_WDTH -1:0] I80d54bec914a5b89de0f5296459b152d,  I4ac93ed29241fee9390fd824452e6632;
reg [fgallag_WDTH -1:0] Ic99c4503bcbcad1099d0c26d3d9161b9,  Id6bb9f52fa37334787904652fbb1bd95;
reg [fgallag_WDTH -1:0] I36119b67ff8b6471d47a6681ce27666b,  I21281177f31dc70c65db2e9a3aa72392;
reg [fgallag_WDTH -1:0] I29103484cf42c813700bcc89a04146c8,  Ia64ddbc7428ff56489b0855ff0fc67a2;
reg [fgallag_WDTH -1:0] I3cef2dada2657f2140d9bdc43f83057b,  I4cebb1a21b9c76387237fe8784f97ac1;
reg [fgallag_WDTH -1:0] I23abb9c83aae42b4b3a330f277ce3c5a,  I3b8cbc445627a75cc4b05aafc8a23cc5;
reg [fgallag_WDTH -1:0] I79b6e7abe2503f1f13195584805dfcb6,  I46c35e4856fb0288a23d9c4c68290ee9;
reg [fgallag_WDTH -1:0] I4d042a3d0026d6b93b5b394034174b00,  I4660e4e54643b4a73afeecea4a4284d5;
reg [fgallag_WDTH -1:0] I92d347131e209dc81a8321d27d38a69e,  I86454d943e7ff4b244882b0f6955d9df;
reg [fgallag_WDTH -1:0] I79c6fd3ceb89abc93f49a67d913505ae,  I3e0245e2c18af49b10a4f2ee38ccdd20;
reg [fgallag_WDTH -1:0] Ieb5038840ac4ab2ebdd9cf6222c15750,  Id34d6ac40408151f201a8b3131463b3b;
reg [fgallag_WDTH -1:0] Id81b8442322f6bdc3728f5459a830aeb,  Ib002905f7b54145ae3dcf7e0f8715b8b;
reg [fgallag_WDTH -1:0] Ie3a852b81ccaf2d520d024dd989caa47,  I3ffe132daa39f108095cd1fd5c38c6d6;
reg [fgallag_WDTH -1:0] I33b0bd948bf4495908c59c2d8f58cf2c,  Ia057defdefe85e4b01cb1acf025fff51;
reg [fgallag_WDTH -1:0] I09a19721c1644f9d1a6eaab84d8dddbe,  I080d693c8cdddee8f9c80ad68d1db1fe;
reg [fgallag_WDTH -1:0] I7065b10d4533cd967733d262d5e5777e,  I55f1644f9601b3553040f8b8ecd84eff;
reg [fgallag_WDTH -1:0] Ie75d8156129eb98d76783e3a6ade280e,  I30ce714aeca130dc1978c6eda3ec0e11;
reg [fgallag_WDTH -1:0] Id3d25ba968ed699bd0b61ee32695edee,  I4ebdb0445ef12223edf4ccf0e4785b01;
reg [fgallag_WDTH -1:0] Ic560d519645177df445db05bad34e60e,  Icd76d18cf8b38caaafc592047ff3b48c;
reg [fgallag_WDTH -1:0] Ia5720f57dcae8ac0b00ac4e4a3c89657,  I51195d2f4e3b638d1f1d226ccf89ccc6;
reg [fgallag_WDTH -1:0] I8cfcf912f60acfc715c63291a8c04729,  Ia29e3ba7f03b070d4381093dcafcdeb9;
reg [fgallag_WDTH -1:0] I6e5f2896cda9b8db3638d2b14cd6ac00,  I2c9a9e255b7ac39f5d6509cdf27f6d4e;
reg [fgallag_WDTH -1:0] I349da988b53307693f1e74a98fa686b6,  I49dd3ecb280e2ea8639a2397343f1700;
reg [fgallag_WDTH -1:0] I47ec23a2e834f9c66f23f1e89eaf8679,  Ia1d516cb29b48f621e47ce669cb9220d;
reg [fgallag_WDTH -1:0] If03782abea72e6519c530636040d2291,  Iecf3c7051c364595cb29b47e8ceae9d7;
reg [fgallag_WDTH -1:0] I512ac9f87b0fc7590f5434fc1e3f0372,  I72fb085a491b61f89d4f95cda02b4b3c;
reg [fgallag_WDTH -1:0] Ia0d98d1391069c78a92be189e60cec14,  I1623b3a676440bab948f5f01c31c87a2;
reg [fgallag_WDTH -1:0] Ic75a566d180368ca17dac6f967fe397d,  Ie83ef8c66f723e3ef386055c5d0b9d8c;
reg [fgallag_WDTH -1:0] Id9acaf5c4d2e0ff41de104ab47e77756,  I858523451a6554f7bc0238638450bb3d;
reg [fgallag_WDTH -1:0] Ic0a4f0637df63f87635fa78c21b2e99e,  I82c65f5d9ca29f356382cf62e638f3a8;
reg [fgallag_WDTH -1:0] I4a61d91e170ec3b767be88ccb343f1ca,  I88222b3d351f2f7334c9f3f22d3f0255;
reg [fgallag_WDTH -1:0] I12a049b431155546b8663137cc66bb9a,  Ide7e980d6331b40896f26f3377d80c32;
reg [fgallag_WDTH -1:0] Ia019f222e96881e643709af1eb85011a,  I2347ec4791ee62d976d13c7c6319e16a;
reg [fgallag_WDTH -1:0] I09be79fb5efca2f460b667770755191b,  Ia5706e1260d5d1b3c625f58c1c2fe509;
reg [fgallag_WDTH -1:0] I53f09f16c58b346a02997b021f882363,  I4c48730b147596406983412e0e6ae556;
reg [fgallag_WDTH -1:0] I19b06a7f2c499994044c7dae5057d8a1,  I7de06231997b971a3acdfe69ebd5a394;
reg [fgallag_WDTH -1:0] Idb57cc9ee60ae36bf3c0117776a46d70,  I70281a4f7bfe2fc5e4a0b91b4194d286;
reg [fgallag_WDTH -1:0] I8c056925751f5cbfd61b1195817d25b1,  Ib95d1aa238c37881c0934c8d22cc79d0;
reg [fgallag_WDTH -1:0] I8b92da1d7f30fa71249623b2bc87b462,  Ib9d8fdfe03633433eab48b80f9d4bae8;
reg [fgallag_WDTH -1:0] I020b3d3e1109655d6f795fd1ecc0a322,  Ibff1757b162a6cba3637e2a0c53d4f57;
reg [fgallag_WDTH -1:0] If0e90362af64ee2a20b44f61aa766fb4,  I69f8f0b916f8d0b4d146e839c19a0756;
reg [fgallag_WDTH -1:0] Ie192f4f4088d17d1f7840213009ca3be,  I0f58fb5960dd9007acf9103e1ef428c0;
reg [fgallag_WDTH -1:0] Ic72e05f3be735d52d9354cb8f43c1cc0,  Ic31af45750c67aca08c2af5f1fdc52d4;
reg [fgallag_WDTH -1:0] I76141646fbd2efad1e121c6e08ac174e,  I81b800210ac62493bcb6993bf20de4f4;
reg [fgallag_WDTH -1:0] I4ac4e1dec3801e462a47f80276b42397,  Idec985d498536ef129885e9baaa69be5;
reg [fgallag_WDTH -1:0] Ifefb5a209dde348266eb66805c0a7d2e,  Ib85fdca5ff6cd6fd13a196d1fb380166;
reg [fgallag_WDTH -1:0] I92c5b8b76f0000bfffa0120f70f1991a,  I64c48585300f968447198fd11396fd71;
reg [fgallag_WDTH -1:0] Ia94fc30c06efdb8ae6f388149d0dad5c,  I9cef63d7e32492a449474355630e84b2;
reg [fgallag_WDTH -1:0] Ifdb73b22fe15d17de645cf8aa3da99e2,  I8d49cc394888a3e49b8e5cd72f2877e5;
reg [fgallag_WDTH -1:0] I0b0e5a5734bd09dfad80a75fca5a763c,  I19030461146fca1f78cdda6d38cd91f1;
reg [fgallag_WDTH -1:0] I73354f6673afdd64f94fe36e146cace0,  I80802c2f239fbc3ed9bff61e9c873550;
reg [fgallag_WDTH -1:0] Ibe0a9cbd6da728e5f7e53081af472ea9,  Idb96776120ec0d249a660e1cdfbf4362;
reg [fgallag_WDTH -1:0] I0edeae6c95ab6198047ded7f3b41efee,  Ib8b1376de13c22be5126d585890438d7;
reg [fgallag_WDTH -1:0] I473cf664c81394c8dab1d7f145b3804b,  I0a617772f4b574bc44555b85eb425b3a;
reg [fgallag_WDTH -1:0] I7201b831890988766bc871eb0fa6e19d,  I3a9c038e7e278e6630b3defab662e10c;
reg [fgallag_WDTH -1:0] Ic772d12c6a9f51ff6cb51bf7d54d1b21,  Ib741e42703c8b7e4ffa9a6fe599e78ec;
reg [fgallag_WDTH -1:0] I16120aeff10370316421751a8f4e9505,  I878e4888b177aa7880c8ab11384db32a;
reg [fgallag_WDTH -1:0] I77146070f8693370d971ec3a91e18f84,  I294424e35f618c68248a468bad92814d;
reg [fgallag_WDTH -1:0] I784fb1f69095ccb95c4bb705539970d8,  If808ebd32478faac57b26b5306292dc4;
reg [fgallag_WDTH -1:0] I2b2174ba9f0956782a3ab584fd11777a,  I122612ac7be83ca897e3d0212c7dcaa1;
reg [fgallag_WDTH -1:0] I8f31a3afb2cc62773332f251278c1153,  I88320212337ea2d63720b17e98675475;
reg [fgallag_WDTH -1:0] Ib2cdf1583fe14fd7b16229572511fd7c,  I777989034e3f2e68b036801349f439ee;
reg [fgallag_WDTH -1:0] Ib04043dbfa7a17abbb728899e2459398,  I20f9fe0be090aee8bf1dcc46f806d73c;
reg [fgallag_WDTH -1:0] Ib1eaa856a32de8ec5107bb40c8611700,  Ie26a8b21d119555a1e9e6b3c41606658;
reg [fgallag_WDTH -1:0] I04ac748d74a312f05ede4d4665042de6,  I47c779e7352c5c5f13cccdd737dc994b;
reg [fgallag_WDTH -1:0] I70ef81ae751a5a7640ce2d4b0ac381c7,  I29f7d07e6ad56f0d6a9b9126d5ebd6bf;
reg [fgallag_WDTH -1:0] I6c64c351f3b91838c0c3c25f3b06d201,  I7ae4796f21cd658ec17c8ff97f369784;
reg [fgallag_WDTH -1:0] I146352e56b780e8cc0f10ac09cee3a2d,  Icae58f7ba349c64263a4465f8de68bd5;
reg [fgallag_WDTH -1:0] I966ffe439dac9390e18e84a65e4b6f11,  Idc1a3fedeccab7f0ee34f79366f5c4e5;
reg [fgallag_WDTH -1:0] Ief16bdfba3e4ab746af015310ebbb6b8,  Ie8117cdb093d8606a07c83ee8e80b388;
reg [fgallag_WDTH -1:0] I0bb8923bb50a4fc7278094a514c79fb6,  I0a65eb60e084d42aa5f5d9d6803068df;
reg [fgallag_WDTH -1:0] I9e93a476f9669fb72f7999a6f0a05c16,  I7f0634ff89c088ca73363e951657ec5a;
reg [fgallag_WDTH -1:0] I0442bb2973db673118791e504be846e4,  Ia45d63e797413cb23c429c7d7a1eef02;
reg [fgallag_WDTH -1:0] Ib00b860d9b3981465aa3bb1f18cfc627,  Ib7b0721390dec3041d5257d0e3df97c3;
reg [fgallag_WDTH -1:0] I6ddab9f5aca020985482b76c25f2f81e,  Ib89de4c510d53bd06fe0f10c7513de04;
reg [fgallag_WDTH -1:0] Idaa6aa87b597a3bcc6275f5f40444057,  I2938e6df94b490c2100ed57268545d36;
reg [fgallag_WDTH -1:0] I1e2ca5efd6735a6e241f9bcade3c2b60,  I8b7353fd85fd2ee67a1df24a9f239f50;
reg [fgallag_WDTH -1:0] I50da8ce0a49993e0b7c16710e68da821,  I66ee7fb42c8ba5991ac6aa8cdb51bf52;
reg [fgallag_WDTH -1:0] Ief43e8dc88393e5a4015033c4021a8e5,  I3ceb68a7f17d021fb3ce01821a19e7d8;
reg [fgallag_WDTH -1:0] Idc4a8277aa0ac4ac35b9fa6b37f198f9,  I649e640596807ec607a1c29006987d98;
reg [fgallag_WDTH -1:0] I4f555c0f5b4b6f79ad394e0f196c8e9f,  Ia67f20bc0f3e32bf1e443bae34efc4b0;
reg [fgallag_WDTH -1:0] I7ddabcd95dfd2719f9e9925598e0cd80,  Ib1af7cd6a6d84431253d818fadb177e4;
reg [fgallag_WDTH -1:0] I007d2500c173825191e1243fc0758203,  I6631364f87a3c0d43c4e1e433b61a132;
reg [fgallag_WDTH -1:0] Icee24ae7d32c16a6b5dd7089f6a63d18,  I8daa733c7e34401a9002dbeef55b89f1;
reg [fgallag_WDTH -1:0] I0d5ad201c17a461d16a13675a0abf874,  Ief1269d4009e33d56efce8d693d3588c;
reg [fgallag_WDTH -1:0] I8cdcb20840d2cafe54bf1a40bb5fdb1c,  I9274d5ddfd1bbfe08138024e1eb81052;
reg [fgallag_WDTH -1:0] I5dce978811c8a3680684eb168992afe7,  If36edf1833e16bf79b7ea16dcc551d2d;
reg [fgallag_WDTH -1:0] Ied4802a1ff9e40f97bd6ed7e5c9af351,  If978d531c028e4c3c00cec8d057703c8;
reg [fgallag_WDTH -1:0] I54c34254efd813baebdff01bb5d9100a,  I1cc0a80d74fe4b030cd838bd32b3cb20;
reg [fgallag_WDTH -1:0] Idf998c5802562dd8ba5cbbe2d8f4eca3,  I0de61810af282ac4baace4ddca69f88c;
reg [fgallag_WDTH -1:0] I5140c93c2312dc879b408cce4db484d3,  I4566be9ae01ab539195295433536bb4e;
reg [fgallag_WDTH -1:0] I0110a5e1c6faa19f5d97ee4b4f763285,  I9ba42ab3f14a648fa7ba73189a272474;
reg [fgallag_WDTH -1:0] I923c20fa85b752d9f31a3476e863c4c5,  I735b9bdb73b8701ec3181c5c08f9637c;
reg [fgallag_WDTH -1:0] I0eb29e587012701bb6ff57aa27d71ecc,  Id88f6239fc5367bf8ce4c1c3bd45f75e;
reg [fgallag_WDTH -1:0] Ib3668e1656878dd9ba2862b988011686,  I78d31cfda6c9de83fbee1581d2cf4330;
reg [fgallag_WDTH -1:0] Id7a758f960bb811f4ebb46662228c33c,  I64ccbe69fe3724b0b97ffc27c7682b0f;
reg [fgallag_WDTH -1:0] I271fa5cfca7bbdafb091c3afcc3a7a41,  Ie29fc0c82ccfe2e936226bbf8a22aa93;
reg [fgallag_WDTH -1:0] I864329472b61fb8580558865bcee6de1,  I9b5a96b0522eb62830257171c98627a0;
reg [fgallag_WDTH -1:0] I78527503b3be9fca973ab9fb7f987f27,  I3b383604747befb7811e7cbda19108f2;
reg [fgallag_WDTH -1:0] I3f50edcfbffa653e39523fb6125d4fd5,  If0b2cc476e6faede63243dc637ef5233;
reg [fgallag_WDTH -1:0] Ib5dd6975eedeed971f4aeaef77f28f1e,  I6e38e23fc4b5a6d9f5990d7f82f6a0c7;
reg [fgallag_WDTH -1:0] Ica77a9f6eb020b850ed2fa38021f33fe,  I0730fb0081845ad1ff057ca56b951d75;
reg [fgallag_WDTH -1:0] I783f912ad4fff3731add8abca943629c,  Id5737f058ffd0a11b2d29f088cf7591b;
reg [fgallag_WDTH -1:0] I1d7c0387f65da7d2ae51250edfc764de,  Ie41e239efec92527dd0d50dbc4dae735;
reg [fgallag_WDTH -1:0] I809a5efeed0db403579d08d520c2c9f1,  Ib906993ed1101ad0992f24c4dae29370;
reg [fgallag_WDTH -1:0] I7649e3988149218a8845000ffe68477f,  Ia9eb0f66bc38056887e1492ee688f373;
reg [fgallag_WDTH -1:0] Iad53806231a0e21d8b1e6b8a22fe3dfb,  I4c6811b2d28239598a23f790a03326fc;
reg [fgallag_WDTH -1:0] I9dcd325f9d12b6495d5b9f050af3c72e,  I29271f07d1108d2c542b60c4296c7195;
reg [fgallag_WDTH -1:0] Ib0d29b4d3693a1487dd507cd4610006f,  I9ac5de9728a0349bdb44341a68adeeec;
reg [fgallag_WDTH -1:0] Ide3d8fa67f76ce3a1762381698b59301,  I3ea1e03eb78be51505b0bdd005aa6e2b;
reg [fgallag_WDTH -1:0] I85818659b37457732130fef9b829758e,  I969fc047ddc46bca31190e0d7f435bd9;
reg [fgallag_WDTH -1:0] Ia8d5826890b3ca20e13dfa917300631b,  I7a23ad071ca3404684d12d2a0f36483d;
reg [fgallag_WDTH -1:0] I6b7c6fa01374134b230ebe6de1602785,  I38083dfdf321de81daef5771d0546525;
reg [fgallag_WDTH -1:0] I4ebeea8273995c7ccb406a5cfedc3ef8,  I894d1f8f86188aea7fea540ac74bd39b;
reg [fgallag_WDTH -1:0] I6521570d5f202bce800b1c49adf3f2ca,  I9d6d3cf2eccd6cba144db2459967a901;
reg [fgallag_WDTH -1:0] Iec61267ecdecf9fe305142fe095a21bb,  I8cec6c5d567ae4efab02118383cbb0cb;
reg [fgallag_WDTH -1:0] Idd383af878d242f7be34d1c9d3efa0e8,  I1cbd09f17301a0bee1cd695a2bde4e1c;
reg [fgallag_WDTH -1:0] I44107557054891b33135a13058e00649,  Ie767f5975b691400b250054bcf08867a;
reg [fgallag_WDTH -1:0] I013496291a38e851842de8ea28b540ba,  I54b29fec4a88bc1e03197a0c55b875db;
reg [fgallag_WDTH -1:0] I54e8b21c865654527ee0720a72ef1cd0,  Ib0c39d1e2cffc0326a30bfd0733075a7;
reg [fgallag_WDTH -1:0] Ia40d6a1517b7b0a79c88646d209263dc,  Ib4dee5c8efd8022bd9c3f9bf8d5e328b;
reg [fgallag_WDTH -1:0] I1e10e22806a41d12b8c6328dbd9471df,  Iae316011740707036b166a712b32f2e2;
reg [fgallag_WDTH -1:0] If96824bc7f67bd2bce941ce96559867e,  I3ae123c41c91d9b53a70aa3e4793be9b;
reg [fgallag_WDTH -1:0] Ib252f7e32a3780abfb1a3e9285d0ed56,  If4ccd39857a7317488e9215271db7210;
reg [fgallag_WDTH -1:0] I192fd55ca87b7cb2277aca900d015b04,  Ief6d7060558cf2ccd8d561ec17b846d5;
reg [fgallag_WDTH -1:0] Ie973db372fd3127653d6c63a551a8c0c,  I2a5d6b55814dbead5a30d961f8f7b478;
reg [fgallag_WDTH -1:0] I3446695b823b258ade0a7ac2aa9d61d7,  Ie03342fcc484bd9f1c934e675c9f6ec4;
reg [fgallag_WDTH -1:0] Iea584b5174273f9082695eec0d7a8ab1,  I195e5182b2d3136ff3ef4572cb4b88da;
reg [fgallag_WDTH -1:0] I6d7f0d64776ea582e326ca3b008f2b35,  Idb2832cb2e894a8c02e7dab1dccdef87;
reg [fgallag_WDTH -1:0] Ifc32a10a9fcddca15eeef7d093d1401a,  I5462aaf13ac6e9761929c998fff0b87a;
reg [fgallag_WDTH -1:0] I84db677284b3e4bf9feddc2af30e9ad3,  I8f9db21a5dea66f9865796d164f689ea;
reg [fgallag_WDTH -1:0] Ia04c9bc6fc469c62a3645e0e691b3897,  I31949043c0e635f71f9785c21d713c96;
reg [fgallag_WDTH -1:0] Ib7457f82785a56cbcb5be6c0432641b7,  I2135e15ed882d1293741fd593369f88d;
reg [fgallag_WDTH -1:0] I42a4d0da5f0b890624310c94b32f1a27,  I8cfec980374c11bdc4947a8c69a55728;
reg [fgallag_WDTH -1:0] I08a589b0a34d88ac456d6cf40da0f5ae,  I5e298171856ae5526301f6d5084f2796;
reg [fgallag_WDTH -1:0] I2f1e3460880499c961fcb244ca935f3b,  Ifc2714ac9c0b998653c2a1b5e9199d5d;
reg [fgallag_WDTH -1:0] Ie7f199c3586f87a1cdba687bd880497e,  I1b7e4002a74d5f33e7d0168ed06aaa2d;
reg [fgallag_WDTH -1:0] Ia3518f4b7c1b0aa2a864d5ce53158ce8,  Ib868c2b4eb4dd68231ed56d937dd4804;
reg [fgallag_WDTH -1:0] Id2616c8625d0a75ea0946506034955ca,  Ibe26ea03448b95798236cf228817dfd0;
reg [fgallag_WDTH -1:0] Ic3c6cbf9171a81f229a0fb9efd57b000,  I4ebe3a4a45add9d58508c58a27a5d46d;
reg [fgallag_WDTH -1:0] If63bcb026b347506aff08fda75ac7c43,  I21d9dac9d09da39f435c7082dca90127;
reg [fgallag_WDTH -1:0] Ia79c0c66c81e60806fe3df0addd5608d,  I69e220ebbcd0c48f5cb1cf16fc33fa57;
reg [fgallag_WDTH -1:0] I0695fe1981c8019decb9873e186934ae,  I8546eab32336885c49882f192be9904c;
reg [fgallag_WDTH -1:0] Ic334a0e64e305848782becce03c85d2b,  Id4da583323a66a1333d836c5f7bba069;
reg [fgallag_WDTH -1:0] If737be717332ee2670d2c6736d9e0a2f,  I8c50bd38d4339a6ae19e13db1a1994e9;
reg [fgallag_WDTH -1:0] I66316458bfbdf6b24cdc0cd7396c84f6,  Ia19b6c2a9b73f96a351eca1700079c42;
reg [fgallag_WDTH -1:0] Ib23a5c11d42408a0f4a6d314a670da51,  Ia98d1ff0d0dac6a253cf48ab85e0eb75;
reg [fgallag_WDTH -1:0] I792738baad12910007da8123fa0ac415,  Ie63e6f9d56e6b192f0703cff4813499d;
reg [fgallag_WDTH -1:0] I64f43975f3065e3c7cfed15d5dbc8d72,  I0b963cc516bb0de18221dd724864d795;
reg [fgallag_WDTH -1:0] I4c0a3a24dcfac4edcdf29847761a8fb8,  If1ede61a06a91d3ae1874816901896de;
reg [fgallag_WDTH -1:0] I65fa0e67f8ee4669bba74ece0c565a0d,  I7f856b89e8b206458e96335076d80c69;
reg [fgallag_WDTH -1:0] I6bea44d0467b461aa22c3ddcb1d8f886,  I8cb21da337ae4059685b273b50116a0d;
reg [fgallag_WDTH -1:0] I582cb5f8b17099f479f297c5475542c1,  I72569b57d65e91bcea79d0682c51c4a7;
reg [fgallag_WDTH -1:0] I6cba6eca48f199379e62726b4ac271f8,  I61e50081c686dfbcb684ae83ed3a53c6;
reg [fgallag_WDTH -1:0] I57cfe42eafe8357ec85906472dec3f36,  Iad3645f6fa7141133b12534c70efc80c;
reg [fgallag_WDTH -1:0] Iec7bf02aeaa8630497275c7eccab7667,  I62c110783203a19c372c6aeda18ee18d;
reg [fgallag_WDTH -1:0] I388c7af9494f4c425621d3abfdf72b63,  Id7216252c1febf54691e626861f6215c;
reg [fgallag_WDTH -1:0] I2622bb3685a7d6a297506eac3efb9c08,  Ide229e0c521de0ffd39c67a6f078766d;
reg [fgallag_WDTH -1:0] If025bad83549d872a3fc9c44248174c8,  Id25c2945168c44ec9f0a4bb2dc6aaf68;
reg [fgallag_WDTH -1:0] I3440574538a5d7dd250fbc98d574548b,  I68a5c8b30e8d3e5b0d710c7f306304ec;
reg [fgallag_WDTH -1:0] Ibe30f2ceb078297737ce1444c1e6c524,  I2b3c4fca6b0feb6fd829e9cbbe9d7142;
reg [fgallag_WDTH -1:0] Ifbd6f1ac3bb594aad652d4e3cac018e1,  Ifec9e94824843f4cd8d623219278f87a;
reg [fgallag_WDTH -1:0] Ie41d26b8a9ac93a09ece53b2af8c855e,  I7858226bb4feb944c5feaa52f2b51034;
reg [fgallag_WDTH -1:0] I497c3961e446544a8031e8013ca80ad5,  I3b39fa7f2ad7920296a8e01cc9c12cd6;
reg [fgallag_WDTH -1:0] I6ab9d8eb7b8e3454b01a8e67a410624c,  I1201c86e1f6f9e890181790896c4afa4;
reg [fgallag_WDTH -1:0] Icd351f2625b163cee904fa4e446d0cc4,  I8280be337ee3709b32502e07241156e3;
reg [fgallag_WDTH -1:0] I79c9be2982685762d0907583f9f459e2,  I3920223ae6d1a6d2ff327f53933ecad4;
reg [fgallag_WDTH -1:0] Idc20427e979f3d5c03d7dd947cb4df84,  Ica4ec266d79edda776095c95c3c20630;
reg [fgallag_WDTH -1:0] Ie8abbb597c8132b8e23936a5bc035041,  Id23811d7cf32f6c5c63ce2782da15720;
reg [fgallag_WDTH -1:0] I42b0c89a558950f658440d8f9916b42f,  I6df32fcf5553d3b899e6a67a35b852b5;
reg [fgallag_WDTH -1:0] I5a4d5a128b1fedabfdc39cb019359106,  I7a01b2b85d70a35d44836e181a22b322;
reg [fgallag_WDTH -1:0] I8227a9907c39647a4cef8e883d487913,  Ib725193cf104f9b56c3211df12867643;
reg [fgallag_WDTH -1:0] Icb2a399b8ac8449ff9ff8e5986aac03d,  I45b1d972b2a5028cc340988f7c37f2e0;
reg [fgallag_WDTH -1:0] I933a5eb08d4d1445f167a74db5fbdc75,  I186a56ca3712df6983eb742d7d80a37e;
reg [fgallag_WDTH -1:0] I9c046caddde3b171774d3eba258190f0,  I389856ba7ca6568e4ead3483c3e52353;
reg [fgallag_WDTH -1:0] Ic8f12fefb9c055923e2842aeca48765f,  I66b39fb4c54ab32b2c876813544ff6bc;
reg [fgallag_WDTH -1:0] I26631e7940eb983e49a9313da628e23a,  I591624fd56ff315e0084af5af206cf8e;
reg [fgallag_WDTH -1:0] I7fac6686ca9a63213ec3cdee4b812daa,  I3994dd74d52d8957e443e869cbbf7184;
reg [fgallag_WDTH -1:0] I1960eba710ca20ef749501b02fd3b0bd,  I92793401ab28d5ed265775c0d165dfe5;
reg [fgallag_WDTH -1:0] Ie1f5cc89163ee091f938a4c3edaca65b,  Ic499c718cc4866eb8536d66ae4fae0e4;
reg [fgallag_WDTH -1:0] I63e7cf958a0de50d3299d2077d8cb192,  I3c28bfe18fb1543683ae264c396a0207;
reg [fgallag_WDTH -1:0] I50c2132c2b5e60af7ba2b9be8c90d9a4,  I083aca08b0d0bd2622d0f7b6b2aaeb99;
reg [fgallag_WDTH -1:0] If1243756e31d0a56b6666cad5b21f731,  I2fd3c0dfd43b65e2fe8afd3368a50fc5;
reg [fgallag_WDTH -1:0] I92c03e59c3f96f63800051762f6949c0,  I58332f7615e647e757033f6b643c21a4;
reg [fgallag_WDTH -1:0] I488d337ed967adebd6c580b7203991b5,  I22bbdf426df953feb5acede78c31b9b2;
reg [fgallag_WDTH -1:0] I32aa0d9a082eb6a595467f3c7f36a3f7,  Ia9f7a93a673c49ef3bfffd6fcadf845a;
reg [fgallag_WDTH -1:0] Iec440f37d189fbcd4c06cf34344c4439,  I687ab1878d38c7c988507163c8a60070;
reg [fgallag_WDTH -1:0] I66d815daa51bcda0d549dbcc9c027195,  I9efb470a3342962583f19eaec3a0ecd7;
reg [fgallag_WDTH -1:0] I192d10feae906d5ef90b4a90398d3ced,  Id7f7499e9b3f529781f4aba6e63490ac;
reg [fgallag_WDTH -1:0] I1d8d269f64d0d3041bc69d879a3654ab,  I88e14285aa13b58457c58439ad1c8c87;
reg [fgallag_WDTH -1:0] I5fce715f064098fe4685479aede832e7,  I730aeccac38e1622c684c468f8cb29f4;
reg [fgallag_WDTH -1:0] I1b65989684c087f328e3fb58d3a3395e,  I9427589efc5ae29474734dcc6e36ea81;
reg [fgallag_WDTH -1:0] I5352562c002801df06f847362d347180,  Iba910435a91ee873f76fa3ec9ac9c3d3;
reg [fgallag_WDTH -1:0] I176397bab05ee39f7d54a28c5f74c3cc,  Ia3c2d3cea56571481655cc77ee025558;
wire start_d_fgallag0x00000;
reg I99ba3451537a2876c9f585f72911bc4f;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 I53846946a877f30f72076ee6f633a0e5 <= 'h0;
 I5d219e3294f2763bc17209a55758ab54 <= 'h0;
 I6273ee09aacad20f733530af1a987ff3 <= 'h0;
 Ie0f63a67c0a6ec07e7bcb943e7804f9a <= 'h0;
 I7b83ef4e45fe20e023e08aa3e56bb21e <= 'h0;
 Ibc8f334cefc147e5c58e7542d26fbe2b <= 'h0;
 I662a566f576ee431bced6f852294713e <= 'h0;
 I2a4bc966b71864a79f582727f122ab60 <= 'h0;
 I23d9f47edf51ff1c2a6275531a1f66be <= 'h0;
 Id46ae2d16f43af3529d91eb4d6bd098e <= 'h0;
 I51298122656d9b893c1dbb33a281f134 <= 'h0;
 I22e0a22ed1768671dbe3caef8ac499cb <= 'h0;
 Ifb9327c663379f77471d460eced9c1b7 <= 'h0;
 Id6080749dda3cd29c1ce36ab39759709 <= 'h0;
 I532fd8f9065e524727e276a1a8408008 <= 'h0;
 I1f0b23c673ff55115f55c80a970172fc <= 'h0;
 I9f99ad4587fb6907b3804c11125f738f <= 'h0;
 I719bd7e94d4289c6fd59bb91ee559980 <= 'h0;
 I9103b57e3550cb68266ba8b102e50dfd <= 'h0;
 I89fca1c1832813b84cafe145377d7b5e <= 'h0;
 Ie17de6e388779502a143212813a50317 <= 'h0;
 Ifcc046128364b8da7bc3d9ddab96a061 <= 'h0;
 Iabe4b7a23f682ed62162dfde9e15d6cf <= 'h0;
 I734eaef0b7d7f6ae5d668ac9b374ff51 <= 'h0;
 I0e0e9fdfeb3e2115deb903b973217384 <= 'h0;
 Ibfd2fd7aa2426054706d0c4e4c0a7cba <= 'h0;
 I0906247e3ba96971232bc42185c9a9b8 <= 'h0;
 Ia3908fda391d7caf1b479d9655164c30 <= 'h0;
 I820e95cdc583108195e8dd0e2d1f4b7f <= 'h0;
 Ibdf5c2c57269da1b04748a59802c8e2a <= 'h0;
 Idd85c8c853438679d99bed4d0ba46af7 <= 'h0;
 I4d617d0b669b3ff1b08dcd4b7440af33 <= 'h0;
 I60d579b60b02f9fc14e98d7d0eb54c18 <= 'h0;
 Ic1a37750fc3d7eb08ad649de157f45a9 <= 'h0;
 I0c13ec63e7208b35a1d4511e1da29fa3 <= 'h0;
 If10c9545a713996735934c5f15cf5365 <= 'h0;
 Ic475963164a956dd24ede91e9d61003d <= 'h0;
 I42001c4b6ab9fb03489ca25defb6c222 <= 'h0;
 Idcfb16adf2996c8cb51e402daafd1734 <= 'h0;
 I924108a2723afd07735574a6f4ebe671 <= 'h0;
 If9fd9ae380997e75ebed2ddd3f93e76f <= 'h0;
 Ief876b7b2af1fbed4d3f457cdb46e0d9 <= 'h0;
 Id2bd196ca25e1a077fb2a9207f143c01 <= 'h0;
 I926e2a038d48db29b5ce215cd6cf6a04 <= 'h0;
 I4ba2cfd94590dee1723ce63afd0926ab <= 'h0;
 I0d42326464ae4c3a55038e0343cebf5a <= 'h0;
 If05fde321fd1456422550f5c3903b826 <= 'h0;
 I41ec48a5a1d657a6266b8f845550d0c2 <= 'h0;
 I76473b4885d423029324fe74ed13d6ed <= 'h0;
 I8ef2366947e3f1352f3874e4ac58d7b2 <= 'h0;
 I874c1e455f85e617a5032ec230fdfdc5 <= 'h0;
 I16d6b6b19890a6bbdf15ddc27717aa30 <= 'h0;
 I6af6d04126eec9eb91e5653cc95c9ef3 <= 'h0;
 If501a668f24fd62a69d0e3c253739c79 <= 'h0;
 I9b70e215a2a1578811b40c669826d41a <= 'h0;
 I26d82966efbe51e03edcd66a5a507ebb <= 'h0;
 I2e4afb94e4af76b4e3d859815bb338fb <= 'h0;
 Ie19faf5d037b74974102c386a13f4946 <= 'h0;
 I2d56338af0755ae5c4ef71ddad3112b1 <= 'h0;
 I99ab212db901b0e65eb33be27c46bd19 <= 'h0;
 If8c09c14d78b1deaf76df6f4de910c64 <= 'h0;
 I1b0ccac0f5cc741403fd6e680899f96f <= 'h0;
 I38153cd88e8b2452977d7dc9b9f44a74 <= 'h0;
 Ic32064fc62eb1cdcdf416a6fe78becfd <= 'h0;
 Ic10eb104fe38a176a51507e748406958 <= 'h0;
 I979fd1b01c99b76a4ff2d0abfb0c2ae9 <= 'h0;
 Ibe530a86c501fbc8dba64ed24806bdf4 <= 'h0;
 If03531315c68272f7de2b0e969770f48 <= 'h0;
 I20160f4e380b0920bcb30a0321b7bfa8 <= 'h0;
 I2bbbe5d3a72af5f654976a7fde2d2d16 <= 'h0;
 I70f4396800d2cb065ad5fe655bacbfd0 <= 'h0;
 If27a0187d1188cf7a8aba100a90cb069 <= 'h0;
 I8994866d080b1befe414fea347e7e74a <= 'h0;
 Iab6971c846299eec0a5cc93ad10e569c <= 'h0;
 I8730924fec54ffaa78a0ffea7e8386ba <= 'h0;
 I338fb9183219691c6b50e6a824fcb14c <= 'h0;
 I1a3d82eaf2fc9235163c0a50765f4ef5 <= 'h0;
 I922539f8d9ffc119ed3a5c92a21f149e <= 'h0;
 I3bc0f1eaad327d5990adb826e54c6d2f <= 'h0;
 I3009d4cc0371f83e6bec8fb38ae461bd <= 'h0;
 I2e0ae02d7a3cdfa36e8645cc7dd0bce6 <= 'h0;
 If2c59f326f3658dee0fd3b048af14cb7 <= 'h0;
 I04431bd4be4601d3cb700c0cd6d9fd24 <= 'h0;
 I7a6fe8c804087a19e32e760f50e3edfa <= 'h0;
 I979817e250e46dcc05f8a6690c2380f9 <= 'h0;
 I3bbb836eee6b5e10fe55879f8620b888 <= 'h0;
 I8bc5128382cbffa289caec56f9b4a3f3 <= 'h0;
 Iee4dafc9d42609fae74410897f29a78d <= 'h0;
 I4ea5b39ed827d8d4618bcfd9283dfa83 <= 'h0;
 I19aa6440394778642eb50f3b94098ea3 <= 'h0;
 I0653a9ef861e5d8af22d120172c2dc03 <= 'h0;
 Ie0aafaeee1abf6d27a70535385ab88b5 <= 'h0;
 I1583cdcd13120f953691a5a60ee72b11 <= 'h0;
 I8080b45a37a3de79ccb338f353f19529 <= 'h0;
 I9bd98a9d18ce7c07e85287f6b80bfd31 <= 'h0;
 Ife85d240c60084dce9b3d7cd87060727 <= 'h0;
 I11f2e4eafc706b43c10a26edc8567052 <= 'h0;
 Iad3a9febf269d9607eedf29912b04af9 <= 'h0;
 I75705fa2cc0ac0577570501510e4e0fc <= 'h0;
 I7674ab7538766e842366dd08ddbbcb28 <= 'h0;
 I8cefcac1f7fa2df45bb8a2f3d64f99c3 <= 'h0;
 I5fd378ba266fd930a839cad56e500ef4 <= 'h0;
 I71a33ca1c7d18d5089d08a8476c8baf7 <= 'h0;
 Ic85b012b9fa77becd419cac0f3692aed <= 'h0;
 I0ae9b4ca5ebb5f3d2e8b02884069e4e7 <= 'h0;
 Ief312304eec0415d1ab208ed6726dd12 <= 'h0;
 Icb9ebf1f5becaede273da59f466506ac <= 'h0;
 I465b9607a8dad0f1c499318d04f42aea <= 'h0;
 I2523c109974807b3b1c0f4b34693e255 <= 'h0;
 Ib4e3121afd90b877b94c4c7cd29e9334 <= 'h0;
 Ibfb66b89c59008f3d4497ee16dad6712 <= 'h0;
 I2d042c4ef15b2f3bdebbc7cbd6c00a1f <= 'h0;
 I489d1b46970800e9684c68b439c15be1 <= 'h0;
 I835143e23243f3fd25cc1ab0ba5c123a <= 'h0;
 I028ef05ea84be3bc45c518f4f45653d2 <= 'h0;
 Ia5a39eeda95dfdb2ab8b55ea9f8b62c5 <= 'h0;
 If5a85945ad1f8d9bdc9213c5ae2c890f <= 'h0;
 I6011a5fc7b168a28fc9a45f796629b59 <= 'h0;
 Ie703b5f1eeedaaaddf56ded14b1765bc <= 'h0;
 I21f34fbc269f5424ea30334ff7ab54f5 <= 'h0;
 I07b47fce56edeb30319038e3a093efd7 <= 'h0;
 I24e7e5c391285f28c20f74820a05b552 <= 'h0;
 Iee1b23b99f7de56829706633297a0513 <= 'h0;
 Ib4b61d3293900c38e8aa7df0a617b476 <= 'h0;
 Ifd5fcb1552fb372ae203fd0166d3df2c <= 'h0;
 Ibb2fb63aef1d336dfa829cd5ab3675b7 <= 'h0;
 I1672371cf33b259cf87210cc49aa35c8 <= 'h0;
 Ia34735ee7f7ca164c2ae71980060f56b <= 'h0;
 I2372d0a72998f0630e994aa3e1c20ff4 <= 'h0;
 I8e363e0bd65cae9725cdd70e46778fee <= 'h0;
 Id6af962a16ff79ac6e9da3b4518b80b2 <= 'h0;
 I7fc8c9245183d05370746c9b2fdabd0f <= 'h0;
 I693f2c9a5d4da90c3105876991c4f4ba <= 'h0;
 Id6c07cd1f9f428b0d971639939b9eb8e <= 'h0;
 Id6561e53aa8f9fd116159969afaa20ae <= 'h0;
 I8267af03225d6d1155142645ad7f53a8 <= 'h0;
 I567872d8892064b62caeb3dcdc39e89c <= 'h0;
 I5072b405191b837596b5efe4ec159519 <= 'h0;
 Ia4e5d30bc160c1f72c8f39cdcd13e5a4 <= 'h0;
 Ic46dd8ff5a79971f7c22f4be0f1f4b23 <= 'h0;
 Ifdd13523ba0ce3329e3aca49a0a36385 <= 'h0;
 Ib449b5d80a7f5a1c5d0d3784d8f236b6 <= 'h0;
 I134d223e71b68cc9c76379f1368fb0f1 <= 'h0;
 Ifa82272c492ce1ed4b223c0cb2b135e1 <= 'h0;
 Ie501d0f392be1309df48c1616ace5a27 <= 'h0;
 I29468f8318cd5bebb5cea27e1ee57b7f <= 'h0;
 Ie3f06a529d5f22198b3b33d649b740e1 <= 'h0;
 I6740505fac3e83de4a6525ac9cf489d1 <= 'h0;
 I0456541b6e82ffeb05fc4052fafc41f7 <= 'h0;
 I6d5739cf589ed46b6f57075a3b2a974d <= 'h0;
 Iabe05603679da24a44565e756adc0881 <= 'h0;
 Icaed4c0a915898eea654ab6f93973ff3 <= 'h0;
 I98805e117c2f4ba4a8f6c2755ebe1fee <= 'h0;
 I766076681dc49b817ec9302eae86d64b <= 'h0;
 Ia82b6e01034a63c2a1a446029f58f1c6 <= 'h0;
 I05de7fd67a0e226201b563fa6c50f362 <= 'h0;
 I8df8f128712fe5445a97566f8f29ecd4 <= 'h0;
 Iae9103582be213e81ea0a25e5d49004f <= 'h0;
 Ibcab213dbb173403005b3d65f780fa2d <= 'h0;
 Ic59b57cadd4b8cbe63f996111e9211b1 <= 'h0;
 Ide1a993a1dfca37107fc81e985714d93 <= 'h0;
 I7004a1bc0ec2272163d33907d21616ea <= 'h0;
 I4ac93ed29241fee9390fd824452e6632 <= 'h0;
 Id6bb9f52fa37334787904652fbb1bd95 <= 'h0;
 I21281177f31dc70c65db2e9a3aa72392 <= 'h0;
 Ia64ddbc7428ff56489b0855ff0fc67a2 <= 'h0;
 I4cebb1a21b9c76387237fe8784f97ac1 <= 'h0;
 I3b8cbc445627a75cc4b05aafc8a23cc5 <= 'h0;
 I46c35e4856fb0288a23d9c4c68290ee9 <= 'h0;
 I4660e4e54643b4a73afeecea4a4284d5 <= 'h0;
 I86454d943e7ff4b244882b0f6955d9df <= 'h0;
 I3e0245e2c18af49b10a4f2ee38ccdd20 <= 'h0;
 Id34d6ac40408151f201a8b3131463b3b <= 'h0;
 Ib002905f7b54145ae3dcf7e0f8715b8b <= 'h0;
 I3ffe132daa39f108095cd1fd5c38c6d6 <= 'h0;
 Ia057defdefe85e4b01cb1acf025fff51 <= 'h0;
 I080d693c8cdddee8f9c80ad68d1db1fe <= 'h0;
 I55f1644f9601b3553040f8b8ecd84eff <= 'h0;
 I30ce714aeca130dc1978c6eda3ec0e11 <= 'h0;
 I4ebdb0445ef12223edf4ccf0e4785b01 <= 'h0;
 Icd76d18cf8b38caaafc592047ff3b48c <= 'h0;
 I51195d2f4e3b638d1f1d226ccf89ccc6 <= 'h0;
 Ia29e3ba7f03b070d4381093dcafcdeb9 <= 'h0;
 I2c9a9e255b7ac39f5d6509cdf27f6d4e <= 'h0;
 I49dd3ecb280e2ea8639a2397343f1700 <= 'h0;
 Ia1d516cb29b48f621e47ce669cb9220d <= 'h0;
 Iecf3c7051c364595cb29b47e8ceae9d7 <= 'h0;
 I72fb085a491b61f89d4f95cda02b4b3c <= 'h0;
 I1623b3a676440bab948f5f01c31c87a2 <= 'h0;
 Ie83ef8c66f723e3ef386055c5d0b9d8c <= 'h0;
 I858523451a6554f7bc0238638450bb3d <= 'h0;
 I82c65f5d9ca29f356382cf62e638f3a8 <= 'h0;
 I88222b3d351f2f7334c9f3f22d3f0255 <= 'h0;
 Ide7e980d6331b40896f26f3377d80c32 <= 'h0;
 I2347ec4791ee62d976d13c7c6319e16a <= 'h0;
 Ia5706e1260d5d1b3c625f58c1c2fe509 <= 'h0;
 I4c48730b147596406983412e0e6ae556 <= 'h0;
 I7de06231997b971a3acdfe69ebd5a394 <= 'h0;
 I70281a4f7bfe2fc5e4a0b91b4194d286 <= 'h0;
 Ib95d1aa238c37881c0934c8d22cc79d0 <= 'h0;
 Ib9d8fdfe03633433eab48b80f9d4bae8 <= 'h0;
 Ibff1757b162a6cba3637e2a0c53d4f57 <= 'h0;
 I69f8f0b916f8d0b4d146e839c19a0756 <= 'h0;
 I0f58fb5960dd9007acf9103e1ef428c0 <= 'h0;
 Ic31af45750c67aca08c2af5f1fdc52d4 <= 'h0;
 I81b800210ac62493bcb6993bf20de4f4 <= 'h0;
 Idec985d498536ef129885e9baaa69be5 <= 'h0;
 Ib85fdca5ff6cd6fd13a196d1fb380166 <= 'h0;
 I64c48585300f968447198fd11396fd71 <= 'h0;
 I9cef63d7e32492a449474355630e84b2 <= 'h0;
 I8d49cc394888a3e49b8e5cd72f2877e5 <= 'h0;
 I19030461146fca1f78cdda6d38cd91f1 <= 'h0;
 I80802c2f239fbc3ed9bff61e9c873550 <= 'h0;
 Idb96776120ec0d249a660e1cdfbf4362 <= 'h0;
 Ib8b1376de13c22be5126d585890438d7 <= 'h0;
 I0a617772f4b574bc44555b85eb425b3a <= 'h0;
 I3a9c038e7e278e6630b3defab662e10c <= 'h0;
 Ib741e42703c8b7e4ffa9a6fe599e78ec <= 'h0;
 I878e4888b177aa7880c8ab11384db32a <= 'h0;
 I294424e35f618c68248a468bad92814d <= 'h0;
 If808ebd32478faac57b26b5306292dc4 <= 'h0;
 I122612ac7be83ca897e3d0212c7dcaa1 <= 'h0;
 I88320212337ea2d63720b17e98675475 <= 'h0;
 I777989034e3f2e68b036801349f439ee <= 'h0;
 I20f9fe0be090aee8bf1dcc46f806d73c <= 'h0;
 Ie26a8b21d119555a1e9e6b3c41606658 <= 'h0;
 I47c779e7352c5c5f13cccdd737dc994b <= 'h0;
 I29f7d07e6ad56f0d6a9b9126d5ebd6bf <= 'h0;
 I7ae4796f21cd658ec17c8ff97f369784 <= 'h0;
 Icae58f7ba349c64263a4465f8de68bd5 <= 'h0;
 Idc1a3fedeccab7f0ee34f79366f5c4e5 <= 'h0;
 Ie8117cdb093d8606a07c83ee8e80b388 <= 'h0;
 I0a65eb60e084d42aa5f5d9d6803068df <= 'h0;
 I7f0634ff89c088ca73363e951657ec5a <= 'h0;
 Ia45d63e797413cb23c429c7d7a1eef02 <= 'h0;
 Ib7b0721390dec3041d5257d0e3df97c3 <= 'h0;
 Ib89de4c510d53bd06fe0f10c7513de04 <= 'h0;
 I2938e6df94b490c2100ed57268545d36 <= 'h0;
 I8b7353fd85fd2ee67a1df24a9f239f50 <= 'h0;
 I66ee7fb42c8ba5991ac6aa8cdb51bf52 <= 'h0;
 I3ceb68a7f17d021fb3ce01821a19e7d8 <= 'h0;
 I649e640596807ec607a1c29006987d98 <= 'h0;
 Ia67f20bc0f3e32bf1e443bae34efc4b0 <= 'h0;
 Ib1af7cd6a6d84431253d818fadb177e4 <= 'h0;
 I6631364f87a3c0d43c4e1e433b61a132 <= 'h0;
 I8daa733c7e34401a9002dbeef55b89f1 <= 'h0;
 Ief1269d4009e33d56efce8d693d3588c <= 'h0;
 I9274d5ddfd1bbfe08138024e1eb81052 <= 'h0;
 If36edf1833e16bf79b7ea16dcc551d2d <= 'h0;
 If978d531c028e4c3c00cec8d057703c8 <= 'h0;
 I1cc0a80d74fe4b030cd838bd32b3cb20 <= 'h0;
 I0de61810af282ac4baace4ddca69f88c <= 'h0;
 I4566be9ae01ab539195295433536bb4e <= 'h0;
 I9ba42ab3f14a648fa7ba73189a272474 <= 'h0;
 I735b9bdb73b8701ec3181c5c08f9637c <= 'h0;
 Id88f6239fc5367bf8ce4c1c3bd45f75e <= 'h0;
 I78d31cfda6c9de83fbee1581d2cf4330 <= 'h0;
 I64ccbe69fe3724b0b97ffc27c7682b0f <= 'h0;
 Ie29fc0c82ccfe2e936226bbf8a22aa93 <= 'h0;
 I9b5a96b0522eb62830257171c98627a0 <= 'h0;
 I3b383604747befb7811e7cbda19108f2 <= 'h0;
 If0b2cc476e6faede63243dc637ef5233 <= 'h0;
 I6e38e23fc4b5a6d9f5990d7f82f6a0c7 <= 'h0;
 I0730fb0081845ad1ff057ca56b951d75 <= 'h0;
 Id5737f058ffd0a11b2d29f088cf7591b <= 'h0;
 Ie41e239efec92527dd0d50dbc4dae735 <= 'h0;
 Ib906993ed1101ad0992f24c4dae29370 <= 'h0;
 Ia9eb0f66bc38056887e1492ee688f373 <= 'h0;
 I4c6811b2d28239598a23f790a03326fc <= 'h0;
 I29271f07d1108d2c542b60c4296c7195 <= 'h0;
 I9ac5de9728a0349bdb44341a68adeeec <= 'h0;
 I3ea1e03eb78be51505b0bdd005aa6e2b <= 'h0;
 I969fc047ddc46bca31190e0d7f435bd9 <= 'h0;
 I7a23ad071ca3404684d12d2a0f36483d <= 'h0;
 I38083dfdf321de81daef5771d0546525 <= 'h0;
 I894d1f8f86188aea7fea540ac74bd39b <= 'h0;
 I9d6d3cf2eccd6cba144db2459967a901 <= 'h0;
 I8cec6c5d567ae4efab02118383cbb0cb <= 'h0;
 I1cbd09f17301a0bee1cd695a2bde4e1c <= 'h0;
 Ie767f5975b691400b250054bcf08867a <= 'h0;
 I54b29fec4a88bc1e03197a0c55b875db <= 'h0;
 Ib0c39d1e2cffc0326a30bfd0733075a7 <= 'h0;
 Ib4dee5c8efd8022bd9c3f9bf8d5e328b <= 'h0;
 Iae316011740707036b166a712b32f2e2 <= 'h0;
 I3ae123c41c91d9b53a70aa3e4793be9b <= 'h0;
 If4ccd39857a7317488e9215271db7210 <= 'h0;
 Ief6d7060558cf2ccd8d561ec17b846d5 <= 'h0;
 I2a5d6b55814dbead5a30d961f8f7b478 <= 'h0;
 Ie03342fcc484bd9f1c934e675c9f6ec4 <= 'h0;
 I195e5182b2d3136ff3ef4572cb4b88da <= 'h0;
 Idb2832cb2e894a8c02e7dab1dccdef87 <= 'h0;
 I5462aaf13ac6e9761929c998fff0b87a <= 'h0;
 I8f9db21a5dea66f9865796d164f689ea <= 'h0;
 I31949043c0e635f71f9785c21d713c96 <= 'h0;
 I2135e15ed882d1293741fd593369f88d <= 'h0;
 I8cfec980374c11bdc4947a8c69a55728 <= 'h0;
 I5e298171856ae5526301f6d5084f2796 <= 'h0;
 Ifc2714ac9c0b998653c2a1b5e9199d5d <= 'h0;
 I1b7e4002a74d5f33e7d0168ed06aaa2d <= 'h0;
 Ib868c2b4eb4dd68231ed56d937dd4804 <= 'h0;
 Ibe26ea03448b95798236cf228817dfd0 <= 'h0;
 I4ebe3a4a45add9d58508c58a27a5d46d <= 'h0;
 I21d9dac9d09da39f435c7082dca90127 <= 'h0;
 I69e220ebbcd0c48f5cb1cf16fc33fa57 <= 'h0;
 I8546eab32336885c49882f192be9904c <= 'h0;
 Id4da583323a66a1333d836c5f7bba069 <= 'h0;
 I8c50bd38d4339a6ae19e13db1a1994e9 <= 'h0;
 Ia19b6c2a9b73f96a351eca1700079c42 <= 'h0;
 Ia98d1ff0d0dac6a253cf48ab85e0eb75 <= 'h0;
 Ie63e6f9d56e6b192f0703cff4813499d <= 'h0;
 I0b963cc516bb0de18221dd724864d795 <= 'h0;
 If1ede61a06a91d3ae1874816901896de <= 'h0;
 I7f856b89e8b206458e96335076d80c69 <= 'h0;
 I8cb21da337ae4059685b273b50116a0d <= 'h0;
 I72569b57d65e91bcea79d0682c51c4a7 <= 'h0;
 I61e50081c686dfbcb684ae83ed3a53c6 <= 'h0;
 Iad3645f6fa7141133b12534c70efc80c <= 'h0;
 I62c110783203a19c372c6aeda18ee18d <= 'h0;
 Id7216252c1febf54691e626861f6215c <= 'h0;
 Ide229e0c521de0ffd39c67a6f078766d <= 'h0;
 Id25c2945168c44ec9f0a4bb2dc6aaf68 <= 'h0;
 I68a5c8b30e8d3e5b0d710c7f306304ec <= 'h0;
 I2b3c4fca6b0feb6fd829e9cbbe9d7142 <= 'h0;
 Ifec9e94824843f4cd8d623219278f87a <= 'h0;
 I7858226bb4feb944c5feaa52f2b51034 <= 'h0;
 I3b39fa7f2ad7920296a8e01cc9c12cd6 <= 'h0;
 I1201c86e1f6f9e890181790896c4afa4 <= 'h0;
 I8280be337ee3709b32502e07241156e3 <= 'h0;
 I3920223ae6d1a6d2ff327f53933ecad4 <= 'h0;
 Ica4ec266d79edda776095c95c3c20630 <= 'h0;
 Id23811d7cf32f6c5c63ce2782da15720 <= 'h0;
 I6df32fcf5553d3b899e6a67a35b852b5 <= 'h0;
 I7a01b2b85d70a35d44836e181a22b322 <= 'h0;
 Ib725193cf104f9b56c3211df12867643 <= 'h0;
 I45b1d972b2a5028cc340988f7c37f2e0 <= 'h0;
 I186a56ca3712df6983eb742d7d80a37e <= 'h0;
 I389856ba7ca6568e4ead3483c3e52353 <= 'h0;
 I66b39fb4c54ab32b2c876813544ff6bc <= 'h0;
 I591624fd56ff315e0084af5af206cf8e <= 'h0;
 I3994dd74d52d8957e443e869cbbf7184 <= 'h0;
 I92793401ab28d5ed265775c0d165dfe5 <= 'h0;
 Ic499c718cc4866eb8536d66ae4fae0e4 <= 'h0;
 I3c28bfe18fb1543683ae264c396a0207 <= 'h0;
 I083aca08b0d0bd2622d0f7b6b2aaeb99 <= 'h0;
 I2fd3c0dfd43b65e2fe8afd3368a50fc5 <= 'h0;
 I58332f7615e647e757033f6b643c21a4 <= 'h0;
 I22bbdf426df953feb5acede78c31b9b2 <= 'h0;
 Ia9f7a93a673c49ef3bfffd6fcadf845a <= 'h0;
 I687ab1878d38c7c988507163c8a60070 <= 'h0;
 I9efb470a3342962583f19eaec3a0ecd7 <= 'h0;
 Id7f7499e9b3f529781f4aba6e63490ac <= 'h0;
 I88e14285aa13b58457c58439ad1c8c87 <= 'h0;
 I730aeccac38e1622c684c468f8cb29f4 <= 'h0;
 I9427589efc5ae29474734dcc6e36ea81 <= 'h0;
 Iba910435a91ee873f76fa3ec9ac9c3d3 <= 'h0;
 Ia3c2d3cea56571481655cc77ee025558 <= 'h0;
 I99ba3451537a2876c9f585f72911bc4f <= 'h0;
end
else
begin
 I53846946a877f30f72076ee6f633a0e5 <= I0b93aca5ef7c84ffba0064eb4a53ec4f;
 I5d219e3294f2763bc17209a55758ab54 <= Id37ee8cb85e5cd05bbe92dd90fd22777;
 I6273ee09aacad20f733530af1a987ff3 <= I41450c30addcb3bb1d2c1c036dc26d2f;
 Ie0f63a67c0a6ec07e7bcb943e7804f9a <= I078a7802a3340b0c207a002a4046a4e3;
 I7b83ef4e45fe20e023e08aa3e56bb21e <= I5a33c28f0bc44840136790663423bd48;
 Ibc8f334cefc147e5c58e7542d26fbe2b <= I777e21d17f74d2fe893977e1654e2c2d;
 I662a566f576ee431bced6f852294713e <= I0b457f5bce1ac08077d7c061655dd03f;
 I2a4bc966b71864a79f582727f122ab60 <= I8d508a837624b899a748b9152f4a787d;
 I23d9f47edf51ff1c2a6275531a1f66be <= Ib226330c1225db758177402a9bcb4848;
 Id46ae2d16f43af3529d91eb4d6bd098e <= Ic9d6b4cdd3bfef73660bcd8319a9a7be;
 I51298122656d9b893c1dbb33a281f134 <= I8e094e0c0b13b04dee8f4f70fdee87c4;
 I22e0a22ed1768671dbe3caef8ac499cb <= I5469abe94b035be8eb8713d061774eb5;
 Ifb9327c663379f77471d460eced9c1b7 <= Ic6dd18ea6082a83222edb24cff9873da;
 Id6080749dda3cd29c1ce36ab39759709 <= If46aa2c29de75a5a44a4d629204b0963;
 I532fd8f9065e524727e276a1a8408008 <= I86f471de37f4d7f2599425d1f7ae60b9;
 I1f0b23c673ff55115f55c80a970172fc <= Id4063c01903ecbf60f39cc2a65c5b73e;
 I9f99ad4587fb6907b3804c11125f738f <= I1be4f732652b930e60cb6bf53fbb7132;
 I719bd7e94d4289c6fd59bb91ee559980 <= I64355c5e822a8d545c6fded925a984b6;
 I9103b57e3550cb68266ba8b102e50dfd <= I865085332575d46654188a23e78a5ab5;
 I89fca1c1832813b84cafe145377d7b5e <= I5a3af3b67e01e19177daaa19b995b876;
 Ie17de6e388779502a143212813a50317 <= Ic82f2a7d5019f0912c100d6336dfb3a8;
 Ifcc046128364b8da7bc3d9ddab96a061 <= Icaa4f34ed9aaa9f1690a03ff7c374de4;
 Iabe4b7a23f682ed62162dfde9e15d6cf <= I7662e29bd142424284880f29b6d32038;
 I734eaef0b7d7f6ae5d668ac9b374ff51 <= Ib9befe6fabe9ca87ddb96713b6c6e0d4;
 I0e0e9fdfeb3e2115deb903b973217384 <= I69bd49e2f242a3c2a32d182a32cf39f8;
 Ibfd2fd7aa2426054706d0c4e4c0a7cba <= I820044a9516905bcd63a9e6d98ec961d;
 I0906247e3ba96971232bc42185c9a9b8 <= I4b1cce4cb416fc1776b09254d2589bfe;
 Ia3908fda391d7caf1b479d9655164c30 <= I9cae305381503e9d92a4a8240bb2aac0;
 I820e95cdc583108195e8dd0e2d1f4b7f <= I5a1301cdc00c141cd57b0c4b90d7dd7a;
 Ibdf5c2c57269da1b04748a59802c8e2a <= I98abd404eafd5efdc2a990f2760fb0d9;
 Idd85c8c853438679d99bed4d0ba46af7 <= I3e8a5169cec2e8120a2ba6b6dc0f5742;
 I4d617d0b669b3ff1b08dcd4b7440af33 <= I8b50f6cf167c2ec62d739f294512c324;
 I60d579b60b02f9fc14e98d7d0eb54c18 <= Ib0fffb83f9af51787fff93443dd10287;
 Ic1a37750fc3d7eb08ad649de157f45a9 <= I3e4d4fb93b28d431849e2dd307f91197;
 I0c13ec63e7208b35a1d4511e1da29fa3 <= I85b43efcd6de020aceb66ed5948fd901;
 If10c9545a713996735934c5f15cf5365 <= Ibf4c9739576bfc4c8d79dcdbdb629a6d;
 Ic475963164a956dd24ede91e9d61003d <= Ib96063e5603755f2354a15d573374fe0;
 I42001c4b6ab9fb03489ca25defb6c222 <= I5f07fe122c1bb26c6805a7f9d31218db;
 Idcfb16adf2996c8cb51e402daafd1734 <= I0ed871a78ca4e2815ce45133571353a1;
 I924108a2723afd07735574a6f4ebe671 <= Ib0ba4dc6303dade812ab25816938899e;
 If9fd9ae380997e75ebed2ddd3f93e76f <= Iea7ffe40a13deb5bfe2903c2965e4b63;
 Ief876b7b2af1fbed4d3f457cdb46e0d9 <= Iad7d1d253ed65347182adf53486dc1de;
 Id2bd196ca25e1a077fb2a9207f143c01 <= Ie4cc734fa69e1b46577b5df885ba3592;
 I926e2a038d48db29b5ce215cd6cf6a04 <= I75554ec87598151940cd118e6ee59741;
 I4ba2cfd94590dee1723ce63afd0926ab <= Ifec751297668f80d860a9d6cc176e5f8;
 I0d42326464ae4c3a55038e0343cebf5a <= I8fcbbdfd901920672268b4d6ca269849;
 If05fde321fd1456422550f5c3903b826 <= Id16656f72b76591b0bd03a3c2750684c;
 I41ec48a5a1d657a6266b8f845550d0c2 <= Iefa235bdb6e83afe1f793787d8dfca2f;
 I76473b4885d423029324fe74ed13d6ed <= Id4fc19c089fa63c1b901fb64c9c0e064;
 I8ef2366947e3f1352f3874e4ac58d7b2 <= Ib22f4bce6db16f279ad4085901174664;
 I874c1e455f85e617a5032ec230fdfdc5 <= I432b06e788f0047c5e66cac253186eca;
 I16d6b6b19890a6bbdf15ddc27717aa30 <= I51d270bbc6e26272e0d6998307c33272;
 I6af6d04126eec9eb91e5653cc95c9ef3 <= I7f0c42c0c3c63ba11cdd3c26093bc3f5;
 If501a668f24fd62a69d0e3c253739c79 <= Ibe2e871186cde032e6ce4de65c0fbf75;
 I9b70e215a2a1578811b40c669826d41a <= I9aaab4112c129c0563c8983c3cb372ba;
 I26d82966efbe51e03edcd66a5a507ebb <= I58b6cde8739d1e98ccbdd13b1a963c8f;
 I2e4afb94e4af76b4e3d859815bb338fb <= I6d3d948976b4f578039a6dbaa8f08642;
 Ie19faf5d037b74974102c386a13f4946 <= I714b8ce615cf088e1ac52a7e22eb69df;
 I2d56338af0755ae5c4ef71ddad3112b1 <= I7672fb8749f7573c27144fffd1721ef7;
 I99ab212db901b0e65eb33be27c46bd19 <= I5fa7ef4e8130409885342236b9f60fcd;
 If8c09c14d78b1deaf76df6f4de910c64 <= I2ab7e691bb0a2f89f9cdbfbad80d7120;
 I1b0ccac0f5cc741403fd6e680899f96f <= Idc22eb4529d6e2f82fd6c23a113809da;
 I38153cd88e8b2452977d7dc9b9f44a74 <= I449ee1a89494568e104c9e29f66d4262;
 Ic32064fc62eb1cdcdf416a6fe78becfd <= I5e8f226f92643e61ad527be4f148de00;
 Ic10eb104fe38a176a51507e748406958 <= I56a2b51825ae20cd1d9b434aa976b4dd;
 I979fd1b01c99b76a4ff2d0abfb0c2ae9 <= I580e0ae47b151812c4373cb1f268e4fe;
 Ibe530a86c501fbc8dba64ed24806bdf4 <= I69e6eeed488ce445421bf458f3d1baaf;
 If03531315c68272f7de2b0e969770f48 <= Ie3781ac0023a6e8091d66990ee3983ff;
 I20160f4e380b0920bcb30a0321b7bfa8 <= Ia6a4c1e9dcb6ab1ad0114e2da7a396bc;
 I2bbbe5d3a72af5f654976a7fde2d2d16 <= I91ed400a23a8aa771dbb930317b63466;
 I70f4396800d2cb065ad5fe655bacbfd0 <= I15c7e1315b03dc87984424245b7e6dab;
 If27a0187d1188cf7a8aba100a90cb069 <= I4ae2e6ccef3d457713203f83eb10d60d;
 I8994866d080b1befe414fea347e7e74a <= I08a273aa764a26045fd205007493d27a;
 Iab6971c846299eec0a5cc93ad10e569c <= Ifae99596becf8c2c7b69fc3e508a362a;
 I8730924fec54ffaa78a0ffea7e8386ba <= Ib080cdead060a391cb67c54d97c7fb0b;
 I338fb9183219691c6b50e6a824fcb14c <= Ie14db629163bf8c01b457b0df3bbb634;
 I1a3d82eaf2fc9235163c0a50765f4ef5 <= Ib4c7a688661be990227b9902dcaa0721;
 I922539f8d9ffc119ed3a5c92a21f149e <= I4b33852fd89354d5eeaaf75dcb84e726;
 I3bc0f1eaad327d5990adb826e54c6d2f <= I982d1672a39f86bf7da5bb7844bd57f9;
 I3009d4cc0371f83e6bec8fb38ae461bd <= I29949584d0bbd464970883cc5724f8a4;
 I2e0ae02d7a3cdfa36e8645cc7dd0bce6 <= I03ec49385def83a3f577d847012976fc;
 If2c59f326f3658dee0fd3b048af14cb7 <= I6bb12bbec43b6315c92ac22f43ef5a60;
 I04431bd4be4601d3cb700c0cd6d9fd24 <= I5c49372712967408ed819ba89624dc98;
 I7a6fe8c804087a19e32e760f50e3edfa <= I477fb86a2ad5f7ed4f225b0c85609bee;
 I979817e250e46dcc05f8a6690c2380f9 <= I67099935c6636fc80d472f193753ba55;
 I3bbb836eee6b5e10fe55879f8620b888 <= Icf692082f362b6bb08f320e2b27853c7;
 I8bc5128382cbffa289caec56f9b4a3f3 <= Iae5385d0436fb1f5c949c0d1e8c3aa96;
 Iee4dafc9d42609fae74410897f29a78d <= I6951d4063e974375523406edae080570;
 I4ea5b39ed827d8d4618bcfd9283dfa83 <= I54e637eae832d289eeba34eda853a657;
 I19aa6440394778642eb50f3b94098ea3 <= I89479946789730c4000d8166356cb964;
 I0653a9ef861e5d8af22d120172c2dc03 <= Ide9c460b12322a14105bd0484d4b9135;
 Ie0aafaeee1abf6d27a70535385ab88b5 <= Icb6633d32c69b880dea230dbae0896cd;
 I1583cdcd13120f953691a5a60ee72b11 <= Icc91b46df090bdc04306996433be6136;
 I8080b45a37a3de79ccb338f353f19529 <= I5ac7c7696f008ebbaf6019fa5ad57302;
 I9bd98a9d18ce7c07e85287f6b80bfd31 <= Iab7f04bf5075b64439bff52f4779ca67;
 Ife85d240c60084dce9b3d7cd87060727 <= I9c3e9f415a26edb9fedf25288a8fa453;
 I11f2e4eafc706b43c10a26edc8567052 <= If0e39a30beb041d9c6b3c168e965a1af;
 Iad3a9febf269d9607eedf29912b04af9 <= Ibb59c086a89025918626f18799e73605;
 I75705fa2cc0ac0577570501510e4e0fc <= Ic436ebe8aa48c3e6e935f6ce0b3f43d5;
 I7674ab7538766e842366dd08ddbbcb28 <= I05239dbfe2cd2ef57477ecb654880bf4;
 I8cefcac1f7fa2df45bb8a2f3d64f99c3 <= I1765216a10c88b6081f34198e8a5d26f;
 I5fd378ba266fd930a839cad56e500ef4 <= I37b9f75cb896a9e45a650b6dadd0b2ff;
 I71a33ca1c7d18d5089d08a8476c8baf7 <= Ib9eeab393231e41cca081394b036bde6;
 Ic85b012b9fa77becd419cac0f3692aed <= I499fb85792bd0c5a73022ac96ac27f13;
 I0ae9b4ca5ebb5f3d2e8b02884069e4e7 <= I3da1d9759bbad87b216b2bc8afc19f8e;
 Ief312304eec0415d1ab208ed6726dd12 <= Ie220bafbf40ee68b7591948b607fcaa0;
 Icb9ebf1f5becaede273da59f466506ac <= I34b7451c43eee381ab7b3f1e2a816b99;
 I465b9607a8dad0f1c499318d04f42aea <= I5a3b2767a2c2b41984b6f2a7f05dfcbc;
 I2523c109974807b3b1c0f4b34693e255 <= I8ad73072ca340501c2b14404b9353b08;
 Ib4e3121afd90b877b94c4c7cd29e9334 <= Id3987a88bcc92458973c9ee529f52a56;
 Ibfb66b89c59008f3d4497ee16dad6712 <= I49666607354671cb5d6ec9c3e6354f42;
 I2d042c4ef15b2f3bdebbc7cbd6c00a1f <= I4da0ec3a6c662f7e76bd3f6c43b40722;
 I489d1b46970800e9684c68b439c15be1 <= I039f5eff8e87d37a9cf7d754a82df849;
 I835143e23243f3fd25cc1ab0ba5c123a <= Ia6fa92e40471f5741d59b8515c67c24b;
 I028ef05ea84be3bc45c518f4f45653d2 <= Ib4ce242cd8f88c4eb147129be5e6785c;
 Ia5a39eeda95dfdb2ab8b55ea9f8b62c5 <= Icc28fa9f2f20d09b439a9553b6e592fa;
 If5a85945ad1f8d9bdc9213c5ae2c890f <= I8b4b437c18f15ae386e0c12371151913;
 I6011a5fc7b168a28fc9a45f796629b59 <= I7c34ca74407090b532ec5f0f65e5dc74;
 Ie703b5f1eeedaaaddf56ded14b1765bc <= I1f69904e43d7fb93f39873efcbbb558b;
 I21f34fbc269f5424ea30334ff7ab54f5 <= Ie1f3985459b6de4b08d14263f5b1aa18;
 I07b47fce56edeb30319038e3a093efd7 <= I3640c422ee8389926afc8108564b593b;
 I24e7e5c391285f28c20f74820a05b552 <= Ie11fa9bb26231d41be8646707525d022;
 Iee1b23b99f7de56829706633297a0513 <= Ibabb39952458fdb3127ed17f3909e043;
 Ib4b61d3293900c38e8aa7df0a617b476 <= I8b1452ad1732c78b5397caddc0d43daa;
 Ifd5fcb1552fb372ae203fd0166d3df2c <= I5adc876cca35af9714a2cb9ca0eb3ae1;
 Ibb2fb63aef1d336dfa829cd5ab3675b7 <= Ia2848a15587c0e23eef1de69c2a238b1;
 I1672371cf33b259cf87210cc49aa35c8 <= Ic4119a74d5a813a98baede5515be91bc;
 Ia34735ee7f7ca164c2ae71980060f56b <= Id3b3231272ef7b602acb9b7dcd5033e8;
 I2372d0a72998f0630e994aa3e1c20ff4 <= I05e604f9ffc573b44538d9d864dd4e92;
 I8e363e0bd65cae9725cdd70e46778fee <= I116d21ad2753927dbf389f373bb1a344;
 Id6af962a16ff79ac6e9da3b4518b80b2 <= I3805a70a8e257eeea2bdc179fba1d185;
 I7fc8c9245183d05370746c9b2fdabd0f <= Ie2d31cc4673f92faf8545984e9b52031;
 I693f2c9a5d4da90c3105876991c4f4ba <= I5bbb1e57ed53613e06ba3fe1cc4fd266;
 Id6c07cd1f9f428b0d971639939b9eb8e <= Ic4e117cdda2e62382412fb1dfb9c850d;
 Id6561e53aa8f9fd116159969afaa20ae <= Iab33d8521b7118693333cb5f624f3904;
 I8267af03225d6d1155142645ad7f53a8 <= I4183bbdffed2418b9190d610ef9c85a5;
 I567872d8892064b62caeb3dcdc39e89c <= Ibee805f0c9d18428759c5ce6c61f4dee;
 I5072b405191b837596b5efe4ec159519 <= Ic8255e62414174e60282be5b4d63c494;
 Ia4e5d30bc160c1f72c8f39cdcd13e5a4 <= Ie76911ee442cfab80022b3a534438350;
 Ic46dd8ff5a79971f7c22f4be0f1f4b23 <= Ie9d09a2059dea91a80a00bdeb56940f2;
 Ifdd13523ba0ce3329e3aca49a0a36385 <= I86ecfe340941ed77c09fd4c69f5c272a;
 Ib449b5d80a7f5a1c5d0d3784d8f236b6 <= I511c8519304a31c10313838c1a053f85;
 I134d223e71b68cc9c76379f1368fb0f1 <= I8824abf0eb1a4d6b48a26abae23d0bff;
 Ifa82272c492ce1ed4b223c0cb2b135e1 <= I5d8953fa34cb14027d8375d02999f132;
 Ie501d0f392be1309df48c1616ace5a27 <= I0d8e31fd51ec5b82c5206c307e0d53f7;
 I29468f8318cd5bebb5cea27e1ee57b7f <= Ie1ea3318d114c790e9343e45555755ab;
 Ie3f06a529d5f22198b3b33d649b740e1 <= I495a91d95803df2b5cfca5053bf13a9b;
 I6740505fac3e83de4a6525ac9cf489d1 <= Ide9b85fb8d57bdfbf9b8de9c18e9c5cd;
 I0456541b6e82ffeb05fc4052fafc41f7 <= I9cd4f5d3b10c25759e7993f9292a7390;
 I6d5739cf589ed46b6f57075a3b2a974d <= I5ea9ea2fd34572dc6833ccf368e52ccb;
 Iabe05603679da24a44565e756adc0881 <= If3883c5646540cf78aee0589c3cd3022;
 Icaed4c0a915898eea654ab6f93973ff3 <= I61df05bea32eda79ed88930bbc84a13f;
 I98805e117c2f4ba4a8f6c2755ebe1fee <= I7f1a2ad313f7af4a0f9eb4311f35ac12;
 I766076681dc49b817ec9302eae86d64b <= I685601482e2bded73351f69f3f5c21b2;
 Ia82b6e01034a63c2a1a446029f58f1c6 <= I484b91ff2256c38308e18bc50afed4ef;
 I05de7fd67a0e226201b563fa6c50f362 <= Id86467d5f10985a00ab65a8b029a8c82;
 I8df8f128712fe5445a97566f8f29ecd4 <= I56110e27931a312345e239eaf42781a2;
 Iae9103582be213e81ea0a25e5d49004f <= Iee57da8134718b73f0598a1884ecf424;
 Ibcab213dbb173403005b3d65f780fa2d <= I7de0f163ab38efee6f9c2f362708f4a0;
 Ic59b57cadd4b8cbe63f996111e9211b1 <= Id397e815fb86c38fbb509692ec4dab0b;
 Ide1a993a1dfca37107fc81e985714d93 <= I2c5e75d48e9ca1a198d70980900bdc41;
 I7004a1bc0ec2272163d33907d21616ea <= If728db81c67f83aab133c8ceaa3a5c7b;
 I4ac93ed29241fee9390fd824452e6632 <= I80d54bec914a5b89de0f5296459b152d;
 Id6bb9f52fa37334787904652fbb1bd95 <= Ic99c4503bcbcad1099d0c26d3d9161b9;
 I21281177f31dc70c65db2e9a3aa72392 <= I36119b67ff8b6471d47a6681ce27666b;
 Ia64ddbc7428ff56489b0855ff0fc67a2 <= I29103484cf42c813700bcc89a04146c8;
 I4cebb1a21b9c76387237fe8784f97ac1 <= I3cef2dada2657f2140d9bdc43f83057b;
 I3b8cbc445627a75cc4b05aafc8a23cc5 <= I23abb9c83aae42b4b3a330f277ce3c5a;
 I46c35e4856fb0288a23d9c4c68290ee9 <= I79b6e7abe2503f1f13195584805dfcb6;
 I4660e4e54643b4a73afeecea4a4284d5 <= I4d042a3d0026d6b93b5b394034174b00;
 I86454d943e7ff4b244882b0f6955d9df <= I92d347131e209dc81a8321d27d38a69e;
 I3e0245e2c18af49b10a4f2ee38ccdd20 <= I79c6fd3ceb89abc93f49a67d913505ae;
 Id34d6ac40408151f201a8b3131463b3b <= Ieb5038840ac4ab2ebdd9cf6222c15750;
 Ib002905f7b54145ae3dcf7e0f8715b8b <= Id81b8442322f6bdc3728f5459a830aeb;
 I3ffe132daa39f108095cd1fd5c38c6d6 <= Ie3a852b81ccaf2d520d024dd989caa47;
 Ia057defdefe85e4b01cb1acf025fff51 <= I33b0bd948bf4495908c59c2d8f58cf2c;
 I080d693c8cdddee8f9c80ad68d1db1fe <= I09a19721c1644f9d1a6eaab84d8dddbe;
 I55f1644f9601b3553040f8b8ecd84eff <= I7065b10d4533cd967733d262d5e5777e;
 I30ce714aeca130dc1978c6eda3ec0e11 <= Ie75d8156129eb98d76783e3a6ade280e;
 I4ebdb0445ef12223edf4ccf0e4785b01 <= Id3d25ba968ed699bd0b61ee32695edee;
 Icd76d18cf8b38caaafc592047ff3b48c <= Ic560d519645177df445db05bad34e60e;
 I51195d2f4e3b638d1f1d226ccf89ccc6 <= Ia5720f57dcae8ac0b00ac4e4a3c89657;
 Ia29e3ba7f03b070d4381093dcafcdeb9 <= I8cfcf912f60acfc715c63291a8c04729;
 I2c9a9e255b7ac39f5d6509cdf27f6d4e <= I6e5f2896cda9b8db3638d2b14cd6ac00;
 I49dd3ecb280e2ea8639a2397343f1700 <= I349da988b53307693f1e74a98fa686b6;
 Ia1d516cb29b48f621e47ce669cb9220d <= I47ec23a2e834f9c66f23f1e89eaf8679;
 Iecf3c7051c364595cb29b47e8ceae9d7 <= If03782abea72e6519c530636040d2291;
 I72fb085a491b61f89d4f95cda02b4b3c <= I512ac9f87b0fc7590f5434fc1e3f0372;
 I1623b3a676440bab948f5f01c31c87a2 <= Ia0d98d1391069c78a92be189e60cec14;
 Ie83ef8c66f723e3ef386055c5d0b9d8c <= Ic75a566d180368ca17dac6f967fe397d;
 I858523451a6554f7bc0238638450bb3d <= Id9acaf5c4d2e0ff41de104ab47e77756;
 I82c65f5d9ca29f356382cf62e638f3a8 <= Ic0a4f0637df63f87635fa78c21b2e99e;
 I88222b3d351f2f7334c9f3f22d3f0255 <= I4a61d91e170ec3b767be88ccb343f1ca;
 Ide7e980d6331b40896f26f3377d80c32 <= I12a049b431155546b8663137cc66bb9a;
 I2347ec4791ee62d976d13c7c6319e16a <= Ia019f222e96881e643709af1eb85011a;
 Ia5706e1260d5d1b3c625f58c1c2fe509 <= I09be79fb5efca2f460b667770755191b;
 I4c48730b147596406983412e0e6ae556 <= I53f09f16c58b346a02997b021f882363;
 I7de06231997b971a3acdfe69ebd5a394 <= I19b06a7f2c499994044c7dae5057d8a1;
 I70281a4f7bfe2fc5e4a0b91b4194d286 <= Idb57cc9ee60ae36bf3c0117776a46d70;
 Ib95d1aa238c37881c0934c8d22cc79d0 <= I8c056925751f5cbfd61b1195817d25b1;
 Ib9d8fdfe03633433eab48b80f9d4bae8 <= I8b92da1d7f30fa71249623b2bc87b462;
 Ibff1757b162a6cba3637e2a0c53d4f57 <= I020b3d3e1109655d6f795fd1ecc0a322;
 I69f8f0b916f8d0b4d146e839c19a0756 <= If0e90362af64ee2a20b44f61aa766fb4;
 I0f58fb5960dd9007acf9103e1ef428c0 <= Ie192f4f4088d17d1f7840213009ca3be;
 Ic31af45750c67aca08c2af5f1fdc52d4 <= Ic72e05f3be735d52d9354cb8f43c1cc0;
 I81b800210ac62493bcb6993bf20de4f4 <= I76141646fbd2efad1e121c6e08ac174e;
 Idec985d498536ef129885e9baaa69be5 <= I4ac4e1dec3801e462a47f80276b42397;
 Ib85fdca5ff6cd6fd13a196d1fb380166 <= Ifefb5a209dde348266eb66805c0a7d2e;
 I64c48585300f968447198fd11396fd71 <= I92c5b8b76f0000bfffa0120f70f1991a;
 I9cef63d7e32492a449474355630e84b2 <= Ia94fc30c06efdb8ae6f388149d0dad5c;
 I8d49cc394888a3e49b8e5cd72f2877e5 <= Ifdb73b22fe15d17de645cf8aa3da99e2;
 I19030461146fca1f78cdda6d38cd91f1 <= I0b0e5a5734bd09dfad80a75fca5a763c;
 I80802c2f239fbc3ed9bff61e9c873550 <= I73354f6673afdd64f94fe36e146cace0;
 Idb96776120ec0d249a660e1cdfbf4362 <= Ibe0a9cbd6da728e5f7e53081af472ea9;
 Ib8b1376de13c22be5126d585890438d7 <= I0edeae6c95ab6198047ded7f3b41efee;
 I0a617772f4b574bc44555b85eb425b3a <= I473cf664c81394c8dab1d7f145b3804b;
 I3a9c038e7e278e6630b3defab662e10c <= I7201b831890988766bc871eb0fa6e19d;
 Ib741e42703c8b7e4ffa9a6fe599e78ec <= Ic772d12c6a9f51ff6cb51bf7d54d1b21;
 I878e4888b177aa7880c8ab11384db32a <= I16120aeff10370316421751a8f4e9505;
 I294424e35f618c68248a468bad92814d <= I77146070f8693370d971ec3a91e18f84;
 If808ebd32478faac57b26b5306292dc4 <= I784fb1f69095ccb95c4bb705539970d8;
 I122612ac7be83ca897e3d0212c7dcaa1 <= I2b2174ba9f0956782a3ab584fd11777a;
 I88320212337ea2d63720b17e98675475 <= I8f31a3afb2cc62773332f251278c1153;
 I777989034e3f2e68b036801349f439ee <= Ib2cdf1583fe14fd7b16229572511fd7c;
 I20f9fe0be090aee8bf1dcc46f806d73c <= Ib04043dbfa7a17abbb728899e2459398;
 Ie26a8b21d119555a1e9e6b3c41606658 <= Ib1eaa856a32de8ec5107bb40c8611700;
 I47c779e7352c5c5f13cccdd737dc994b <= I04ac748d74a312f05ede4d4665042de6;
 I29f7d07e6ad56f0d6a9b9126d5ebd6bf <= I70ef81ae751a5a7640ce2d4b0ac381c7;
 I7ae4796f21cd658ec17c8ff97f369784 <= I6c64c351f3b91838c0c3c25f3b06d201;
 Icae58f7ba349c64263a4465f8de68bd5 <= I146352e56b780e8cc0f10ac09cee3a2d;
 Idc1a3fedeccab7f0ee34f79366f5c4e5 <= I966ffe439dac9390e18e84a65e4b6f11;
 Ie8117cdb093d8606a07c83ee8e80b388 <= Ief16bdfba3e4ab746af015310ebbb6b8;
 I0a65eb60e084d42aa5f5d9d6803068df <= I0bb8923bb50a4fc7278094a514c79fb6;
 I7f0634ff89c088ca73363e951657ec5a <= I9e93a476f9669fb72f7999a6f0a05c16;
 Ia45d63e797413cb23c429c7d7a1eef02 <= I0442bb2973db673118791e504be846e4;
 Ib7b0721390dec3041d5257d0e3df97c3 <= Ib00b860d9b3981465aa3bb1f18cfc627;
 Ib89de4c510d53bd06fe0f10c7513de04 <= I6ddab9f5aca020985482b76c25f2f81e;
 I2938e6df94b490c2100ed57268545d36 <= Idaa6aa87b597a3bcc6275f5f40444057;
 I8b7353fd85fd2ee67a1df24a9f239f50 <= I1e2ca5efd6735a6e241f9bcade3c2b60;
 I66ee7fb42c8ba5991ac6aa8cdb51bf52 <= I50da8ce0a49993e0b7c16710e68da821;
 I3ceb68a7f17d021fb3ce01821a19e7d8 <= Ief43e8dc88393e5a4015033c4021a8e5;
 I649e640596807ec607a1c29006987d98 <= Idc4a8277aa0ac4ac35b9fa6b37f198f9;
 Ia67f20bc0f3e32bf1e443bae34efc4b0 <= I4f555c0f5b4b6f79ad394e0f196c8e9f;
 Ib1af7cd6a6d84431253d818fadb177e4 <= I7ddabcd95dfd2719f9e9925598e0cd80;
 I6631364f87a3c0d43c4e1e433b61a132 <= I007d2500c173825191e1243fc0758203;
 I8daa733c7e34401a9002dbeef55b89f1 <= Icee24ae7d32c16a6b5dd7089f6a63d18;
 Ief1269d4009e33d56efce8d693d3588c <= I0d5ad201c17a461d16a13675a0abf874;
 I9274d5ddfd1bbfe08138024e1eb81052 <= I8cdcb20840d2cafe54bf1a40bb5fdb1c;
 If36edf1833e16bf79b7ea16dcc551d2d <= I5dce978811c8a3680684eb168992afe7;
 If978d531c028e4c3c00cec8d057703c8 <= Ied4802a1ff9e40f97bd6ed7e5c9af351;
 I1cc0a80d74fe4b030cd838bd32b3cb20 <= I54c34254efd813baebdff01bb5d9100a;
 I0de61810af282ac4baace4ddca69f88c <= Idf998c5802562dd8ba5cbbe2d8f4eca3;
 I4566be9ae01ab539195295433536bb4e <= I5140c93c2312dc879b408cce4db484d3;
 I9ba42ab3f14a648fa7ba73189a272474 <= I0110a5e1c6faa19f5d97ee4b4f763285;
 I735b9bdb73b8701ec3181c5c08f9637c <= I923c20fa85b752d9f31a3476e863c4c5;
 Id88f6239fc5367bf8ce4c1c3bd45f75e <= I0eb29e587012701bb6ff57aa27d71ecc;
 I78d31cfda6c9de83fbee1581d2cf4330 <= Ib3668e1656878dd9ba2862b988011686;
 I64ccbe69fe3724b0b97ffc27c7682b0f <= Id7a758f960bb811f4ebb46662228c33c;
 Ie29fc0c82ccfe2e936226bbf8a22aa93 <= I271fa5cfca7bbdafb091c3afcc3a7a41;
 I9b5a96b0522eb62830257171c98627a0 <= I864329472b61fb8580558865bcee6de1;
 I3b383604747befb7811e7cbda19108f2 <= I78527503b3be9fca973ab9fb7f987f27;
 If0b2cc476e6faede63243dc637ef5233 <= I3f50edcfbffa653e39523fb6125d4fd5;
 I6e38e23fc4b5a6d9f5990d7f82f6a0c7 <= Ib5dd6975eedeed971f4aeaef77f28f1e;
 I0730fb0081845ad1ff057ca56b951d75 <= Ica77a9f6eb020b850ed2fa38021f33fe;
 Id5737f058ffd0a11b2d29f088cf7591b <= I783f912ad4fff3731add8abca943629c;
 Ie41e239efec92527dd0d50dbc4dae735 <= I1d7c0387f65da7d2ae51250edfc764de;
 Ib906993ed1101ad0992f24c4dae29370 <= I809a5efeed0db403579d08d520c2c9f1;
 Ia9eb0f66bc38056887e1492ee688f373 <= I7649e3988149218a8845000ffe68477f;
 I4c6811b2d28239598a23f790a03326fc <= Iad53806231a0e21d8b1e6b8a22fe3dfb;
 I29271f07d1108d2c542b60c4296c7195 <= I9dcd325f9d12b6495d5b9f050af3c72e;
 I9ac5de9728a0349bdb44341a68adeeec <= Ib0d29b4d3693a1487dd507cd4610006f;
 I3ea1e03eb78be51505b0bdd005aa6e2b <= Ide3d8fa67f76ce3a1762381698b59301;
 I969fc047ddc46bca31190e0d7f435bd9 <= I85818659b37457732130fef9b829758e;
 I7a23ad071ca3404684d12d2a0f36483d <= Ia8d5826890b3ca20e13dfa917300631b;
 I38083dfdf321de81daef5771d0546525 <= I6b7c6fa01374134b230ebe6de1602785;
 I894d1f8f86188aea7fea540ac74bd39b <= I4ebeea8273995c7ccb406a5cfedc3ef8;
 I9d6d3cf2eccd6cba144db2459967a901 <= I6521570d5f202bce800b1c49adf3f2ca;
 I8cec6c5d567ae4efab02118383cbb0cb <= Iec61267ecdecf9fe305142fe095a21bb;
 I1cbd09f17301a0bee1cd695a2bde4e1c <= Idd383af878d242f7be34d1c9d3efa0e8;
 Ie767f5975b691400b250054bcf08867a <= I44107557054891b33135a13058e00649;
 I54b29fec4a88bc1e03197a0c55b875db <= I013496291a38e851842de8ea28b540ba;
 Ib0c39d1e2cffc0326a30bfd0733075a7 <= I54e8b21c865654527ee0720a72ef1cd0;
 Ib4dee5c8efd8022bd9c3f9bf8d5e328b <= Ia40d6a1517b7b0a79c88646d209263dc;
 Iae316011740707036b166a712b32f2e2 <= I1e10e22806a41d12b8c6328dbd9471df;
 I3ae123c41c91d9b53a70aa3e4793be9b <= If96824bc7f67bd2bce941ce96559867e;
 If4ccd39857a7317488e9215271db7210 <= Ib252f7e32a3780abfb1a3e9285d0ed56;
 Ief6d7060558cf2ccd8d561ec17b846d5 <= I192fd55ca87b7cb2277aca900d015b04;
 I2a5d6b55814dbead5a30d961f8f7b478 <= Ie973db372fd3127653d6c63a551a8c0c;
 Ie03342fcc484bd9f1c934e675c9f6ec4 <= I3446695b823b258ade0a7ac2aa9d61d7;
 I195e5182b2d3136ff3ef4572cb4b88da <= Iea584b5174273f9082695eec0d7a8ab1;
 Idb2832cb2e894a8c02e7dab1dccdef87 <= I6d7f0d64776ea582e326ca3b008f2b35;
 I5462aaf13ac6e9761929c998fff0b87a <= Ifc32a10a9fcddca15eeef7d093d1401a;
 I8f9db21a5dea66f9865796d164f689ea <= I84db677284b3e4bf9feddc2af30e9ad3;
 I31949043c0e635f71f9785c21d713c96 <= Ia04c9bc6fc469c62a3645e0e691b3897;
 I2135e15ed882d1293741fd593369f88d <= Ib7457f82785a56cbcb5be6c0432641b7;
 I8cfec980374c11bdc4947a8c69a55728 <= I42a4d0da5f0b890624310c94b32f1a27;
 I5e298171856ae5526301f6d5084f2796 <= I08a589b0a34d88ac456d6cf40da0f5ae;
 Ifc2714ac9c0b998653c2a1b5e9199d5d <= I2f1e3460880499c961fcb244ca935f3b;
 I1b7e4002a74d5f33e7d0168ed06aaa2d <= Ie7f199c3586f87a1cdba687bd880497e;
 Ib868c2b4eb4dd68231ed56d937dd4804 <= Ia3518f4b7c1b0aa2a864d5ce53158ce8;
 Ibe26ea03448b95798236cf228817dfd0 <= Id2616c8625d0a75ea0946506034955ca;
 I4ebe3a4a45add9d58508c58a27a5d46d <= Ic3c6cbf9171a81f229a0fb9efd57b000;
 I21d9dac9d09da39f435c7082dca90127 <= If63bcb026b347506aff08fda75ac7c43;
 I69e220ebbcd0c48f5cb1cf16fc33fa57 <= Ia79c0c66c81e60806fe3df0addd5608d;
 I8546eab32336885c49882f192be9904c <= I0695fe1981c8019decb9873e186934ae;
 Id4da583323a66a1333d836c5f7bba069 <= Ic334a0e64e305848782becce03c85d2b;
 I8c50bd38d4339a6ae19e13db1a1994e9 <= If737be717332ee2670d2c6736d9e0a2f;
 Ia19b6c2a9b73f96a351eca1700079c42 <= I66316458bfbdf6b24cdc0cd7396c84f6;
 Ia98d1ff0d0dac6a253cf48ab85e0eb75 <= Ib23a5c11d42408a0f4a6d314a670da51;
 Ie63e6f9d56e6b192f0703cff4813499d <= I792738baad12910007da8123fa0ac415;
 I0b963cc516bb0de18221dd724864d795 <= I64f43975f3065e3c7cfed15d5dbc8d72;
 If1ede61a06a91d3ae1874816901896de <= I4c0a3a24dcfac4edcdf29847761a8fb8;
 I7f856b89e8b206458e96335076d80c69 <= I65fa0e67f8ee4669bba74ece0c565a0d;
 I8cb21da337ae4059685b273b50116a0d <= I6bea44d0467b461aa22c3ddcb1d8f886;
 I72569b57d65e91bcea79d0682c51c4a7 <= I582cb5f8b17099f479f297c5475542c1;
 I61e50081c686dfbcb684ae83ed3a53c6 <= I6cba6eca48f199379e62726b4ac271f8;
 Iad3645f6fa7141133b12534c70efc80c <= I57cfe42eafe8357ec85906472dec3f36;
 I62c110783203a19c372c6aeda18ee18d <= Iec7bf02aeaa8630497275c7eccab7667;
 Id7216252c1febf54691e626861f6215c <= I388c7af9494f4c425621d3abfdf72b63;
 Ide229e0c521de0ffd39c67a6f078766d <= I2622bb3685a7d6a297506eac3efb9c08;
 Id25c2945168c44ec9f0a4bb2dc6aaf68 <= If025bad83549d872a3fc9c44248174c8;
 I68a5c8b30e8d3e5b0d710c7f306304ec <= I3440574538a5d7dd250fbc98d574548b;
 I2b3c4fca6b0feb6fd829e9cbbe9d7142 <= Ibe30f2ceb078297737ce1444c1e6c524;
 Ifec9e94824843f4cd8d623219278f87a <= Ifbd6f1ac3bb594aad652d4e3cac018e1;
 I7858226bb4feb944c5feaa52f2b51034 <= Ie41d26b8a9ac93a09ece53b2af8c855e;
 I3b39fa7f2ad7920296a8e01cc9c12cd6 <= I497c3961e446544a8031e8013ca80ad5;
 I1201c86e1f6f9e890181790896c4afa4 <= I6ab9d8eb7b8e3454b01a8e67a410624c;
 I8280be337ee3709b32502e07241156e3 <= Icd351f2625b163cee904fa4e446d0cc4;
 I3920223ae6d1a6d2ff327f53933ecad4 <= I79c9be2982685762d0907583f9f459e2;
 Ica4ec266d79edda776095c95c3c20630 <= Idc20427e979f3d5c03d7dd947cb4df84;
 Id23811d7cf32f6c5c63ce2782da15720 <= Ie8abbb597c8132b8e23936a5bc035041;
 I6df32fcf5553d3b899e6a67a35b852b5 <= I42b0c89a558950f658440d8f9916b42f;
 I7a01b2b85d70a35d44836e181a22b322 <= I5a4d5a128b1fedabfdc39cb019359106;
 Ib725193cf104f9b56c3211df12867643 <= I8227a9907c39647a4cef8e883d487913;
 I45b1d972b2a5028cc340988f7c37f2e0 <= Icb2a399b8ac8449ff9ff8e5986aac03d;
 I186a56ca3712df6983eb742d7d80a37e <= I933a5eb08d4d1445f167a74db5fbdc75;
 I389856ba7ca6568e4ead3483c3e52353 <= I9c046caddde3b171774d3eba258190f0;
 I66b39fb4c54ab32b2c876813544ff6bc <= Ic8f12fefb9c055923e2842aeca48765f;
 I591624fd56ff315e0084af5af206cf8e <= I26631e7940eb983e49a9313da628e23a;
 I3994dd74d52d8957e443e869cbbf7184 <= I7fac6686ca9a63213ec3cdee4b812daa;
 I92793401ab28d5ed265775c0d165dfe5 <= I1960eba710ca20ef749501b02fd3b0bd;
 Ic499c718cc4866eb8536d66ae4fae0e4 <= Ie1f5cc89163ee091f938a4c3edaca65b;
 I3c28bfe18fb1543683ae264c396a0207 <= I63e7cf958a0de50d3299d2077d8cb192;
 I083aca08b0d0bd2622d0f7b6b2aaeb99 <= I50c2132c2b5e60af7ba2b9be8c90d9a4;
 I2fd3c0dfd43b65e2fe8afd3368a50fc5 <= If1243756e31d0a56b6666cad5b21f731;
 I58332f7615e647e757033f6b643c21a4 <= I92c03e59c3f96f63800051762f6949c0;
 I22bbdf426df953feb5acede78c31b9b2 <= I488d337ed967adebd6c580b7203991b5;
 Ia9f7a93a673c49ef3bfffd6fcadf845a <= I32aa0d9a082eb6a595467f3c7f36a3f7;
 I687ab1878d38c7c988507163c8a60070 <= Iec440f37d189fbcd4c06cf34344c4439;
 I9efb470a3342962583f19eaec3a0ecd7 <= I66d815daa51bcda0d549dbcc9c027195;
 Id7f7499e9b3f529781f4aba6e63490ac <= I192d10feae906d5ef90b4a90398d3ced;
 I88e14285aa13b58457c58439ad1c8c87 <= I1d8d269f64d0d3041bc69d879a3654ab;
 I730aeccac38e1622c684c468f8cb29f4 <= I5fce715f064098fe4685479aede832e7;
 I9427589efc5ae29474734dcc6e36ea81 <= I1b65989684c087f328e3fb58d3a3395e;
 Iba910435a91ee873f76fa3ec9ac9c3d3 <= I5352562c002801df06f847362d347180;
 Ia3c2d3cea56571481655cc77ee025558 <= I176397bab05ee39f7d54a28c5f74c3cc;
 I99ba3451537a2876c9f585f72911bc4f <=  start_d_fgallag0x00000;
end
