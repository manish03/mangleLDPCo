 reg  ['h0:0] [$clog2('h7000+1)-1:0] Ib10d67e2c07b1438e202f7b58974fa8e94cfa1651476e39e36cd90f61705d1c2 ;
