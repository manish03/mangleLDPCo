 reg  ['h3fff:0] [$clog2('h7000+1)-1:0] Ifd35529b44c957737bf422127283c08e ;
