//`include "GF2_LDPC_flogtanh_0x00006_assign_inc.sv"
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00000] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00000] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00001] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00001] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00002] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00003] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00002] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00004] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00005] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00003] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00006] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00007] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00004] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00008] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00009] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00005] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0000a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0000b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00006] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0000c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0000d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00007] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0000e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0000f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00008] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00010] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00011] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00009] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00012] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00013] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000a] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00014] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00015] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000b] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00016] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00017] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000c] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00018] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00019] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000d] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0001a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0001b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000e] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0001c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0001d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0000f] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0001e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0001f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00010] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00020] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00021] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00011] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00022] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00023] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00012] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00024] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00025] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00013] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00026] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00027] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00014] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00028] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00029] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00015] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0002a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0002b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00016] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0002c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0002d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00017] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0002e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0002f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00018] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00030] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00031] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00019] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00032] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00033] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001a] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00034] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00035] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001b] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00036] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00037] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001c] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00038] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00039] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001d] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0003a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0003b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001e] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0003c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0003d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0001f] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0003e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0003f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00020] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00040] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00041] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00021] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00042] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00043] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00022] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00044] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00045] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00023] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00046] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00047] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00024] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00048] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00049] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00025] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0004a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0004b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00026] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0004c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0004d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00027] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0004e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0004f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00028] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00050] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00051] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00029] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00052] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00053] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002a] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00054] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00055] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002b] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00056] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00057] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002c] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00058] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00059] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002d] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0005a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0005b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002e] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0005c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0005d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0002f] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0005e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0005f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00030] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00060] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00061] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00031] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00062] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00063] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00032] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00064] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00065] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00033] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00066] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00067] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00034] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00068] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00069] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00035] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0006a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0006b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00036] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0006c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0006d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00037] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0006e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0006f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00038] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00070] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00071] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00039] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00072] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00073] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003a] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00074] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00075] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003b] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00076] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00077] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003c] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00078] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00079] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003d] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0007a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0007b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003e] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0007c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0007d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0003f] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0007e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0007f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00040] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00080] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00081] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00041] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00082] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00083] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00042] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00084] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00085] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00043] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00086] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00087] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00044] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00088] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00089] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00045] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0008a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0008b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00046] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0008c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0008d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00047] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0008e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0008f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00048] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00090] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00091] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00049] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00092] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00093] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004a] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00094] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00095] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004b] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00096] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00097] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004c] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00098] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00099] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004d] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0009a] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0009b] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004e] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0009c] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0009d] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0004f] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h0009e] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h0009f] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00050] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a0] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a1] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00051] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a2] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a3] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00052] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a4] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a5] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00053] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a6] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a7] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00054] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a8] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000a9] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00055] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000aa] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000ab] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00056] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000ac] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000ad] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00057] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000ae] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000af] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00058] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b0] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b1] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00059] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b2] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b3] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005a] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b4] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b5] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005b] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b6] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b7] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005c] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b8] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000b9] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005d] =  Ifcca41d795dde8a35d1654b9520c92e7['h000ba] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005e] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000bc] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000bd] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0005f] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000be] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000bf] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00060] =  Ifcca41d795dde8a35d1654b9520c92e7['h000c0] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00061] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000c2] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000c3] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00062] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000c4] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000c5] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00063] =  Ifcca41d795dde8a35d1654b9520c92e7['h000c6] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00064] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000c8] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000c9] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00065] =  Ifcca41d795dde8a35d1654b9520c92e7['h000ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00066] =  Ifcca41d795dde8a35d1654b9520c92e7['h000cc] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00067] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000ce] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000cf] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00068] =  Ifcca41d795dde8a35d1654b9520c92e7['h000d0] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00069] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000d2] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000d3] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006a] =  Ifcca41d795dde8a35d1654b9520c92e7['h000d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006b] =  Ifcca41d795dde8a35d1654b9520c92e7['h000d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006c] =  Ifcca41d795dde8a35d1654b9520c92e7['h000d8] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006d] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000da] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000db] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006e] =  Ifcca41d795dde8a35d1654b9520c92e7['h000dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0006f] =  Ifcca41d795dde8a35d1654b9520c92e7['h000de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00070] =  Ifcca41d795dde8a35d1654b9520c92e7['h000e0] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00071] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000e2] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000e3] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00072] =  Ifcca41d795dde8a35d1654b9520c92e7['h000e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00073] =  Ifcca41d795dde8a35d1654b9520c92e7['h000e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00074] =  Ifcca41d795dde8a35d1654b9520c92e7['h000e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00075] =  Ifcca41d795dde8a35d1654b9520c92e7['h000ea] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00076] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000ec] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000ed] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00077] =  Ifcca41d795dde8a35d1654b9520c92e7['h000ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00078] =  Ifcca41d795dde8a35d1654b9520c92e7['h000f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00079] =  Ifcca41d795dde8a35d1654b9520c92e7['h000f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007a] =  Ifcca41d795dde8a35d1654b9520c92e7['h000f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007b] =  Ifcca41d795dde8a35d1654b9520c92e7['h000f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007c] =  Ifcca41d795dde8a35d1654b9520c92e7['h000f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007d] =  Ifcca41d795dde8a35d1654b9520c92e7['h000fa] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007e] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h000fc] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h000fd] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0007f] =  Ifcca41d795dde8a35d1654b9520c92e7['h000fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00080] =  Ifcca41d795dde8a35d1654b9520c92e7['h00100] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00081] =  Ifcca41d795dde8a35d1654b9520c92e7['h00102] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00082] =  Ifcca41d795dde8a35d1654b9520c92e7['h00104] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00083] =  Ifcca41d795dde8a35d1654b9520c92e7['h00106] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00084] =  Ifcca41d795dde8a35d1654b9520c92e7['h00108] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00085] =  Ifcca41d795dde8a35d1654b9520c92e7['h0010a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00086] =  Ifcca41d795dde8a35d1654b9520c92e7['h0010c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00087] =  Ifcca41d795dde8a35d1654b9520c92e7['h0010e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00088] =  Ifcca41d795dde8a35d1654b9520c92e7['h00110] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00089] =  Ifcca41d795dde8a35d1654b9520c92e7['h00112] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00114] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00116] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00118] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0011a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0011c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0008f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0011e] ;
//end
//always_comb begin
              I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00090] = 
          (!flogtanh_sel['h00006]) ? 
                       Ifcca41d795dde8a35d1654b9520c92e7['h00120] : //%
                       Ifcca41d795dde8a35d1654b9520c92e7['h00121] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00091] =  Ifcca41d795dde8a35d1654b9520c92e7['h00122] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00092] =  Ifcca41d795dde8a35d1654b9520c92e7['h00124] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00093] =  Ifcca41d795dde8a35d1654b9520c92e7['h00126] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00094] =  Ifcca41d795dde8a35d1654b9520c92e7['h00128] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00095] =  Ifcca41d795dde8a35d1654b9520c92e7['h0012a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00096] =  Ifcca41d795dde8a35d1654b9520c92e7['h0012c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00097] =  Ifcca41d795dde8a35d1654b9520c92e7['h0012e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00098] =  Ifcca41d795dde8a35d1654b9520c92e7['h00130] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00099] =  Ifcca41d795dde8a35d1654b9520c92e7['h00132] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00134] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00136] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00138] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0013a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0013c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0009f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0013e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00140] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00142] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00144] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00146] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00148] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0014a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0014c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0014e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00150] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00152] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00154] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h00156] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h00158] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0015a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0015c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000af] =  Ifcca41d795dde8a35d1654b9520c92e7['h0015e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00160] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00162] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00164] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00166] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00168] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0016a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0016c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0016e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00170] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00172] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h00174] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00176] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00178] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0017a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000be] =  Ifcca41d795dde8a35d1654b9520c92e7['h0017c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0017e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00180] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00182] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00184] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00186] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00188] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0018a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0018c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0018e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00190] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00192] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h00194] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00196] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00198] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0019a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0019c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0019e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h001a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h001a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h001a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h001a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h001a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h001aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h001ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h001ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h001b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h001b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000da] =  Ifcca41d795dde8a35d1654b9520c92e7['h001b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000db] =  Ifcca41d795dde8a35d1654b9520c92e7['h001b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h001b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h001ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000de] =  Ifcca41d795dde8a35d1654b9520c92e7['h001bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000df] =  Ifcca41d795dde8a35d1654b9520c92e7['h001be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h001c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h001c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h001c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h001c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h001c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h001ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h001cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h001ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h001d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h001d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h001d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h001d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h001d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h001da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h001dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h001de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h001e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h001e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h001e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h001e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h001e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h001ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h001ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h001ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h001f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h001f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h001f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h001f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h001f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h001fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h001fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h000ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h001fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00100] =  Ifcca41d795dde8a35d1654b9520c92e7['h00200] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00101] =  Ifcca41d795dde8a35d1654b9520c92e7['h00202] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00102] =  Ifcca41d795dde8a35d1654b9520c92e7['h00204] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00103] =  Ifcca41d795dde8a35d1654b9520c92e7['h00206] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00104] =  Ifcca41d795dde8a35d1654b9520c92e7['h00208] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00105] =  Ifcca41d795dde8a35d1654b9520c92e7['h0020a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00106] =  Ifcca41d795dde8a35d1654b9520c92e7['h0020c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00107] =  Ifcca41d795dde8a35d1654b9520c92e7['h0020e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00108] =  Ifcca41d795dde8a35d1654b9520c92e7['h00210] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00109] =  Ifcca41d795dde8a35d1654b9520c92e7['h00212] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00214] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00216] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00218] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0021a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0021c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0010f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0021e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00110] =  Ifcca41d795dde8a35d1654b9520c92e7['h00220] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00111] =  Ifcca41d795dde8a35d1654b9520c92e7['h00222] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00112] =  Ifcca41d795dde8a35d1654b9520c92e7['h00224] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00113] =  Ifcca41d795dde8a35d1654b9520c92e7['h00226] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00114] =  Ifcca41d795dde8a35d1654b9520c92e7['h00228] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00115] =  Ifcca41d795dde8a35d1654b9520c92e7['h0022a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00116] =  Ifcca41d795dde8a35d1654b9520c92e7['h0022c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00117] =  Ifcca41d795dde8a35d1654b9520c92e7['h0022e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00118] =  Ifcca41d795dde8a35d1654b9520c92e7['h00230] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00119] =  Ifcca41d795dde8a35d1654b9520c92e7['h00232] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00234] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00236] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00238] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0023a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0023c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0011f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0023e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00120] =  Ifcca41d795dde8a35d1654b9520c92e7['h00240] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00121] =  Ifcca41d795dde8a35d1654b9520c92e7['h00242] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00122] =  Ifcca41d795dde8a35d1654b9520c92e7['h00244] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00123] =  Ifcca41d795dde8a35d1654b9520c92e7['h00246] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00124] =  Ifcca41d795dde8a35d1654b9520c92e7['h00248] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00125] =  Ifcca41d795dde8a35d1654b9520c92e7['h0024a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00126] =  Ifcca41d795dde8a35d1654b9520c92e7['h0024c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00127] =  Ifcca41d795dde8a35d1654b9520c92e7['h0024e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00128] =  Ifcca41d795dde8a35d1654b9520c92e7['h00250] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00129] =  Ifcca41d795dde8a35d1654b9520c92e7['h00252] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00254] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00256] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00258] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0025a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0025c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0012f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0025e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00130] =  Ifcca41d795dde8a35d1654b9520c92e7['h00260] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00131] =  Ifcca41d795dde8a35d1654b9520c92e7['h00262] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00132] =  Ifcca41d795dde8a35d1654b9520c92e7['h00264] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00133] =  Ifcca41d795dde8a35d1654b9520c92e7['h00266] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00134] =  Ifcca41d795dde8a35d1654b9520c92e7['h00268] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00135] =  Ifcca41d795dde8a35d1654b9520c92e7['h0026a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00136] =  Ifcca41d795dde8a35d1654b9520c92e7['h0026c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00137] =  Ifcca41d795dde8a35d1654b9520c92e7['h0026e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00138] =  Ifcca41d795dde8a35d1654b9520c92e7['h00270] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00139] =  Ifcca41d795dde8a35d1654b9520c92e7['h00272] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00274] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00276] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00278] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0027a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0027c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0013f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0027e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00140] =  Ifcca41d795dde8a35d1654b9520c92e7['h00280] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00141] =  Ifcca41d795dde8a35d1654b9520c92e7['h00282] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00142] =  Ifcca41d795dde8a35d1654b9520c92e7['h00284] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00143] =  Ifcca41d795dde8a35d1654b9520c92e7['h00286] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00144] =  Ifcca41d795dde8a35d1654b9520c92e7['h00288] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00145] =  Ifcca41d795dde8a35d1654b9520c92e7['h0028a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00146] =  Ifcca41d795dde8a35d1654b9520c92e7['h0028c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00147] =  Ifcca41d795dde8a35d1654b9520c92e7['h0028e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00148] =  Ifcca41d795dde8a35d1654b9520c92e7['h00290] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00149] =  Ifcca41d795dde8a35d1654b9520c92e7['h00292] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00294] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00296] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00298] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0029a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0029c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0014f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0029e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00150] =  Ifcca41d795dde8a35d1654b9520c92e7['h002a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00151] =  Ifcca41d795dde8a35d1654b9520c92e7['h002a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00152] =  Ifcca41d795dde8a35d1654b9520c92e7['h002a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00153] =  Ifcca41d795dde8a35d1654b9520c92e7['h002a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00154] =  Ifcca41d795dde8a35d1654b9520c92e7['h002a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00155] =  Ifcca41d795dde8a35d1654b9520c92e7['h002aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00156] =  Ifcca41d795dde8a35d1654b9520c92e7['h002ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00157] =  Ifcca41d795dde8a35d1654b9520c92e7['h002ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00158] =  Ifcca41d795dde8a35d1654b9520c92e7['h002b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00159] =  Ifcca41d795dde8a35d1654b9520c92e7['h002b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015a] =  Ifcca41d795dde8a35d1654b9520c92e7['h002b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015b] =  Ifcca41d795dde8a35d1654b9520c92e7['h002b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015c] =  Ifcca41d795dde8a35d1654b9520c92e7['h002b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015d] =  Ifcca41d795dde8a35d1654b9520c92e7['h002ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015e] =  Ifcca41d795dde8a35d1654b9520c92e7['h002bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0015f] =  Ifcca41d795dde8a35d1654b9520c92e7['h002be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00160] =  Ifcca41d795dde8a35d1654b9520c92e7['h002c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00161] =  Ifcca41d795dde8a35d1654b9520c92e7['h002c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00162] =  Ifcca41d795dde8a35d1654b9520c92e7['h002c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00163] =  Ifcca41d795dde8a35d1654b9520c92e7['h002c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00164] =  Ifcca41d795dde8a35d1654b9520c92e7['h002c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00165] =  Ifcca41d795dde8a35d1654b9520c92e7['h002ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00166] =  Ifcca41d795dde8a35d1654b9520c92e7['h002cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00167] =  Ifcca41d795dde8a35d1654b9520c92e7['h002ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00168] =  Ifcca41d795dde8a35d1654b9520c92e7['h002d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00169] =  Ifcca41d795dde8a35d1654b9520c92e7['h002d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016a] =  Ifcca41d795dde8a35d1654b9520c92e7['h002d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016b] =  Ifcca41d795dde8a35d1654b9520c92e7['h002d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016c] =  Ifcca41d795dde8a35d1654b9520c92e7['h002d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016d] =  Ifcca41d795dde8a35d1654b9520c92e7['h002da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016e] =  Ifcca41d795dde8a35d1654b9520c92e7['h002dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0016f] =  Ifcca41d795dde8a35d1654b9520c92e7['h002de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00170] =  Ifcca41d795dde8a35d1654b9520c92e7['h002e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00171] =  Ifcca41d795dde8a35d1654b9520c92e7['h002e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00172] =  Ifcca41d795dde8a35d1654b9520c92e7['h002e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00173] =  Ifcca41d795dde8a35d1654b9520c92e7['h002e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00174] =  Ifcca41d795dde8a35d1654b9520c92e7['h002e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00175] =  Ifcca41d795dde8a35d1654b9520c92e7['h002ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00176] =  Ifcca41d795dde8a35d1654b9520c92e7['h002ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00177] =  Ifcca41d795dde8a35d1654b9520c92e7['h002ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00178] =  Ifcca41d795dde8a35d1654b9520c92e7['h002f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00179] =  Ifcca41d795dde8a35d1654b9520c92e7['h002f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017a] =  Ifcca41d795dde8a35d1654b9520c92e7['h002f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017b] =  Ifcca41d795dde8a35d1654b9520c92e7['h002f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017c] =  Ifcca41d795dde8a35d1654b9520c92e7['h002f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017d] =  Ifcca41d795dde8a35d1654b9520c92e7['h002fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017e] =  Ifcca41d795dde8a35d1654b9520c92e7['h002fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0017f] =  Ifcca41d795dde8a35d1654b9520c92e7['h002fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00180] =  Ifcca41d795dde8a35d1654b9520c92e7['h00300] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00181] =  Ifcca41d795dde8a35d1654b9520c92e7['h00302] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00182] =  Ifcca41d795dde8a35d1654b9520c92e7['h00304] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00183] =  Ifcca41d795dde8a35d1654b9520c92e7['h00306] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00184] =  Ifcca41d795dde8a35d1654b9520c92e7['h00308] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00185] =  Ifcca41d795dde8a35d1654b9520c92e7['h0030a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00186] =  Ifcca41d795dde8a35d1654b9520c92e7['h0030c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00187] =  Ifcca41d795dde8a35d1654b9520c92e7['h0030e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00188] =  Ifcca41d795dde8a35d1654b9520c92e7['h00310] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00189] =  Ifcca41d795dde8a35d1654b9520c92e7['h00312] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00314] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00316] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00318] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0031a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0031c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0018f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0031e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00190] =  Ifcca41d795dde8a35d1654b9520c92e7['h00320] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00191] =  Ifcca41d795dde8a35d1654b9520c92e7['h00322] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00192] =  Ifcca41d795dde8a35d1654b9520c92e7['h00324] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00193] =  Ifcca41d795dde8a35d1654b9520c92e7['h00326] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00194] =  Ifcca41d795dde8a35d1654b9520c92e7['h00328] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00195] =  Ifcca41d795dde8a35d1654b9520c92e7['h0032a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00196] =  Ifcca41d795dde8a35d1654b9520c92e7['h0032c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00197] =  Ifcca41d795dde8a35d1654b9520c92e7['h0032e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00198] =  Ifcca41d795dde8a35d1654b9520c92e7['h00330] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00199] =  Ifcca41d795dde8a35d1654b9520c92e7['h00332] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00334] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00336] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00338] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0033a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0033c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0019f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0033e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00340] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00342] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00344] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00346] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00348] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0034a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0034c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0034e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00350] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00352] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00354] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h00356] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h00358] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0035a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0035c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001af] =  Ifcca41d795dde8a35d1654b9520c92e7['h0035e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00360] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00362] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00364] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00366] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00368] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0036a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0036c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0036e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00370] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00372] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h00374] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00376] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00378] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0037a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001be] =  Ifcca41d795dde8a35d1654b9520c92e7['h0037c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0037e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00380] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00382] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00384] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00386] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00388] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0038a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0038c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0038e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00390] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00392] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h00394] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00396] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00398] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0039a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0039c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0039e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h003a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h003a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h003a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h003a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h003a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h003aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h003ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h003ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h003b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h003b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001da] =  Ifcca41d795dde8a35d1654b9520c92e7['h003b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001db] =  Ifcca41d795dde8a35d1654b9520c92e7['h003b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h003b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h003ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001de] =  Ifcca41d795dde8a35d1654b9520c92e7['h003bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001df] =  Ifcca41d795dde8a35d1654b9520c92e7['h003be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h003c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h003c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h003c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h003c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h003c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h003ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h003cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h003ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h003d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h003d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h003d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h003d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h003d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h003da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h003dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h003de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h003e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h003e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h003e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h003e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h003e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h003ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h003ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h003ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h003f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h003f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h003f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h003f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h003f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h003fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h003fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h001ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h003fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00200] =  Ifcca41d795dde8a35d1654b9520c92e7['h00400] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00201] =  Ifcca41d795dde8a35d1654b9520c92e7['h00402] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00202] =  Ifcca41d795dde8a35d1654b9520c92e7['h00404] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00203] =  Ifcca41d795dde8a35d1654b9520c92e7['h00406] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00204] =  Ifcca41d795dde8a35d1654b9520c92e7['h00408] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00205] =  Ifcca41d795dde8a35d1654b9520c92e7['h0040a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00206] =  Ifcca41d795dde8a35d1654b9520c92e7['h0040c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00207] =  Ifcca41d795dde8a35d1654b9520c92e7['h0040e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00208] =  Ifcca41d795dde8a35d1654b9520c92e7['h00410] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00209] =  Ifcca41d795dde8a35d1654b9520c92e7['h00412] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00414] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00416] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00418] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0041a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0041c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0020f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0041e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00210] =  Ifcca41d795dde8a35d1654b9520c92e7['h00420] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00211] =  Ifcca41d795dde8a35d1654b9520c92e7['h00422] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00212] =  Ifcca41d795dde8a35d1654b9520c92e7['h00424] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00213] =  Ifcca41d795dde8a35d1654b9520c92e7['h00426] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00214] =  Ifcca41d795dde8a35d1654b9520c92e7['h00428] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00215] =  Ifcca41d795dde8a35d1654b9520c92e7['h0042a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00216] =  Ifcca41d795dde8a35d1654b9520c92e7['h0042c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00217] =  Ifcca41d795dde8a35d1654b9520c92e7['h0042e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00218] =  Ifcca41d795dde8a35d1654b9520c92e7['h00430] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00219] =  Ifcca41d795dde8a35d1654b9520c92e7['h00432] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00434] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00436] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00438] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0043a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0043c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0021f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0043e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00220] =  Ifcca41d795dde8a35d1654b9520c92e7['h00440] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00221] =  Ifcca41d795dde8a35d1654b9520c92e7['h00442] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00222] =  Ifcca41d795dde8a35d1654b9520c92e7['h00444] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00223] =  Ifcca41d795dde8a35d1654b9520c92e7['h00446] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00224] =  Ifcca41d795dde8a35d1654b9520c92e7['h00448] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00225] =  Ifcca41d795dde8a35d1654b9520c92e7['h0044a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00226] =  Ifcca41d795dde8a35d1654b9520c92e7['h0044c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00227] =  Ifcca41d795dde8a35d1654b9520c92e7['h0044e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00228] =  Ifcca41d795dde8a35d1654b9520c92e7['h00450] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00229] =  Ifcca41d795dde8a35d1654b9520c92e7['h00452] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00454] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00456] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00458] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0045a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0045c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0022f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0045e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00230] =  Ifcca41d795dde8a35d1654b9520c92e7['h00460] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00231] =  Ifcca41d795dde8a35d1654b9520c92e7['h00462] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00232] =  Ifcca41d795dde8a35d1654b9520c92e7['h00464] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00233] =  Ifcca41d795dde8a35d1654b9520c92e7['h00466] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00234] =  Ifcca41d795dde8a35d1654b9520c92e7['h00468] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00235] =  Ifcca41d795dde8a35d1654b9520c92e7['h0046a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00236] =  Ifcca41d795dde8a35d1654b9520c92e7['h0046c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00237] =  Ifcca41d795dde8a35d1654b9520c92e7['h0046e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00238] =  Ifcca41d795dde8a35d1654b9520c92e7['h00470] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00239] =  Ifcca41d795dde8a35d1654b9520c92e7['h00472] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00474] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00476] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00478] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0047a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0047c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0023f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0047e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00240] =  Ifcca41d795dde8a35d1654b9520c92e7['h00480] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00241] =  Ifcca41d795dde8a35d1654b9520c92e7['h00482] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00242] =  Ifcca41d795dde8a35d1654b9520c92e7['h00484] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00243] =  Ifcca41d795dde8a35d1654b9520c92e7['h00486] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00244] =  Ifcca41d795dde8a35d1654b9520c92e7['h00488] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00245] =  Ifcca41d795dde8a35d1654b9520c92e7['h0048a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00246] =  Ifcca41d795dde8a35d1654b9520c92e7['h0048c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00247] =  Ifcca41d795dde8a35d1654b9520c92e7['h0048e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00248] =  Ifcca41d795dde8a35d1654b9520c92e7['h00490] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00249] =  Ifcca41d795dde8a35d1654b9520c92e7['h00492] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00494] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00496] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00498] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0049a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0049c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0024f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0049e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00250] =  Ifcca41d795dde8a35d1654b9520c92e7['h004a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00251] =  Ifcca41d795dde8a35d1654b9520c92e7['h004a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00252] =  Ifcca41d795dde8a35d1654b9520c92e7['h004a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00253] =  Ifcca41d795dde8a35d1654b9520c92e7['h004a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00254] =  Ifcca41d795dde8a35d1654b9520c92e7['h004a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00255] =  Ifcca41d795dde8a35d1654b9520c92e7['h004aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00256] =  Ifcca41d795dde8a35d1654b9520c92e7['h004ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00257] =  Ifcca41d795dde8a35d1654b9520c92e7['h004ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00258] =  Ifcca41d795dde8a35d1654b9520c92e7['h004b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00259] =  Ifcca41d795dde8a35d1654b9520c92e7['h004b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025a] =  Ifcca41d795dde8a35d1654b9520c92e7['h004b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025b] =  Ifcca41d795dde8a35d1654b9520c92e7['h004b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025c] =  Ifcca41d795dde8a35d1654b9520c92e7['h004b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025d] =  Ifcca41d795dde8a35d1654b9520c92e7['h004ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025e] =  Ifcca41d795dde8a35d1654b9520c92e7['h004bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0025f] =  Ifcca41d795dde8a35d1654b9520c92e7['h004be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00260] =  Ifcca41d795dde8a35d1654b9520c92e7['h004c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00261] =  Ifcca41d795dde8a35d1654b9520c92e7['h004c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00262] =  Ifcca41d795dde8a35d1654b9520c92e7['h004c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00263] =  Ifcca41d795dde8a35d1654b9520c92e7['h004c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00264] =  Ifcca41d795dde8a35d1654b9520c92e7['h004c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00265] =  Ifcca41d795dde8a35d1654b9520c92e7['h004ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00266] =  Ifcca41d795dde8a35d1654b9520c92e7['h004cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00267] =  Ifcca41d795dde8a35d1654b9520c92e7['h004ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00268] =  Ifcca41d795dde8a35d1654b9520c92e7['h004d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00269] =  Ifcca41d795dde8a35d1654b9520c92e7['h004d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026a] =  Ifcca41d795dde8a35d1654b9520c92e7['h004d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026b] =  Ifcca41d795dde8a35d1654b9520c92e7['h004d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026c] =  Ifcca41d795dde8a35d1654b9520c92e7['h004d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026d] =  Ifcca41d795dde8a35d1654b9520c92e7['h004da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026e] =  Ifcca41d795dde8a35d1654b9520c92e7['h004dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0026f] =  Ifcca41d795dde8a35d1654b9520c92e7['h004de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00270] =  Ifcca41d795dde8a35d1654b9520c92e7['h004e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00271] =  Ifcca41d795dde8a35d1654b9520c92e7['h004e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00272] =  Ifcca41d795dde8a35d1654b9520c92e7['h004e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00273] =  Ifcca41d795dde8a35d1654b9520c92e7['h004e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00274] =  Ifcca41d795dde8a35d1654b9520c92e7['h004e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00275] =  Ifcca41d795dde8a35d1654b9520c92e7['h004ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00276] =  Ifcca41d795dde8a35d1654b9520c92e7['h004ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00277] =  Ifcca41d795dde8a35d1654b9520c92e7['h004ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00278] =  Ifcca41d795dde8a35d1654b9520c92e7['h004f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00279] =  Ifcca41d795dde8a35d1654b9520c92e7['h004f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027a] =  Ifcca41d795dde8a35d1654b9520c92e7['h004f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027b] =  Ifcca41d795dde8a35d1654b9520c92e7['h004f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027c] =  Ifcca41d795dde8a35d1654b9520c92e7['h004f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027d] =  Ifcca41d795dde8a35d1654b9520c92e7['h004fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027e] =  Ifcca41d795dde8a35d1654b9520c92e7['h004fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0027f] =  Ifcca41d795dde8a35d1654b9520c92e7['h004fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00280] =  Ifcca41d795dde8a35d1654b9520c92e7['h00500] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00281] =  Ifcca41d795dde8a35d1654b9520c92e7['h00502] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00282] =  Ifcca41d795dde8a35d1654b9520c92e7['h00504] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00283] =  Ifcca41d795dde8a35d1654b9520c92e7['h00506] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00284] =  Ifcca41d795dde8a35d1654b9520c92e7['h00508] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00285] =  Ifcca41d795dde8a35d1654b9520c92e7['h0050a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00286] =  Ifcca41d795dde8a35d1654b9520c92e7['h0050c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00287] =  Ifcca41d795dde8a35d1654b9520c92e7['h0050e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00288] =  Ifcca41d795dde8a35d1654b9520c92e7['h00510] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00289] =  Ifcca41d795dde8a35d1654b9520c92e7['h00512] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00514] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00516] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00518] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0051a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0051c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0028f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0051e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00290] =  Ifcca41d795dde8a35d1654b9520c92e7['h00520] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00291] =  Ifcca41d795dde8a35d1654b9520c92e7['h00522] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00292] =  Ifcca41d795dde8a35d1654b9520c92e7['h00524] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00293] =  Ifcca41d795dde8a35d1654b9520c92e7['h00526] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00294] =  Ifcca41d795dde8a35d1654b9520c92e7['h00528] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00295] =  Ifcca41d795dde8a35d1654b9520c92e7['h0052a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00296] =  Ifcca41d795dde8a35d1654b9520c92e7['h0052c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00297] =  Ifcca41d795dde8a35d1654b9520c92e7['h0052e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00298] =  Ifcca41d795dde8a35d1654b9520c92e7['h00530] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00299] =  Ifcca41d795dde8a35d1654b9520c92e7['h00532] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00534] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00536] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00538] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0053a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0053c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0029f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0053e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00540] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00542] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00544] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00546] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00548] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0054a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0054c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0054e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00550] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00552] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00554] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h00556] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h00558] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0055a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0055c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002af] =  Ifcca41d795dde8a35d1654b9520c92e7['h0055e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00560] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00562] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00564] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00566] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00568] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0056a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0056c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0056e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00570] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00572] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h00574] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00576] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00578] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0057a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002be] =  Ifcca41d795dde8a35d1654b9520c92e7['h0057c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0057e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00580] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00582] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00584] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00586] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00588] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0058a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0058c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0058e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00590] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00592] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h00594] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00596] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00598] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0059a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0059c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0059e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h005a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h005a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h005a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h005a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h005a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h005aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h005ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h005ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h005b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h005b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002da] =  Ifcca41d795dde8a35d1654b9520c92e7['h005b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002db] =  Ifcca41d795dde8a35d1654b9520c92e7['h005b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h005b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h005ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002de] =  Ifcca41d795dde8a35d1654b9520c92e7['h005bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002df] =  Ifcca41d795dde8a35d1654b9520c92e7['h005be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h005c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h005c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h005c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h005c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h005c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h005ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h005cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h005ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h005d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h005d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h005d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h005d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h005d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h005da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h005dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h005de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h005e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h005e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h005e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h005e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h005e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h005ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h005ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h005ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h005f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h005f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h005f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h005f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h005f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h005fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h005fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h002ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h005fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00300] =  Ifcca41d795dde8a35d1654b9520c92e7['h00600] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00301] =  Ifcca41d795dde8a35d1654b9520c92e7['h00602] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00302] =  Ifcca41d795dde8a35d1654b9520c92e7['h00604] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00303] =  Ifcca41d795dde8a35d1654b9520c92e7['h00606] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00304] =  Ifcca41d795dde8a35d1654b9520c92e7['h00608] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00305] =  Ifcca41d795dde8a35d1654b9520c92e7['h0060a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00306] =  Ifcca41d795dde8a35d1654b9520c92e7['h0060c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00307] =  Ifcca41d795dde8a35d1654b9520c92e7['h0060e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00308] =  Ifcca41d795dde8a35d1654b9520c92e7['h00610] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00309] =  Ifcca41d795dde8a35d1654b9520c92e7['h00612] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00614] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00616] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00618] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0061a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0061c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0030f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0061e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00310] =  Ifcca41d795dde8a35d1654b9520c92e7['h00620] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00311] =  Ifcca41d795dde8a35d1654b9520c92e7['h00622] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00312] =  Ifcca41d795dde8a35d1654b9520c92e7['h00624] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00313] =  Ifcca41d795dde8a35d1654b9520c92e7['h00626] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00314] =  Ifcca41d795dde8a35d1654b9520c92e7['h00628] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00315] =  Ifcca41d795dde8a35d1654b9520c92e7['h0062a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00316] =  Ifcca41d795dde8a35d1654b9520c92e7['h0062c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00317] =  Ifcca41d795dde8a35d1654b9520c92e7['h0062e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00318] =  Ifcca41d795dde8a35d1654b9520c92e7['h00630] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00319] =  Ifcca41d795dde8a35d1654b9520c92e7['h00632] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00634] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00636] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00638] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0063a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0063c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0031f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0063e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00320] =  Ifcca41d795dde8a35d1654b9520c92e7['h00640] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00321] =  Ifcca41d795dde8a35d1654b9520c92e7['h00642] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00322] =  Ifcca41d795dde8a35d1654b9520c92e7['h00644] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00323] =  Ifcca41d795dde8a35d1654b9520c92e7['h00646] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00324] =  Ifcca41d795dde8a35d1654b9520c92e7['h00648] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00325] =  Ifcca41d795dde8a35d1654b9520c92e7['h0064a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00326] =  Ifcca41d795dde8a35d1654b9520c92e7['h0064c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00327] =  Ifcca41d795dde8a35d1654b9520c92e7['h0064e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00328] =  Ifcca41d795dde8a35d1654b9520c92e7['h00650] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00329] =  Ifcca41d795dde8a35d1654b9520c92e7['h00652] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00654] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00656] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00658] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0065a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0065c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0032f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0065e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00330] =  Ifcca41d795dde8a35d1654b9520c92e7['h00660] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00331] =  Ifcca41d795dde8a35d1654b9520c92e7['h00662] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00332] =  Ifcca41d795dde8a35d1654b9520c92e7['h00664] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00333] =  Ifcca41d795dde8a35d1654b9520c92e7['h00666] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00334] =  Ifcca41d795dde8a35d1654b9520c92e7['h00668] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00335] =  Ifcca41d795dde8a35d1654b9520c92e7['h0066a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00336] =  Ifcca41d795dde8a35d1654b9520c92e7['h0066c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00337] =  Ifcca41d795dde8a35d1654b9520c92e7['h0066e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00338] =  Ifcca41d795dde8a35d1654b9520c92e7['h00670] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00339] =  Ifcca41d795dde8a35d1654b9520c92e7['h00672] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00674] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00676] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00678] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0067a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0067c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0033f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0067e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00340] =  Ifcca41d795dde8a35d1654b9520c92e7['h00680] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00341] =  Ifcca41d795dde8a35d1654b9520c92e7['h00682] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00342] =  Ifcca41d795dde8a35d1654b9520c92e7['h00684] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00343] =  Ifcca41d795dde8a35d1654b9520c92e7['h00686] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00344] =  Ifcca41d795dde8a35d1654b9520c92e7['h00688] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00345] =  Ifcca41d795dde8a35d1654b9520c92e7['h0068a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00346] =  Ifcca41d795dde8a35d1654b9520c92e7['h0068c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00347] =  Ifcca41d795dde8a35d1654b9520c92e7['h0068e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00348] =  Ifcca41d795dde8a35d1654b9520c92e7['h00690] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00349] =  Ifcca41d795dde8a35d1654b9520c92e7['h00692] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00694] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00696] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00698] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0069a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0069c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0034f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0069e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00350] =  Ifcca41d795dde8a35d1654b9520c92e7['h006a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00351] =  Ifcca41d795dde8a35d1654b9520c92e7['h006a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00352] =  Ifcca41d795dde8a35d1654b9520c92e7['h006a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00353] =  Ifcca41d795dde8a35d1654b9520c92e7['h006a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00354] =  Ifcca41d795dde8a35d1654b9520c92e7['h006a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00355] =  Ifcca41d795dde8a35d1654b9520c92e7['h006aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00356] =  Ifcca41d795dde8a35d1654b9520c92e7['h006ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00357] =  Ifcca41d795dde8a35d1654b9520c92e7['h006ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00358] =  Ifcca41d795dde8a35d1654b9520c92e7['h006b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00359] =  Ifcca41d795dde8a35d1654b9520c92e7['h006b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035a] =  Ifcca41d795dde8a35d1654b9520c92e7['h006b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035b] =  Ifcca41d795dde8a35d1654b9520c92e7['h006b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035c] =  Ifcca41d795dde8a35d1654b9520c92e7['h006b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035d] =  Ifcca41d795dde8a35d1654b9520c92e7['h006ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035e] =  Ifcca41d795dde8a35d1654b9520c92e7['h006bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0035f] =  Ifcca41d795dde8a35d1654b9520c92e7['h006be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00360] =  Ifcca41d795dde8a35d1654b9520c92e7['h006c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00361] =  Ifcca41d795dde8a35d1654b9520c92e7['h006c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00362] =  Ifcca41d795dde8a35d1654b9520c92e7['h006c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00363] =  Ifcca41d795dde8a35d1654b9520c92e7['h006c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00364] =  Ifcca41d795dde8a35d1654b9520c92e7['h006c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00365] =  Ifcca41d795dde8a35d1654b9520c92e7['h006ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00366] =  Ifcca41d795dde8a35d1654b9520c92e7['h006cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00367] =  Ifcca41d795dde8a35d1654b9520c92e7['h006ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00368] =  Ifcca41d795dde8a35d1654b9520c92e7['h006d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00369] =  Ifcca41d795dde8a35d1654b9520c92e7['h006d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036a] =  Ifcca41d795dde8a35d1654b9520c92e7['h006d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036b] =  Ifcca41d795dde8a35d1654b9520c92e7['h006d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036c] =  Ifcca41d795dde8a35d1654b9520c92e7['h006d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036d] =  Ifcca41d795dde8a35d1654b9520c92e7['h006da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036e] =  Ifcca41d795dde8a35d1654b9520c92e7['h006dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0036f] =  Ifcca41d795dde8a35d1654b9520c92e7['h006de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00370] =  Ifcca41d795dde8a35d1654b9520c92e7['h006e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00371] =  Ifcca41d795dde8a35d1654b9520c92e7['h006e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00372] =  Ifcca41d795dde8a35d1654b9520c92e7['h006e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00373] =  Ifcca41d795dde8a35d1654b9520c92e7['h006e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00374] =  Ifcca41d795dde8a35d1654b9520c92e7['h006e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00375] =  Ifcca41d795dde8a35d1654b9520c92e7['h006ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00376] =  Ifcca41d795dde8a35d1654b9520c92e7['h006ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00377] =  Ifcca41d795dde8a35d1654b9520c92e7['h006ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00378] =  Ifcca41d795dde8a35d1654b9520c92e7['h006f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00379] =  Ifcca41d795dde8a35d1654b9520c92e7['h006f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037a] =  Ifcca41d795dde8a35d1654b9520c92e7['h006f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037b] =  Ifcca41d795dde8a35d1654b9520c92e7['h006f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037c] =  Ifcca41d795dde8a35d1654b9520c92e7['h006f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037d] =  Ifcca41d795dde8a35d1654b9520c92e7['h006fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037e] =  Ifcca41d795dde8a35d1654b9520c92e7['h006fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0037f] =  Ifcca41d795dde8a35d1654b9520c92e7['h006fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00380] =  Ifcca41d795dde8a35d1654b9520c92e7['h00700] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00381] =  Ifcca41d795dde8a35d1654b9520c92e7['h00702] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00382] =  Ifcca41d795dde8a35d1654b9520c92e7['h00704] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00383] =  Ifcca41d795dde8a35d1654b9520c92e7['h00706] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00384] =  Ifcca41d795dde8a35d1654b9520c92e7['h00708] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00385] =  Ifcca41d795dde8a35d1654b9520c92e7['h0070a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00386] =  Ifcca41d795dde8a35d1654b9520c92e7['h0070c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00387] =  Ifcca41d795dde8a35d1654b9520c92e7['h0070e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00388] =  Ifcca41d795dde8a35d1654b9520c92e7['h00710] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00389] =  Ifcca41d795dde8a35d1654b9520c92e7['h00712] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00714] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00716] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00718] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0071a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0071c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0038f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0071e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00390] =  Ifcca41d795dde8a35d1654b9520c92e7['h00720] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00391] =  Ifcca41d795dde8a35d1654b9520c92e7['h00722] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00392] =  Ifcca41d795dde8a35d1654b9520c92e7['h00724] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00393] =  Ifcca41d795dde8a35d1654b9520c92e7['h00726] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00394] =  Ifcca41d795dde8a35d1654b9520c92e7['h00728] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00395] =  Ifcca41d795dde8a35d1654b9520c92e7['h0072a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00396] =  Ifcca41d795dde8a35d1654b9520c92e7['h0072c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00397] =  Ifcca41d795dde8a35d1654b9520c92e7['h0072e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00398] =  Ifcca41d795dde8a35d1654b9520c92e7['h00730] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00399] =  Ifcca41d795dde8a35d1654b9520c92e7['h00732] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00734] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00736] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00738] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0073a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0073c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0039f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0073e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00740] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00742] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00744] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00746] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00748] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0074a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0074c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0074e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00750] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00752] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00754] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h00756] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h00758] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0075a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0075c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003af] =  Ifcca41d795dde8a35d1654b9520c92e7['h0075e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00760] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00762] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00764] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00766] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00768] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0076a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0076c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0076e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00770] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00772] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h00774] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00776] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00778] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0077a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003be] =  Ifcca41d795dde8a35d1654b9520c92e7['h0077c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0077e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00780] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00782] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00784] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00786] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00788] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0078a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0078c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0078e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00790] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00792] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h00794] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00796] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00798] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0079a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0079c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0079e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h007a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h007a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h007a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h007a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h007a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h007aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h007ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h007ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h007b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h007b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003da] =  Ifcca41d795dde8a35d1654b9520c92e7['h007b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003db] =  Ifcca41d795dde8a35d1654b9520c92e7['h007b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h007b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h007ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003de] =  Ifcca41d795dde8a35d1654b9520c92e7['h007bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003df] =  Ifcca41d795dde8a35d1654b9520c92e7['h007be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h007c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h007c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h007c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h007c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h007c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h007ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h007cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h007ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h007d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h007d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h007d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h007d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h007d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h007da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h007dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h007de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h007e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h007e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h007e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h007e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h007e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h007ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h007ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h007ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h007f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h007f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h007f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h007f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h007f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h007fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h007fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h003ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h007fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00400] =  Ifcca41d795dde8a35d1654b9520c92e7['h00800] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00401] =  Ifcca41d795dde8a35d1654b9520c92e7['h00802] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00402] =  Ifcca41d795dde8a35d1654b9520c92e7['h00804] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00403] =  Ifcca41d795dde8a35d1654b9520c92e7['h00806] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00404] =  Ifcca41d795dde8a35d1654b9520c92e7['h00808] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00405] =  Ifcca41d795dde8a35d1654b9520c92e7['h0080a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00406] =  Ifcca41d795dde8a35d1654b9520c92e7['h0080c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00407] =  Ifcca41d795dde8a35d1654b9520c92e7['h0080e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00408] =  Ifcca41d795dde8a35d1654b9520c92e7['h00810] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00409] =  Ifcca41d795dde8a35d1654b9520c92e7['h00812] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00814] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00816] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00818] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0081a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0081c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0040f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0081e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00410] =  Ifcca41d795dde8a35d1654b9520c92e7['h00820] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00411] =  Ifcca41d795dde8a35d1654b9520c92e7['h00822] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00412] =  Ifcca41d795dde8a35d1654b9520c92e7['h00824] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00413] =  Ifcca41d795dde8a35d1654b9520c92e7['h00826] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00414] =  Ifcca41d795dde8a35d1654b9520c92e7['h00828] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00415] =  Ifcca41d795dde8a35d1654b9520c92e7['h0082a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00416] =  Ifcca41d795dde8a35d1654b9520c92e7['h0082c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00417] =  Ifcca41d795dde8a35d1654b9520c92e7['h0082e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00418] =  Ifcca41d795dde8a35d1654b9520c92e7['h00830] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00419] =  Ifcca41d795dde8a35d1654b9520c92e7['h00832] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00834] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00836] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00838] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0083a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0083c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0041f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0083e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00420] =  Ifcca41d795dde8a35d1654b9520c92e7['h00840] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00421] =  Ifcca41d795dde8a35d1654b9520c92e7['h00842] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00422] =  Ifcca41d795dde8a35d1654b9520c92e7['h00844] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00423] =  Ifcca41d795dde8a35d1654b9520c92e7['h00846] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00424] =  Ifcca41d795dde8a35d1654b9520c92e7['h00848] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00425] =  Ifcca41d795dde8a35d1654b9520c92e7['h0084a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00426] =  Ifcca41d795dde8a35d1654b9520c92e7['h0084c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00427] =  Ifcca41d795dde8a35d1654b9520c92e7['h0084e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00428] =  Ifcca41d795dde8a35d1654b9520c92e7['h00850] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00429] =  Ifcca41d795dde8a35d1654b9520c92e7['h00852] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00854] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00856] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00858] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0085a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0085c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0042f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0085e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00430] =  Ifcca41d795dde8a35d1654b9520c92e7['h00860] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00431] =  Ifcca41d795dde8a35d1654b9520c92e7['h00862] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00432] =  Ifcca41d795dde8a35d1654b9520c92e7['h00864] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00433] =  Ifcca41d795dde8a35d1654b9520c92e7['h00866] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00434] =  Ifcca41d795dde8a35d1654b9520c92e7['h00868] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00435] =  Ifcca41d795dde8a35d1654b9520c92e7['h0086a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00436] =  Ifcca41d795dde8a35d1654b9520c92e7['h0086c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00437] =  Ifcca41d795dde8a35d1654b9520c92e7['h0086e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00438] =  Ifcca41d795dde8a35d1654b9520c92e7['h00870] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00439] =  Ifcca41d795dde8a35d1654b9520c92e7['h00872] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00874] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00876] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00878] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0087a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0087c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0043f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0087e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00440] =  Ifcca41d795dde8a35d1654b9520c92e7['h00880] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00441] =  Ifcca41d795dde8a35d1654b9520c92e7['h00882] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00442] =  Ifcca41d795dde8a35d1654b9520c92e7['h00884] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00443] =  Ifcca41d795dde8a35d1654b9520c92e7['h00886] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00444] =  Ifcca41d795dde8a35d1654b9520c92e7['h00888] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00445] =  Ifcca41d795dde8a35d1654b9520c92e7['h0088a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00446] =  Ifcca41d795dde8a35d1654b9520c92e7['h0088c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00447] =  Ifcca41d795dde8a35d1654b9520c92e7['h0088e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00448] =  Ifcca41d795dde8a35d1654b9520c92e7['h00890] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00449] =  Ifcca41d795dde8a35d1654b9520c92e7['h00892] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00894] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00896] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00898] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0089a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0089c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0044f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0089e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00450] =  Ifcca41d795dde8a35d1654b9520c92e7['h008a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00451] =  Ifcca41d795dde8a35d1654b9520c92e7['h008a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00452] =  Ifcca41d795dde8a35d1654b9520c92e7['h008a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00453] =  Ifcca41d795dde8a35d1654b9520c92e7['h008a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00454] =  Ifcca41d795dde8a35d1654b9520c92e7['h008a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00455] =  Ifcca41d795dde8a35d1654b9520c92e7['h008aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00456] =  Ifcca41d795dde8a35d1654b9520c92e7['h008ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00457] =  Ifcca41d795dde8a35d1654b9520c92e7['h008ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00458] =  Ifcca41d795dde8a35d1654b9520c92e7['h008b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00459] =  Ifcca41d795dde8a35d1654b9520c92e7['h008b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045a] =  Ifcca41d795dde8a35d1654b9520c92e7['h008b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045b] =  Ifcca41d795dde8a35d1654b9520c92e7['h008b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045c] =  Ifcca41d795dde8a35d1654b9520c92e7['h008b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045d] =  Ifcca41d795dde8a35d1654b9520c92e7['h008ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045e] =  Ifcca41d795dde8a35d1654b9520c92e7['h008bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0045f] =  Ifcca41d795dde8a35d1654b9520c92e7['h008be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00460] =  Ifcca41d795dde8a35d1654b9520c92e7['h008c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00461] =  Ifcca41d795dde8a35d1654b9520c92e7['h008c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00462] =  Ifcca41d795dde8a35d1654b9520c92e7['h008c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00463] =  Ifcca41d795dde8a35d1654b9520c92e7['h008c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00464] =  Ifcca41d795dde8a35d1654b9520c92e7['h008c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00465] =  Ifcca41d795dde8a35d1654b9520c92e7['h008ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00466] =  Ifcca41d795dde8a35d1654b9520c92e7['h008cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00467] =  Ifcca41d795dde8a35d1654b9520c92e7['h008ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00468] =  Ifcca41d795dde8a35d1654b9520c92e7['h008d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00469] =  Ifcca41d795dde8a35d1654b9520c92e7['h008d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046a] =  Ifcca41d795dde8a35d1654b9520c92e7['h008d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046b] =  Ifcca41d795dde8a35d1654b9520c92e7['h008d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046c] =  Ifcca41d795dde8a35d1654b9520c92e7['h008d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046d] =  Ifcca41d795dde8a35d1654b9520c92e7['h008da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046e] =  Ifcca41d795dde8a35d1654b9520c92e7['h008dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0046f] =  Ifcca41d795dde8a35d1654b9520c92e7['h008de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00470] =  Ifcca41d795dde8a35d1654b9520c92e7['h008e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00471] =  Ifcca41d795dde8a35d1654b9520c92e7['h008e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00472] =  Ifcca41d795dde8a35d1654b9520c92e7['h008e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00473] =  Ifcca41d795dde8a35d1654b9520c92e7['h008e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00474] =  Ifcca41d795dde8a35d1654b9520c92e7['h008e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00475] =  Ifcca41d795dde8a35d1654b9520c92e7['h008ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00476] =  Ifcca41d795dde8a35d1654b9520c92e7['h008ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00477] =  Ifcca41d795dde8a35d1654b9520c92e7['h008ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00478] =  Ifcca41d795dde8a35d1654b9520c92e7['h008f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00479] =  Ifcca41d795dde8a35d1654b9520c92e7['h008f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047a] =  Ifcca41d795dde8a35d1654b9520c92e7['h008f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047b] =  Ifcca41d795dde8a35d1654b9520c92e7['h008f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047c] =  Ifcca41d795dde8a35d1654b9520c92e7['h008f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047d] =  Ifcca41d795dde8a35d1654b9520c92e7['h008fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047e] =  Ifcca41d795dde8a35d1654b9520c92e7['h008fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0047f] =  Ifcca41d795dde8a35d1654b9520c92e7['h008fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00480] =  Ifcca41d795dde8a35d1654b9520c92e7['h00900] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00481] =  Ifcca41d795dde8a35d1654b9520c92e7['h00902] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00482] =  Ifcca41d795dde8a35d1654b9520c92e7['h00904] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00483] =  Ifcca41d795dde8a35d1654b9520c92e7['h00906] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00484] =  Ifcca41d795dde8a35d1654b9520c92e7['h00908] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00485] =  Ifcca41d795dde8a35d1654b9520c92e7['h0090a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00486] =  Ifcca41d795dde8a35d1654b9520c92e7['h0090c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00487] =  Ifcca41d795dde8a35d1654b9520c92e7['h0090e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00488] =  Ifcca41d795dde8a35d1654b9520c92e7['h00910] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00489] =  Ifcca41d795dde8a35d1654b9520c92e7['h00912] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00914] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00916] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00918] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0091a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0091c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0048f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0091e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00490] =  Ifcca41d795dde8a35d1654b9520c92e7['h00920] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00491] =  Ifcca41d795dde8a35d1654b9520c92e7['h00922] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00492] =  Ifcca41d795dde8a35d1654b9520c92e7['h00924] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00493] =  Ifcca41d795dde8a35d1654b9520c92e7['h00926] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00494] =  Ifcca41d795dde8a35d1654b9520c92e7['h00928] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00495] =  Ifcca41d795dde8a35d1654b9520c92e7['h0092a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00496] =  Ifcca41d795dde8a35d1654b9520c92e7['h0092c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00497] =  Ifcca41d795dde8a35d1654b9520c92e7['h0092e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00498] =  Ifcca41d795dde8a35d1654b9520c92e7['h00930] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00499] =  Ifcca41d795dde8a35d1654b9520c92e7['h00932] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00934] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00936] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00938] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0093a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0093c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0049f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0093e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00940] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00942] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00944] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00946] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00948] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0094a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0094c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0094e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00950] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00952] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00954] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h00956] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h00958] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0095a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0095c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004af] =  Ifcca41d795dde8a35d1654b9520c92e7['h0095e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00960] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00962] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00964] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00966] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00968] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0096a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0096c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0096e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00970] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00972] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h00974] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00976] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00978] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0097a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004be] =  Ifcca41d795dde8a35d1654b9520c92e7['h0097c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0097e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00980] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00982] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00984] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00986] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00988] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0098a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0098c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0098e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00990] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00992] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h00994] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00996] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00998] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0099a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0099c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0099e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h009a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h009a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h009a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h009a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h009a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h009aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h009ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h009ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h009b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h009b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004da] =  Ifcca41d795dde8a35d1654b9520c92e7['h009b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004db] =  Ifcca41d795dde8a35d1654b9520c92e7['h009b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h009b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h009ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004de] =  Ifcca41d795dde8a35d1654b9520c92e7['h009bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004df] =  Ifcca41d795dde8a35d1654b9520c92e7['h009be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h009c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h009c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h009c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h009c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h009c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h009ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h009cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h009ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h009d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h009d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h009d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h009d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h009d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h009da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h009dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h009de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h009e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h009e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h009e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h009e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h009e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h009ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h009ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h009ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h009f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h009f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h009f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h009f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h009f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h009fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h009fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h004ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h009fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00500] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00501] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00502] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00503] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00504] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00505] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00506] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00507] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00508] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00509] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0050f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00510] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00511] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00512] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00513] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00514] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00515] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00516] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00517] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00518] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00519] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0051f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00520] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00521] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00522] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00523] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00524] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00525] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00526] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00527] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00528] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00529] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0052f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00530] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00531] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00532] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00533] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00534] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00535] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00536] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00537] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00538] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00539] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0053f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00540] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00541] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00542] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00543] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00544] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00545] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00546] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00547] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00548] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00549] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0054f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00a9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00550] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aa0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00551] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aa2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00552] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aa4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00553] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aa6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00554] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aa8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00555] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aaa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00556] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00557] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00558] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ab0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00559] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ab2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ab4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ab6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ab8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00abc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0055f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00abe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00560] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ac0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00561] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ac2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00562] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ac4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00563] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ac6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00564] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ac8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00565] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00566] =  Ifcca41d795dde8a35d1654b9520c92e7['h00acc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00567] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ace] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00568] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ad0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00569] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ad2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ad4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ad6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ad8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ada] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00adc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0056f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ade] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00570] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ae0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00571] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ae2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00572] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ae4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00573] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ae6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00574] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ae8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00575] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00576] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00577] =  Ifcca41d795dde8a35d1654b9520c92e7['h00aee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00578] =  Ifcca41d795dde8a35d1654b9520c92e7['h00af0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00579] =  Ifcca41d795dde8a35d1654b9520c92e7['h00af2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00af4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00af6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00af8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00afa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00afc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0057f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00afe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00580] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00581] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00582] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00583] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00584] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00585] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00586] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00587] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00588] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00589] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0058f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00590] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00591] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00592] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00593] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00594] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00595] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00596] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00597] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00598] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00599] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0059f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005af] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005be] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h00b9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ba0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ba2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ba4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ba6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ba8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00baa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bb0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bb2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005da] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bb4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005db] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bb6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bb8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005de] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bbc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005df] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bbe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bc0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bc2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bc4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bc6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bc8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bcc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bd0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bd2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bd4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bd6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bd8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bdc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bde] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00be0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00be2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00be4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00be6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00be8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bf0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bf2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bf4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bf6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bf8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bfa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bfc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h005ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h00bfe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00600] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00601] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00602] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00603] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00604] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00605] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00606] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00607] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00608] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00609] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0060f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00610] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00611] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00612] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00613] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00614] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00615] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00616] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00617] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00618] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00619] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0061f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00620] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00621] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00622] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00623] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00624] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00625] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00626] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00627] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00628] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00629] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0062f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00630] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00631] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00632] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00633] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00634] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00635] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00636] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00637] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00638] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00639] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0063f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00640] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00641] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00642] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00643] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00644] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00645] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00646] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00647] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00648] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00649] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0064f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00c9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00650] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ca0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00651] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ca2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00652] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ca4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00653] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ca6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00654] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ca8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00655] =  Ifcca41d795dde8a35d1654b9520c92e7['h00caa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00656] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00657] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00658] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cb0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00659] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cb2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cb4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cb6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cb8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cbc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0065f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cbe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00660] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cc0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00661] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cc2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00662] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cc4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00663] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cc6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00664] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cc8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00665] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00666] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ccc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00667] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00668] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cd0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00669] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cd2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cd4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cd6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cd8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cdc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0066f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cde] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00670] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ce0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00671] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ce2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00672] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ce4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00673] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ce6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00674] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ce8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00675] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00676] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00677] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00678] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cf0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00679] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cf2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cf4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cf6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cf8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cfa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cfc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0067f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00cfe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00680] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00681] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00682] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00683] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00684] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00685] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00686] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00687] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00688] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00689] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0068f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00690] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00691] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00692] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00693] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00694] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00695] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00696] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00697] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00698] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00699] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0069f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006af] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006be] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h00d9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00da0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00da2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00da4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00da6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00da8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00daa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00db0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00db2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006da] =  Ifcca41d795dde8a35d1654b9520c92e7['h00db4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006db] =  Ifcca41d795dde8a35d1654b9520c92e7['h00db6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00db8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006de] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dbc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006df] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dbe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dc0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dc2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dc4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dc6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dc8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dcc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dd0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dd2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dd4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dd6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dd8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ddc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dde] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00de0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00de2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00de4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00de6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00de8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00df0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00df2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00df4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00df6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00df8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dfa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dfc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h006ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h00dfe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00700] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00701] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00702] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00703] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00704] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00705] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00706] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00707] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00708] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00709] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0070f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00710] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00711] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00712] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00713] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00714] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00715] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00716] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00717] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00718] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00719] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0071f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00720] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00721] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00722] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00723] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00724] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00725] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00726] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00727] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00728] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00729] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0072f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00730] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00731] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00732] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00733] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00734] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00735] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00736] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00737] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00738] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00739] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0073f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00740] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00741] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00742] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00743] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00744] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00745] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00746] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00747] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00748] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00749] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0074f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00e9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00750] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ea0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00751] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ea2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00752] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ea4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00753] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ea6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00754] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ea8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00755] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eaa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00756] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00757] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00758] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eb0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00759] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eb2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eb4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eb6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eb8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ebc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0075f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ebe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00760] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ec0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00761] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ec2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00762] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ec4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00763] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ec6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00764] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ec8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00765] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00766] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ecc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00767] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ece] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00768] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ed0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00769] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ed2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ed4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ed6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ed8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00edc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0076f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ede] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00770] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ee0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00771] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ee2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00772] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ee4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00773] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ee6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00774] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ee8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00775] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00776] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00777] =  Ifcca41d795dde8a35d1654b9520c92e7['h00eee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00778] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ef0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00779] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ef2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ef4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ef6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ef8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00efa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00efc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0077f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00efe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00780] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00781] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00782] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00783] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00784] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00785] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00786] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00787] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00788] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00789] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0078f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00790] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00791] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00792] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00793] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00794] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00795] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00796] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00797] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00798] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00799] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079a] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079b] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079c] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079d] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079e] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0079f] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007af] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007be] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h00f9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fa0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fa2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fa4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fa6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fa8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00faa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fb0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fb2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007da] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fb4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007db] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fb6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fb8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007de] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fbc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007df] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fbe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fc0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fc2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fc4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fc6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fc8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fcc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fd0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fd2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fd4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fd6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fd8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fdc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fde] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fe0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fe2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fe4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fe6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fe8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h00fee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ff0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ff2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ff4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ff6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ff8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ffa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ffc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h007ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h00ffe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00800] =  Ifcca41d795dde8a35d1654b9520c92e7['h01000] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00801] =  Ifcca41d795dde8a35d1654b9520c92e7['h01002] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00802] =  Ifcca41d795dde8a35d1654b9520c92e7['h01004] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00803] =  Ifcca41d795dde8a35d1654b9520c92e7['h01006] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00804] =  Ifcca41d795dde8a35d1654b9520c92e7['h01008] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00805] =  Ifcca41d795dde8a35d1654b9520c92e7['h0100a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00806] =  Ifcca41d795dde8a35d1654b9520c92e7['h0100c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00807] =  Ifcca41d795dde8a35d1654b9520c92e7['h0100e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00808] =  Ifcca41d795dde8a35d1654b9520c92e7['h01010] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00809] =  Ifcca41d795dde8a35d1654b9520c92e7['h01012] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01014] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01016] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01018] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0101a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0101c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0080f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0101e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00810] =  Ifcca41d795dde8a35d1654b9520c92e7['h01020] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00811] =  Ifcca41d795dde8a35d1654b9520c92e7['h01022] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00812] =  Ifcca41d795dde8a35d1654b9520c92e7['h01024] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00813] =  Ifcca41d795dde8a35d1654b9520c92e7['h01026] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00814] =  Ifcca41d795dde8a35d1654b9520c92e7['h01028] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00815] =  Ifcca41d795dde8a35d1654b9520c92e7['h0102a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00816] =  Ifcca41d795dde8a35d1654b9520c92e7['h0102c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00817] =  Ifcca41d795dde8a35d1654b9520c92e7['h0102e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00818] =  Ifcca41d795dde8a35d1654b9520c92e7['h01030] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00819] =  Ifcca41d795dde8a35d1654b9520c92e7['h01032] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01034] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01036] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01038] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0103a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0103c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0081f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0103e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00820] =  Ifcca41d795dde8a35d1654b9520c92e7['h01040] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00821] =  Ifcca41d795dde8a35d1654b9520c92e7['h01042] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00822] =  Ifcca41d795dde8a35d1654b9520c92e7['h01044] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00823] =  Ifcca41d795dde8a35d1654b9520c92e7['h01046] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00824] =  Ifcca41d795dde8a35d1654b9520c92e7['h01048] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00825] =  Ifcca41d795dde8a35d1654b9520c92e7['h0104a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00826] =  Ifcca41d795dde8a35d1654b9520c92e7['h0104c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00827] =  Ifcca41d795dde8a35d1654b9520c92e7['h0104e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00828] =  Ifcca41d795dde8a35d1654b9520c92e7['h01050] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00829] =  Ifcca41d795dde8a35d1654b9520c92e7['h01052] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01054] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01056] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01058] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0105a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0105c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0082f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0105e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00830] =  Ifcca41d795dde8a35d1654b9520c92e7['h01060] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00831] =  Ifcca41d795dde8a35d1654b9520c92e7['h01062] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00832] =  Ifcca41d795dde8a35d1654b9520c92e7['h01064] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00833] =  Ifcca41d795dde8a35d1654b9520c92e7['h01066] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00834] =  Ifcca41d795dde8a35d1654b9520c92e7['h01068] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00835] =  Ifcca41d795dde8a35d1654b9520c92e7['h0106a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00836] =  Ifcca41d795dde8a35d1654b9520c92e7['h0106c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00837] =  Ifcca41d795dde8a35d1654b9520c92e7['h0106e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00838] =  Ifcca41d795dde8a35d1654b9520c92e7['h01070] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00839] =  Ifcca41d795dde8a35d1654b9520c92e7['h01072] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01074] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01076] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01078] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0107a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0107c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0083f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0107e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00840] =  Ifcca41d795dde8a35d1654b9520c92e7['h01080] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00841] =  Ifcca41d795dde8a35d1654b9520c92e7['h01082] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00842] =  Ifcca41d795dde8a35d1654b9520c92e7['h01084] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00843] =  Ifcca41d795dde8a35d1654b9520c92e7['h01086] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00844] =  Ifcca41d795dde8a35d1654b9520c92e7['h01088] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00845] =  Ifcca41d795dde8a35d1654b9520c92e7['h0108a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00846] =  Ifcca41d795dde8a35d1654b9520c92e7['h0108c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00847] =  Ifcca41d795dde8a35d1654b9520c92e7['h0108e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00848] =  Ifcca41d795dde8a35d1654b9520c92e7['h01090] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00849] =  Ifcca41d795dde8a35d1654b9520c92e7['h01092] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01094] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01096] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01098] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0109a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0109c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0084f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0109e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00850] =  Ifcca41d795dde8a35d1654b9520c92e7['h010a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00851] =  Ifcca41d795dde8a35d1654b9520c92e7['h010a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00852] =  Ifcca41d795dde8a35d1654b9520c92e7['h010a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00853] =  Ifcca41d795dde8a35d1654b9520c92e7['h010a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00854] =  Ifcca41d795dde8a35d1654b9520c92e7['h010a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00855] =  Ifcca41d795dde8a35d1654b9520c92e7['h010aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00856] =  Ifcca41d795dde8a35d1654b9520c92e7['h010ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00857] =  Ifcca41d795dde8a35d1654b9520c92e7['h010ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00858] =  Ifcca41d795dde8a35d1654b9520c92e7['h010b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00859] =  Ifcca41d795dde8a35d1654b9520c92e7['h010b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085a] =  Ifcca41d795dde8a35d1654b9520c92e7['h010b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085b] =  Ifcca41d795dde8a35d1654b9520c92e7['h010b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085c] =  Ifcca41d795dde8a35d1654b9520c92e7['h010b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085d] =  Ifcca41d795dde8a35d1654b9520c92e7['h010ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085e] =  Ifcca41d795dde8a35d1654b9520c92e7['h010bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0085f] =  Ifcca41d795dde8a35d1654b9520c92e7['h010be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00860] =  Ifcca41d795dde8a35d1654b9520c92e7['h010c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00861] =  Ifcca41d795dde8a35d1654b9520c92e7['h010c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00862] =  Ifcca41d795dde8a35d1654b9520c92e7['h010c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00863] =  Ifcca41d795dde8a35d1654b9520c92e7['h010c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00864] =  Ifcca41d795dde8a35d1654b9520c92e7['h010c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00865] =  Ifcca41d795dde8a35d1654b9520c92e7['h010ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00866] =  Ifcca41d795dde8a35d1654b9520c92e7['h010cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00867] =  Ifcca41d795dde8a35d1654b9520c92e7['h010ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00868] =  Ifcca41d795dde8a35d1654b9520c92e7['h010d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00869] =  Ifcca41d795dde8a35d1654b9520c92e7['h010d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086a] =  Ifcca41d795dde8a35d1654b9520c92e7['h010d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086b] =  Ifcca41d795dde8a35d1654b9520c92e7['h010d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086c] =  Ifcca41d795dde8a35d1654b9520c92e7['h010d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086d] =  Ifcca41d795dde8a35d1654b9520c92e7['h010da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086e] =  Ifcca41d795dde8a35d1654b9520c92e7['h010dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0086f] =  Ifcca41d795dde8a35d1654b9520c92e7['h010de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00870] =  Ifcca41d795dde8a35d1654b9520c92e7['h010e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00871] =  Ifcca41d795dde8a35d1654b9520c92e7['h010e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00872] =  Ifcca41d795dde8a35d1654b9520c92e7['h010e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00873] =  Ifcca41d795dde8a35d1654b9520c92e7['h010e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00874] =  Ifcca41d795dde8a35d1654b9520c92e7['h010e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00875] =  Ifcca41d795dde8a35d1654b9520c92e7['h010ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00876] =  Ifcca41d795dde8a35d1654b9520c92e7['h010ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00877] =  Ifcca41d795dde8a35d1654b9520c92e7['h010ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00878] =  Ifcca41d795dde8a35d1654b9520c92e7['h010f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00879] =  Ifcca41d795dde8a35d1654b9520c92e7['h010f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087a] =  Ifcca41d795dde8a35d1654b9520c92e7['h010f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087b] =  Ifcca41d795dde8a35d1654b9520c92e7['h010f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087c] =  Ifcca41d795dde8a35d1654b9520c92e7['h010f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087d] =  Ifcca41d795dde8a35d1654b9520c92e7['h010fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087e] =  Ifcca41d795dde8a35d1654b9520c92e7['h010fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0087f] =  Ifcca41d795dde8a35d1654b9520c92e7['h010fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00880] =  Ifcca41d795dde8a35d1654b9520c92e7['h01100] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00881] =  Ifcca41d795dde8a35d1654b9520c92e7['h01102] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00882] =  Ifcca41d795dde8a35d1654b9520c92e7['h01104] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00883] =  Ifcca41d795dde8a35d1654b9520c92e7['h01106] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00884] =  Ifcca41d795dde8a35d1654b9520c92e7['h01108] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00885] =  Ifcca41d795dde8a35d1654b9520c92e7['h0110a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00886] =  Ifcca41d795dde8a35d1654b9520c92e7['h0110c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00887] =  Ifcca41d795dde8a35d1654b9520c92e7['h0110e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00888] =  Ifcca41d795dde8a35d1654b9520c92e7['h01110] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00889] =  Ifcca41d795dde8a35d1654b9520c92e7['h01112] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01114] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01116] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01118] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0111a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0111c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0088f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0111e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00890] =  Ifcca41d795dde8a35d1654b9520c92e7['h01120] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00891] =  Ifcca41d795dde8a35d1654b9520c92e7['h01122] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00892] =  Ifcca41d795dde8a35d1654b9520c92e7['h01124] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00893] =  Ifcca41d795dde8a35d1654b9520c92e7['h01126] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00894] =  Ifcca41d795dde8a35d1654b9520c92e7['h01128] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00895] =  Ifcca41d795dde8a35d1654b9520c92e7['h0112a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00896] =  Ifcca41d795dde8a35d1654b9520c92e7['h0112c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00897] =  Ifcca41d795dde8a35d1654b9520c92e7['h0112e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00898] =  Ifcca41d795dde8a35d1654b9520c92e7['h01130] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00899] =  Ifcca41d795dde8a35d1654b9520c92e7['h01132] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01134] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01136] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01138] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0113a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0113c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0089f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0113e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01140] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01142] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01144] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01146] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01148] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0114a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0114c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0114e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01150] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01152] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01154] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h01156] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h01158] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0115a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0115c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008af] =  Ifcca41d795dde8a35d1654b9520c92e7['h0115e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01160] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01162] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01164] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01166] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01168] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0116a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0116c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0116e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01170] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01172] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h01174] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01176] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01178] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0117a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008be] =  Ifcca41d795dde8a35d1654b9520c92e7['h0117c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0117e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01180] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01182] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01184] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01186] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01188] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0118a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0118c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0118e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01190] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01192] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h01194] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01196] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01198] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0119a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0119c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0119e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h011a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h011a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h011a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h011a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h011a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h011aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h011ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h011ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h011b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h011b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008da] =  Ifcca41d795dde8a35d1654b9520c92e7['h011b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008db] =  Ifcca41d795dde8a35d1654b9520c92e7['h011b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h011b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h011ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008de] =  Ifcca41d795dde8a35d1654b9520c92e7['h011bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008df] =  Ifcca41d795dde8a35d1654b9520c92e7['h011be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h011c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h011c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h011c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h011c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h011c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h011ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h011cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h011ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h011d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h011d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h011d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h011d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h011d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h011da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h011dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h011de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h011e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h011e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h011e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h011e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h011e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h011ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h011ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h011ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h011f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h011f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h011f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h011f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h011f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h011fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h011fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h008ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h011fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00900] =  Ifcca41d795dde8a35d1654b9520c92e7['h01200] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00901] =  Ifcca41d795dde8a35d1654b9520c92e7['h01202] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00902] =  Ifcca41d795dde8a35d1654b9520c92e7['h01204] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00903] =  Ifcca41d795dde8a35d1654b9520c92e7['h01206] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00904] =  Ifcca41d795dde8a35d1654b9520c92e7['h01208] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00905] =  Ifcca41d795dde8a35d1654b9520c92e7['h0120a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00906] =  Ifcca41d795dde8a35d1654b9520c92e7['h0120c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00907] =  Ifcca41d795dde8a35d1654b9520c92e7['h0120e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00908] =  Ifcca41d795dde8a35d1654b9520c92e7['h01210] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00909] =  Ifcca41d795dde8a35d1654b9520c92e7['h01212] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01214] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01216] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01218] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0121a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0121c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0090f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0121e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00910] =  Ifcca41d795dde8a35d1654b9520c92e7['h01220] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00911] =  Ifcca41d795dde8a35d1654b9520c92e7['h01222] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00912] =  Ifcca41d795dde8a35d1654b9520c92e7['h01224] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00913] =  Ifcca41d795dde8a35d1654b9520c92e7['h01226] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00914] =  Ifcca41d795dde8a35d1654b9520c92e7['h01228] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00915] =  Ifcca41d795dde8a35d1654b9520c92e7['h0122a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00916] =  Ifcca41d795dde8a35d1654b9520c92e7['h0122c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00917] =  Ifcca41d795dde8a35d1654b9520c92e7['h0122e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00918] =  Ifcca41d795dde8a35d1654b9520c92e7['h01230] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00919] =  Ifcca41d795dde8a35d1654b9520c92e7['h01232] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01234] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01236] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01238] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0123a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0123c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0091f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0123e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00920] =  Ifcca41d795dde8a35d1654b9520c92e7['h01240] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00921] =  Ifcca41d795dde8a35d1654b9520c92e7['h01242] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00922] =  Ifcca41d795dde8a35d1654b9520c92e7['h01244] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00923] =  Ifcca41d795dde8a35d1654b9520c92e7['h01246] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00924] =  Ifcca41d795dde8a35d1654b9520c92e7['h01248] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00925] =  Ifcca41d795dde8a35d1654b9520c92e7['h0124a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00926] =  Ifcca41d795dde8a35d1654b9520c92e7['h0124c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00927] =  Ifcca41d795dde8a35d1654b9520c92e7['h0124e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00928] =  Ifcca41d795dde8a35d1654b9520c92e7['h01250] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00929] =  Ifcca41d795dde8a35d1654b9520c92e7['h01252] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01254] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01256] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01258] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0125a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0125c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0092f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0125e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00930] =  Ifcca41d795dde8a35d1654b9520c92e7['h01260] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00931] =  Ifcca41d795dde8a35d1654b9520c92e7['h01262] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00932] =  Ifcca41d795dde8a35d1654b9520c92e7['h01264] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00933] =  Ifcca41d795dde8a35d1654b9520c92e7['h01266] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00934] =  Ifcca41d795dde8a35d1654b9520c92e7['h01268] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00935] =  Ifcca41d795dde8a35d1654b9520c92e7['h0126a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00936] =  Ifcca41d795dde8a35d1654b9520c92e7['h0126c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00937] =  Ifcca41d795dde8a35d1654b9520c92e7['h0126e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00938] =  Ifcca41d795dde8a35d1654b9520c92e7['h01270] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00939] =  Ifcca41d795dde8a35d1654b9520c92e7['h01272] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01274] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01276] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01278] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0127a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0127c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0093f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0127e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00940] =  Ifcca41d795dde8a35d1654b9520c92e7['h01280] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00941] =  Ifcca41d795dde8a35d1654b9520c92e7['h01282] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00942] =  Ifcca41d795dde8a35d1654b9520c92e7['h01284] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00943] =  Ifcca41d795dde8a35d1654b9520c92e7['h01286] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00944] =  Ifcca41d795dde8a35d1654b9520c92e7['h01288] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00945] =  Ifcca41d795dde8a35d1654b9520c92e7['h0128a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00946] =  Ifcca41d795dde8a35d1654b9520c92e7['h0128c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00947] =  Ifcca41d795dde8a35d1654b9520c92e7['h0128e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00948] =  Ifcca41d795dde8a35d1654b9520c92e7['h01290] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00949] =  Ifcca41d795dde8a35d1654b9520c92e7['h01292] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01294] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01296] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01298] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0129a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0129c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0094f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0129e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00950] =  Ifcca41d795dde8a35d1654b9520c92e7['h012a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00951] =  Ifcca41d795dde8a35d1654b9520c92e7['h012a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00952] =  Ifcca41d795dde8a35d1654b9520c92e7['h012a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00953] =  Ifcca41d795dde8a35d1654b9520c92e7['h012a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00954] =  Ifcca41d795dde8a35d1654b9520c92e7['h012a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00955] =  Ifcca41d795dde8a35d1654b9520c92e7['h012aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00956] =  Ifcca41d795dde8a35d1654b9520c92e7['h012ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00957] =  Ifcca41d795dde8a35d1654b9520c92e7['h012ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00958] =  Ifcca41d795dde8a35d1654b9520c92e7['h012b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00959] =  Ifcca41d795dde8a35d1654b9520c92e7['h012b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095a] =  Ifcca41d795dde8a35d1654b9520c92e7['h012b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095b] =  Ifcca41d795dde8a35d1654b9520c92e7['h012b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095c] =  Ifcca41d795dde8a35d1654b9520c92e7['h012b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095d] =  Ifcca41d795dde8a35d1654b9520c92e7['h012ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095e] =  Ifcca41d795dde8a35d1654b9520c92e7['h012bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0095f] =  Ifcca41d795dde8a35d1654b9520c92e7['h012be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00960] =  Ifcca41d795dde8a35d1654b9520c92e7['h012c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00961] =  Ifcca41d795dde8a35d1654b9520c92e7['h012c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00962] =  Ifcca41d795dde8a35d1654b9520c92e7['h012c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00963] =  Ifcca41d795dde8a35d1654b9520c92e7['h012c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00964] =  Ifcca41d795dde8a35d1654b9520c92e7['h012c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00965] =  Ifcca41d795dde8a35d1654b9520c92e7['h012ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00966] =  Ifcca41d795dde8a35d1654b9520c92e7['h012cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00967] =  Ifcca41d795dde8a35d1654b9520c92e7['h012ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00968] =  Ifcca41d795dde8a35d1654b9520c92e7['h012d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00969] =  Ifcca41d795dde8a35d1654b9520c92e7['h012d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096a] =  Ifcca41d795dde8a35d1654b9520c92e7['h012d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096b] =  Ifcca41d795dde8a35d1654b9520c92e7['h012d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096c] =  Ifcca41d795dde8a35d1654b9520c92e7['h012d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096d] =  Ifcca41d795dde8a35d1654b9520c92e7['h012da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096e] =  Ifcca41d795dde8a35d1654b9520c92e7['h012dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0096f] =  Ifcca41d795dde8a35d1654b9520c92e7['h012de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00970] =  Ifcca41d795dde8a35d1654b9520c92e7['h012e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00971] =  Ifcca41d795dde8a35d1654b9520c92e7['h012e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00972] =  Ifcca41d795dde8a35d1654b9520c92e7['h012e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00973] =  Ifcca41d795dde8a35d1654b9520c92e7['h012e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00974] =  Ifcca41d795dde8a35d1654b9520c92e7['h012e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00975] =  Ifcca41d795dde8a35d1654b9520c92e7['h012ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00976] =  Ifcca41d795dde8a35d1654b9520c92e7['h012ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00977] =  Ifcca41d795dde8a35d1654b9520c92e7['h012ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00978] =  Ifcca41d795dde8a35d1654b9520c92e7['h012f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00979] =  Ifcca41d795dde8a35d1654b9520c92e7['h012f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097a] =  Ifcca41d795dde8a35d1654b9520c92e7['h012f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097b] =  Ifcca41d795dde8a35d1654b9520c92e7['h012f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097c] =  Ifcca41d795dde8a35d1654b9520c92e7['h012f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097d] =  Ifcca41d795dde8a35d1654b9520c92e7['h012fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097e] =  Ifcca41d795dde8a35d1654b9520c92e7['h012fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0097f] =  Ifcca41d795dde8a35d1654b9520c92e7['h012fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00980] =  Ifcca41d795dde8a35d1654b9520c92e7['h01300] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00981] =  Ifcca41d795dde8a35d1654b9520c92e7['h01302] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00982] =  Ifcca41d795dde8a35d1654b9520c92e7['h01304] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00983] =  Ifcca41d795dde8a35d1654b9520c92e7['h01306] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00984] =  Ifcca41d795dde8a35d1654b9520c92e7['h01308] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00985] =  Ifcca41d795dde8a35d1654b9520c92e7['h0130a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00986] =  Ifcca41d795dde8a35d1654b9520c92e7['h0130c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00987] =  Ifcca41d795dde8a35d1654b9520c92e7['h0130e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00988] =  Ifcca41d795dde8a35d1654b9520c92e7['h01310] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00989] =  Ifcca41d795dde8a35d1654b9520c92e7['h01312] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01314] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01316] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01318] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0131a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0131c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0098f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0131e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00990] =  Ifcca41d795dde8a35d1654b9520c92e7['h01320] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00991] =  Ifcca41d795dde8a35d1654b9520c92e7['h01322] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00992] =  Ifcca41d795dde8a35d1654b9520c92e7['h01324] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00993] =  Ifcca41d795dde8a35d1654b9520c92e7['h01326] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00994] =  Ifcca41d795dde8a35d1654b9520c92e7['h01328] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00995] =  Ifcca41d795dde8a35d1654b9520c92e7['h0132a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00996] =  Ifcca41d795dde8a35d1654b9520c92e7['h0132c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00997] =  Ifcca41d795dde8a35d1654b9520c92e7['h0132e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00998] =  Ifcca41d795dde8a35d1654b9520c92e7['h01330] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00999] =  Ifcca41d795dde8a35d1654b9520c92e7['h01332] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01334] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01336] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01338] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0133a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0133c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h0099f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0133e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01340] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01342] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01344] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01346] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01348] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0134a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0134c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0134e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01350] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009a9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01352] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009aa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01354] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ab] =  Ifcca41d795dde8a35d1654b9520c92e7['h01356] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ac] =  Ifcca41d795dde8a35d1654b9520c92e7['h01358] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0135a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0135c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009af] =  Ifcca41d795dde8a35d1654b9520c92e7['h0135e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01360] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01362] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01364] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01366] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01368] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0136a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0136c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0136e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01370] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009b9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01372] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ba] =  Ifcca41d795dde8a35d1654b9520c92e7['h01374] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009bb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01376] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009bc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01378] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009bd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0137a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009be] =  Ifcca41d795dde8a35d1654b9520c92e7['h0137c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009bf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0137e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01380] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01382] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01384] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01386] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01388] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0138a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0138c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0138e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01390] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009c9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01392] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ca] =  Ifcca41d795dde8a35d1654b9520c92e7['h01394] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009cb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01396] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009cc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01398] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009cd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0139a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0139c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009cf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0139e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d0] =  Ifcca41d795dde8a35d1654b9520c92e7['h013a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d1] =  Ifcca41d795dde8a35d1654b9520c92e7['h013a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d2] =  Ifcca41d795dde8a35d1654b9520c92e7['h013a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d3] =  Ifcca41d795dde8a35d1654b9520c92e7['h013a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d4] =  Ifcca41d795dde8a35d1654b9520c92e7['h013a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d5] =  Ifcca41d795dde8a35d1654b9520c92e7['h013aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d6] =  Ifcca41d795dde8a35d1654b9520c92e7['h013ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d7] =  Ifcca41d795dde8a35d1654b9520c92e7['h013ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d8] =  Ifcca41d795dde8a35d1654b9520c92e7['h013b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009d9] =  Ifcca41d795dde8a35d1654b9520c92e7['h013b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009da] =  Ifcca41d795dde8a35d1654b9520c92e7['h013b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009db] =  Ifcca41d795dde8a35d1654b9520c92e7['h013b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009dc] =  Ifcca41d795dde8a35d1654b9520c92e7['h013b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009dd] =  Ifcca41d795dde8a35d1654b9520c92e7['h013ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009de] =  Ifcca41d795dde8a35d1654b9520c92e7['h013bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009df] =  Ifcca41d795dde8a35d1654b9520c92e7['h013be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e0] =  Ifcca41d795dde8a35d1654b9520c92e7['h013c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e1] =  Ifcca41d795dde8a35d1654b9520c92e7['h013c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e2] =  Ifcca41d795dde8a35d1654b9520c92e7['h013c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e3] =  Ifcca41d795dde8a35d1654b9520c92e7['h013c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e4] =  Ifcca41d795dde8a35d1654b9520c92e7['h013c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e5] =  Ifcca41d795dde8a35d1654b9520c92e7['h013ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e6] =  Ifcca41d795dde8a35d1654b9520c92e7['h013cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e7] =  Ifcca41d795dde8a35d1654b9520c92e7['h013ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e8] =  Ifcca41d795dde8a35d1654b9520c92e7['h013d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009e9] =  Ifcca41d795dde8a35d1654b9520c92e7['h013d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ea] =  Ifcca41d795dde8a35d1654b9520c92e7['h013d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009eb] =  Ifcca41d795dde8a35d1654b9520c92e7['h013d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ec] =  Ifcca41d795dde8a35d1654b9520c92e7['h013d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ed] =  Ifcca41d795dde8a35d1654b9520c92e7['h013da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ee] =  Ifcca41d795dde8a35d1654b9520c92e7['h013dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ef] =  Ifcca41d795dde8a35d1654b9520c92e7['h013de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f0] =  Ifcca41d795dde8a35d1654b9520c92e7['h013e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f1] =  Ifcca41d795dde8a35d1654b9520c92e7['h013e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f2] =  Ifcca41d795dde8a35d1654b9520c92e7['h013e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f3] =  Ifcca41d795dde8a35d1654b9520c92e7['h013e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f4] =  Ifcca41d795dde8a35d1654b9520c92e7['h013e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f5] =  Ifcca41d795dde8a35d1654b9520c92e7['h013ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f6] =  Ifcca41d795dde8a35d1654b9520c92e7['h013ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f7] =  Ifcca41d795dde8a35d1654b9520c92e7['h013ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f8] =  Ifcca41d795dde8a35d1654b9520c92e7['h013f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009f9] =  Ifcca41d795dde8a35d1654b9520c92e7['h013f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009fa] =  Ifcca41d795dde8a35d1654b9520c92e7['h013f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009fb] =  Ifcca41d795dde8a35d1654b9520c92e7['h013f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009fc] =  Ifcca41d795dde8a35d1654b9520c92e7['h013f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009fd] =  Ifcca41d795dde8a35d1654b9520c92e7['h013fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009fe] =  Ifcca41d795dde8a35d1654b9520c92e7['h013fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h009ff] =  Ifcca41d795dde8a35d1654b9520c92e7['h013fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a00] =  Ifcca41d795dde8a35d1654b9520c92e7['h01400] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a01] =  Ifcca41d795dde8a35d1654b9520c92e7['h01402] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a02] =  Ifcca41d795dde8a35d1654b9520c92e7['h01404] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a03] =  Ifcca41d795dde8a35d1654b9520c92e7['h01406] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a04] =  Ifcca41d795dde8a35d1654b9520c92e7['h01408] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a05] =  Ifcca41d795dde8a35d1654b9520c92e7['h0140a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a06] =  Ifcca41d795dde8a35d1654b9520c92e7['h0140c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a07] =  Ifcca41d795dde8a35d1654b9520c92e7['h0140e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a08] =  Ifcca41d795dde8a35d1654b9520c92e7['h01410] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a09] =  Ifcca41d795dde8a35d1654b9520c92e7['h01412] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01414] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01416] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01418] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0141a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0141c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a0f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0141e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a10] =  Ifcca41d795dde8a35d1654b9520c92e7['h01420] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a11] =  Ifcca41d795dde8a35d1654b9520c92e7['h01422] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a12] =  Ifcca41d795dde8a35d1654b9520c92e7['h01424] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a13] =  Ifcca41d795dde8a35d1654b9520c92e7['h01426] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a14] =  Ifcca41d795dde8a35d1654b9520c92e7['h01428] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a15] =  Ifcca41d795dde8a35d1654b9520c92e7['h0142a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a16] =  Ifcca41d795dde8a35d1654b9520c92e7['h0142c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a17] =  Ifcca41d795dde8a35d1654b9520c92e7['h0142e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a18] =  Ifcca41d795dde8a35d1654b9520c92e7['h01430] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a19] =  Ifcca41d795dde8a35d1654b9520c92e7['h01432] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01434] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01436] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01438] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0143a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0143c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a1f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0143e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a20] =  Ifcca41d795dde8a35d1654b9520c92e7['h01440] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a21] =  Ifcca41d795dde8a35d1654b9520c92e7['h01442] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a22] =  Ifcca41d795dde8a35d1654b9520c92e7['h01444] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a23] =  Ifcca41d795dde8a35d1654b9520c92e7['h01446] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a24] =  Ifcca41d795dde8a35d1654b9520c92e7['h01448] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a25] =  Ifcca41d795dde8a35d1654b9520c92e7['h0144a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a26] =  Ifcca41d795dde8a35d1654b9520c92e7['h0144c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a27] =  Ifcca41d795dde8a35d1654b9520c92e7['h0144e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a28] =  Ifcca41d795dde8a35d1654b9520c92e7['h01450] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a29] =  Ifcca41d795dde8a35d1654b9520c92e7['h01452] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01454] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01456] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01458] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0145a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0145c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a2f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0145e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a30] =  Ifcca41d795dde8a35d1654b9520c92e7['h01460] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a31] =  Ifcca41d795dde8a35d1654b9520c92e7['h01462] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a32] =  Ifcca41d795dde8a35d1654b9520c92e7['h01464] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a33] =  Ifcca41d795dde8a35d1654b9520c92e7['h01466] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a34] =  Ifcca41d795dde8a35d1654b9520c92e7['h01468] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a35] =  Ifcca41d795dde8a35d1654b9520c92e7['h0146a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a36] =  Ifcca41d795dde8a35d1654b9520c92e7['h0146c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a37] =  Ifcca41d795dde8a35d1654b9520c92e7['h0146e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a38] =  Ifcca41d795dde8a35d1654b9520c92e7['h01470] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a39] =  Ifcca41d795dde8a35d1654b9520c92e7['h01472] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01474] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01476] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01478] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0147a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0147c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a3f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0147e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a40] =  Ifcca41d795dde8a35d1654b9520c92e7['h01480] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a41] =  Ifcca41d795dde8a35d1654b9520c92e7['h01482] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a42] =  Ifcca41d795dde8a35d1654b9520c92e7['h01484] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a43] =  Ifcca41d795dde8a35d1654b9520c92e7['h01486] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a44] =  Ifcca41d795dde8a35d1654b9520c92e7['h01488] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a45] =  Ifcca41d795dde8a35d1654b9520c92e7['h0148a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a46] =  Ifcca41d795dde8a35d1654b9520c92e7['h0148c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a47] =  Ifcca41d795dde8a35d1654b9520c92e7['h0148e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a48] =  Ifcca41d795dde8a35d1654b9520c92e7['h01490] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a49] =  Ifcca41d795dde8a35d1654b9520c92e7['h01492] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01494] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01496] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01498] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0149a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0149c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a4f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0149e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a50] =  Ifcca41d795dde8a35d1654b9520c92e7['h014a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a51] =  Ifcca41d795dde8a35d1654b9520c92e7['h014a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a52] =  Ifcca41d795dde8a35d1654b9520c92e7['h014a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a53] =  Ifcca41d795dde8a35d1654b9520c92e7['h014a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a54] =  Ifcca41d795dde8a35d1654b9520c92e7['h014a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a55] =  Ifcca41d795dde8a35d1654b9520c92e7['h014aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a56] =  Ifcca41d795dde8a35d1654b9520c92e7['h014ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a57] =  Ifcca41d795dde8a35d1654b9520c92e7['h014ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a58] =  Ifcca41d795dde8a35d1654b9520c92e7['h014b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a59] =  Ifcca41d795dde8a35d1654b9520c92e7['h014b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5a] =  Ifcca41d795dde8a35d1654b9520c92e7['h014b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5b] =  Ifcca41d795dde8a35d1654b9520c92e7['h014b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5c] =  Ifcca41d795dde8a35d1654b9520c92e7['h014b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5d] =  Ifcca41d795dde8a35d1654b9520c92e7['h014ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5e] =  Ifcca41d795dde8a35d1654b9520c92e7['h014bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a5f] =  Ifcca41d795dde8a35d1654b9520c92e7['h014be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a60] =  Ifcca41d795dde8a35d1654b9520c92e7['h014c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a61] =  Ifcca41d795dde8a35d1654b9520c92e7['h014c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a62] =  Ifcca41d795dde8a35d1654b9520c92e7['h014c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a63] =  Ifcca41d795dde8a35d1654b9520c92e7['h014c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a64] =  Ifcca41d795dde8a35d1654b9520c92e7['h014c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a65] =  Ifcca41d795dde8a35d1654b9520c92e7['h014ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a66] =  Ifcca41d795dde8a35d1654b9520c92e7['h014cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a67] =  Ifcca41d795dde8a35d1654b9520c92e7['h014ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a68] =  Ifcca41d795dde8a35d1654b9520c92e7['h014d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a69] =  Ifcca41d795dde8a35d1654b9520c92e7['h014d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6a] =  Ifcca41d795dde8a35d1654b9520c92e7['h014d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6b] =  Ifcca41d795dde8a35d1654b9520c92e7['h014d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6c] =  Ifcca41d795dde8a35d1654b9520c92e7['h014d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6d] =  Ifcca41d795dde8a35d1654b9520c92e7['h014da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6e] =  Ifcca41d795dde8a35d1654b9520c92e7['h014dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a6f] =  Ifcca41d795dde8a35d1654b9520c92e7['h014de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a70] =  Ifcca41d795dde8a35d1654b9520c92e7['h014e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a71] =  Ifcca41d795dde8a35d1654b9520c92e7['h014e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a72] =  Ifcca41d795dde8a35d1654b9520c92e7['h014e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a73] =  Ifcca41d795dde8a35d1654b9520c92e7['h014e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a74] =  Ifcca41d795dde8a35d1654b9520c92e7['h014e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a75] =  Ifcca41d795dde8a35d1654b9520c92e7['h014ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a76] =  Ifcca41d795dde8a35d1654b9520c92e7['h014ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a77] =  Ifcca41d795dde8a35d1654b9520c92e7['h014ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a78] =  Ifcca41d795dde8a35d1654b9520c92e7['h014f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a79] =  Ifcca41d795dde8a35d1654b9520c92e7['h014f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7a] =  Ifcca41d795dde8a35d1654b9520c92e7['h014f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7b] =  Ifcca41d795dde8a35d1654b9520c92e7['h014f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7c] =  Ifcca41d795dde8a35d1654b9520c92e7['h014f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7d] =  Ifcca41d795dde8a35d1654b9520c92e7['h014fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7e] =  Ifcca41d795dde8a35d1654b9520c92e7['h014fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a7f] =  Ifcca41d795dde8a35d1654b9520c92e7['h014fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a80] =  Ifcca41d795dde8a35d1654b9520c92e7['h01500] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a81] =  Ifcca41d795dde8a35d1654b9520c92e7['h01502] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a82] =  Ifcca41d795dde8a35d1654b9520c92e7['h01504] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a83] =  Ifcca41d795dde8a35d1654b9520c92e7['h01506] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a84] =  Ifcca41d795dde8a35d1654b9520c92e7['h01508] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a85] =  Ifcca41d795dde8a35d1654b9520c92e7['h0150a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a86] =  Ifcca41d795dde8a35d1654b9520c92e7['h0150c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a87] =  Ifcca41d795dde8a35d1654b9520c92e7['h0150e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a88] =  Ifcca41d795dde8a35d1654b9520c92e7['h01510] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a89] =  Ifcca41d795dde8a35d1654b9520c92e7['h01512] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01514] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01516] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01518] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0151a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0151c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a8f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0151e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a90] =  Ifcca41d795dde8a35d1654b9520c92e7['h01520] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a91] =  Ifcca41d795dde8a35d1654b9520c92e7['h01522] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a92] =  Ifcca41d795dde8a35d1654b9520c92e7['h01524] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a93] =  Ifcca41d795dde8a35d1654b9520c92e7['h01526] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a94] =  Ifcca41d795dde8a35d1654b9520c92e7['h01528] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a95] =  Ifcca41d795dde8a35d1654b9520c92e7['h0152a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a96] =  Ifcca41d795dde8a35d1654b9520c92e7['h0152c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a97] =  Ifcca41d795dde8a35d1654b9520c92e7['h0152e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a98] =  Ifcca41d795dde8a35d1654b9520c92e7['h01530] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a99] =  Ifcca41d795dde8a35d1654b9520c92e7['h01532] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01534] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01536] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01538] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0153a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0153c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00a9f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0153e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01540] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01542] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01544] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01546] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01548] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0154a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0154c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0154e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01550] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aa9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01552] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aaa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01554] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aab] =  Ifcca41d795dde8a35d1654b9520c92e7['h01556] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aac] =  Ifcca41d795dde8a35d1654b9520c92e7['h01558] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0155a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0155c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aaf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0155e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01560] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01562] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01564] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01566] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01568] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0156a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0156c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0156e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01570] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ab9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01572] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aba] =  Ifcca41d795dde8a35d1654b9520c92e7['h01574] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00abb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01576] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00abc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01578] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00abd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0157a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00abe] =  Ifcca41d795dde8a35d1654b9520c92e7['h0157c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00abf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0157e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01580] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01582] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01584] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01586] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01588] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0158a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0158c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0158e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01590] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ac9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01592] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aca] =  Ifcca41d795dde8a35d1654b9520c92e7['h01594] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00acb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01596] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00acc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01598] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00acd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0159a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ace] =  Ifcca41d795dde8a35d1654b9520c92e7['h0159c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00acf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0159e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad0] =  Ifcca41d795dde8a35d1654b9520c92e7['h015a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad1] =  Ifcca41d795dde8a35d1654b9520c92e7['h015a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad2] =  Ifcca41d795dde8a35d1654b9520c92e7['h015a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad3] =  Ifcca41d795dde8a35d1654b9520c92e7['h015a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad4] =  Ifcca41d795dde8a35d1654b9520c92e7['h015a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad5] =  Ifcca41d795dde8a35d1654b9520c92e7['h015aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad6] =  Ifcca41d795dde8a35d1654b9520c92e7['h015ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad7] =  Ifcca41d795dde8a35d1654b9520c92e7['h015ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad8] =  Ifcca41d795dde8a35d1654b9520c92e7['h015b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ad9] =  Ifcca41d795dde8a35d1654b9520c92e7['h015b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ada] =  Ifcca41d795dde8a35d1654b9520c92e7['h015b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00adb] =  Ifcca41d795dde8a35d1654b9520c92e7['h015b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00adc] =  Ifcca41d795dde8a35d1654b9520c92e7['h015b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00add] =  Ifcca41d795dde8a35d1654b9520c92e7['h015ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ade] =  Ifcca41d795dde8a35d1654b9520c92e7['h015bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00adf] =  Ifcca41d795dde8a35d1654b9520c92e7['h015be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae0] =  Ifcca41d795dde8a35d1654b9520c92e7['h015c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae1] =  Ifcca41d795dde8a35d1654b9520c92e7['h015c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae2] =  Ifcca41d795dde8a35d1654b9520c92e7['h015c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae3] =  Ifcca41d795dde8a35d1654b9520c92e7['h015c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae4] =  Ifcca41d795dde8a35d1654b9520c92e7['h015c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae5] =  Ifcca41d795dde8a35d1654b9520c92e7['h015ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae6] =  Ifcca41d795dde8a35d1654b9520c92e7['h015cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae7] =  Ifcca41d795dde8a35d1654b9520c92e7['h015ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae8] =  Ifcca41d795dde8a35d1654b9520c92e7['h015d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ae9] =  Ifcca41d795dde8a35d1654b9520c92e7['h015d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aea] =  Ifcca41d795dde8a35d1654b9520c92e7['h015d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aeb] =  Ifcca41d795dde8a35d1654b9520c92e7['h015d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aec] =  Ifcca41d795dde8a35d1654b9520c92e7['h015d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aed] =  Ifcca41d795dde8a35d1654b9520c92e7['h015da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aee] =  Ifcca41d795dde8a35d1654b9520c92e7['h015dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aef] =  Ifcca41d795dde8a35d1654b9520c92e7['h015de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af0] =  Ifcca41d795dde8a35d1654b9520c92e7['h015e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af1] =  Ifcca41d795dde8a35d1654b9520c92e7['h015e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af2] =  Ifcca41d795dde8a35d1654b9520c92e7['h015e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af3] =  Ifcca41d795dde8a35d1654b9520c92e7['h015e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af4] =  Ifcca41d795dde8a35d1654b9520c92e7['h015e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af5] =  Ifcca41d795dde8a35d1654b9520c92e7['h015ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af6] =  Ifcca41d795dde8a35d1654b9520c92e7['h015ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af7] =  Ifcca41d795dde8a35d1654b9520c92e7['h015ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af8] =  Ifcca41d795dde8a35d1654b9520c92e7['h015f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00af9] =  Ifcca41d795dde8a35d1654b9520c92e7['h015f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00afa] =  Ifcca41d795dde8a35d1654b9520c92e7['h015f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00afb] =  Ifcca41d795dde8a35d1654b9520c92e7['h015f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00afc] =  Ifcca41d795dde8a35d1654b9520c92e7['h015f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00afd] =  Ifcca41d795dde8a35d1654b9520c92e7['h015fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00afe] =  Ifcca41d795dde8a35d1654b9520c92e7['h015fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00aff] =  Ifcca41d795dde8a35d1654b9520c92e7['h015fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b00] =  Ifcca41d795dde8a35d1654b9520c92e7['h01600] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b01] =  Ifcca41d795dde8a35d1654b9520c92e7['h01602] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b02] =  Ifcca41d795dde8a35d1654b9520c92e7['h01604] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b03] =  Ifcca41d795dde8a35d1654b9520c92e7['h01606] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b04] =  Ifcca41d795dde8a35d1654b9520c92e7['h01608] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b05] =  Ifcca41d795dde8a35d1654b9520c92e7['h0160a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b06] =  Ifcca41d795dde8a35d1654b9520c92e7['h0160c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b07] =  Ifcca41d795dde8a35d1654b9520c92e7['h0160e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b08] =  Ifcca41d795dde8a35d1654b9520c92e7['h01610] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b09] =  Ifcca41d795dde8a35d1654b9520c92e7['h01612] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01614] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01616] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01618] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0161a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0161c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b0f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0161e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b10] =  Ifcca41d795dde8a35d1654b9520c92e7['h01620] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b11] =  Ifcca41d795dde8a35d1654b9520c92e7['h01622] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b12] =  Ifcca41d795dde8a35d1654b9520c92e7['h01624] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b13] =  Ifcca41d795dde8a35d1654b9520c92e7['h01626] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b14] =  Ifcca41d795dde8a35d1654b9520c92e7['h01628] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b15] =  Ifcca41d795dde8a35d1654b9520c92e7['h0162a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b16] =  Ifcca41d795dde8a35d1654b9520c92e7['h0162c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b17] =  Ifcca41d795dde8a35d1654b9520c92e7['h0162e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b18] =  Ifcca41d795dde8a35d1654b9520c92e7['h01630] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b19] =  Ifcca41d795dde8a35d1654b9520c92e7['h01632] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01634] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01636] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01638] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0163a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0163c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b1f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0163e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b20] =  Ifcca41d795dde8a35d1654b9520c92e7['h01640] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b21] =  Ifcca41d795dde8a35d1654b9520c92e7['h01642] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b22] =  Ifcca41d795dde8a35d1654b9520c92e7['h01644] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b23] =  Ifcca41d795dde8a35d1654b9520c92e7['h01646] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b24] =  Ifcca41d795dde8a35d1654b9520c92e7['h01648] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b25] =  Ifcca41d795dde8a35d1654b9520c92e7['h0164a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b26] =  Ifcca41d795dde8a35d1654b9520c92e7['h0164c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b27] =  Ifcca41d795dde8a35d1654b9520c92e7['h0164e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b28] =  Ifcca41d795dde8a35d1654b9520c92e7['h01650] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b29] =  Ifcca41d795dde8a35d1654b9520c92e7['h01652] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01654] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01656] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01658] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0165a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0165c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b2f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0165e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b30] =  Ifcca41d795dde8a35d1654b9520c92e7['h01660] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b31] =  Ifcca41d795dde8a35d1654b9520c92e7['h01662] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b32] =  Ifcca41d795dde8a35d1654b9520c92e7['h01664] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b33] =  Ifcca41d795dde8a35d1654b9520c92e7['h01666] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b34] =  Ifcca41d795dde8a35d1654b9520c92e7['h01668] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b35] =  Ifcca41d795dde8a35d1654b9520c92e7['h0166a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b36] =  Ifcca41d795dde8a35d1654b9520c92e7['h0166c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b37] =  Ifcca41d795dde8a35d1654b9520c92e7['h0166e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b38] =  Ifcca41d795dde8a35d1654b9520c92e7['h01670] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b39] =  Ifcca41d795dde8a35d1654b9520c92e7['h01672] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01674] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01676] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01678] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0167a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0167c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b3f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0167e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b40] =  Ifcca41d795dde8a35d1654b9520c92e7['h01680] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b41] =  Ifcca41d795dde8a35d1654b9520c92e7['h01682] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b42] =  Ifcca41d795dde8a35d1654b9520c92e7['h01684] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b43] =  Ifcca41d795dde8a35d1654b9520c92e7['h01686] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b44] =  Ifcca41d795dde8a35d1654b9520c92e7['h01688] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b45] =  Ifcca41d795dde8a35d1654b9520c92e7['h0168a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b46] =  Ifcca41d795dde8a35d1654b9520c92e7['h0168c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b47] =  Ifcca41d795dde8a35d1654b9520c92e7['h0168e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b48] =  Ifcca41d795dde8a35d1654b9520c92e7['h01690] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b49] =  Ifcca41d795dde8a35d1654b9520c92e7['h01692] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01694] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01696] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01698] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0169a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0169c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b4f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0169e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b50] =  Ifcca41d795dde8a35d1654b9520c92e7['h016a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b51] =  Ifcca41d795dde8a35d1654b9520c92e7['h016a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b52] =  Ifcca41d795dde8a35d1654b9520c92e7['h016a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b53] =  Ifcca41d795dde8a35d1654b9520c92e7['h016a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b54] =  Ifcca41d795dde8a35d1654b9520c92e7['h016a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b55] =  Ifcca41d795dde8a35d1654b9520c92e7['h016aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b56] =  Ifcca41d795dde8a35d1654b9520c92e7['h016ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b57] =  Ifcca41d795dde8a35d1654b9520c92e7['h016ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b58] =  Ifcca41d795dde8a35d1654b9520c92e7['h016b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b59] =  Ifcca41d795dde8a35d1654b9520c92e7['h016b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5a] =  Ifcca41d795dde8a35d1654b9520c92e7['h016b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5b] =  Ifcca41d795dde8a35d1654b9520c92e7['h016b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5c] =  Ifcca41d795dde8a35d1654b9520c92e7['h016b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5d] =  Ifcca41d795dde8a35d1654b9520c92e7['h016ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5e] =  Ifcca41d795dde8a35d1654b9520c92e7['h016bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b5f] =  Ifcca41d795dde8a35d1654b9520c92e7['h016be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b60] =  Ifcca41d795dde8a35d1654b9520c92e7['h016c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b61] =  Ifcca41d795dde8a35d1654b9520c92e7['h016c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b62] =  Ifcca41d795dde8a35d1654b9520c92e7['h016c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b63] =  Ifcca41d795dde8a35d1654b9520c92e7['h016c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b64] =  Ifcca41d795dde8a35d1654b9520c92e7['h016c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b65] =  Ifcca41d795dde8a35d1654b9520c92e7['h016ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b66] =  Ifcca41d795dde8a35d1654b9520c92e7['h016cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b67] =  Ifcca41d795dde8a35d1654b9520c92e7['h016ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b68] =  Ifcca41d795dde8a35d1654b9520c92e7['h016d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b69] =  Ifcca41d795dde8a35d1654b9520c92e7['h016d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6a] =  Ifcca41d795dde8a35d1654b9520c92e7['h016d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6b] =  Ifcca41d795dde8a35d1654b9520c92e7['h016d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6c] =  Ifcca41d795dde8a35d1654b9520c92e7['h016d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6d] =  Ifcca41d795dde8a35d1654b9520c92e7['h016da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6e] =  Ifcca41d795dde8a35d1654b9520c92e7['h016dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b6f] =  Ifcca41d795dde8a35d1654b9520c92e7['h016de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b70] =  Ifcca41d795dde8a35d1654b9520c92e7['h016e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b71] =  Ifcca41d795dde8a35d1654b9520c92e7['h016e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b72] =  Ifcca41d795dde8a35d1654b9520c92e7['h016e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b73] =  Ifcca41d795dde8a35d1654b9520c92e7['h016e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b74] =  Ifcca41d795dde8a35d1654b9520c92e7['h016e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b75] =  Ifcca41d795dde8a35d1654b9520c92e7['h016ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b76] =  Ifcca41d795dde8a35d1654b9520c92e7['h016ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b77] =  Ifcca41d795dde8a35d1654b9520c92e7['h016ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b78] =  Ifcca41d795dde8a35d1654b9520c92e7['h016f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b79] =  Ifcca41d795dde8a35d1654b9520c92e7['h016f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7a] =  Ifcca41d795dde8a35d1654b9520c92e7['h016f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7b] =  Ifcca41d795dde8a35d1654b9520c92e7['h016f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7c] =  Ifcca41d795dde8a35d1654b9520c92e7['h016f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7d] =  Ifcca41d795dde8a35d1654b9520c92e7['h016fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7e] =  Ifcca41d795dde8a35d1654b9520c92e7['h016fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b7f] =  Ifcca41d795dde8a35d1654b9520c92e7['h016fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b80] =  Ifcca41d795dde8a35d1654b9520c92e7['h01700] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b81] =  Ifcca41d795dde8a35d1654b9520c92e7['h01702] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b82] =  Ifcca41d795dde8a35d1654b9520c92e7['h01704] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b83] =  Ifcca41d795dde8a35d1654b9520c92e7['h01706] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b84] =  Ifcca41d795dde8a35d1654b9520c92e7['h01708] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b85] =  Ifcca41d795dde8a35d1654b9520c92e7['h0170a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b86] =  Ifcca41d795dde8a35d1654b9520c92e7['h0170c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b87] =  Ifcca41d795dde8a35d1654b9520c92e7['h0170e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b88] =  Ifcca41d795dde8a35d1654b9520c92e7['h01710] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b89] =  Ifcca41d795dde8a35d1654b9520c92e7['h01712] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01714] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01716] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01718] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0171a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0171c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b8f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0171e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b90] =  Ifcca41d795dde8a35d1654b9520c92e7['h01720] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b91] =  Ifcca41d795dde8a35d1654b9520c92e7['h01722] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b92] =  Ifcca41d795dde8a35d1654b9520c92e7['h01724] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b93] =  Ifcca41d795dde8a35d1654b9520c92e7['h01726] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b94] =  Ifcca41d795dde8a35d1654b9520c92e7['h01728] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b95] =  Ifcca41d795dde8a35d1654b9520c92e7['h0172a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b96] =  Ifcca41d795dde8a35d1654b9520c92e7['h0172c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b97] =  Ifcca41d795dde8a35d1654b9520c92e7['h0172e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b98] =  Ifcca41d795dde8a35d1654b9520c92e7['h01730] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b99] =  Ifcca41d795dde8a35d1654b9520c92e7['h01732] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01734] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01736] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01738] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0173a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0173c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00b9f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0173e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01740] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01742] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01744] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01746] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01748] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0174a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0174c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0174e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01750] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ba9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01752] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00baa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01754] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bab] =  Ifcca41d795dde8a35d1654b9520c92e7['h01756] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bac] =  Ifcca41d795dde8a35d1654b9520c92e7['h01758] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0175a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0175c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00baf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0175e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01760] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01762] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01764] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01766] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01768] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0176a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0176c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0176e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01770] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bb9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01772] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bba] =  Ifcca41d795dde8a35d1654b9520c92e7['h01774] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bbb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01776] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bbc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01778] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bbd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0177a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bbe] =  Ifcca41d795dde8a35d1654b9520c92e7['h0177c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bbf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0177e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01780] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01782] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01784] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01786] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01788] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0178a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0178c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0178e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01790] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bc9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01792] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bca] =  Ifcca41d795dde8a35d1654b9520c92e7['h01794] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bcb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01796] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bcc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01798] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bcd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0179a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0179c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bcf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0179e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd0] =  Ifcca41d795dde8a35d1654b9520c92e7['h017a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd1] =  Ifcca41d795dde8a35d1654b9520c92e7['h017a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd2] =  Ifcca41d795dde8a35d1654b9520c92e7['h017a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd3] =  Ifcca41d795dde8a35d1654b9520c92e7['h017a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd4] =  Ifcca41d795dde8a35d1654b9520c92e7['h017a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd5] =  Ifcca41d795dde8a35d1654b9520c92e7['h017aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd6] =  Ifcca41d795dde8a35d1654b9520c92e7['h017ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd7] =  Ifcca41d795dde8a35d1654b9520c92e7['h017ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd8] =  Ifcca41d795dde8a35d1654b9520c92e7['h017b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bd9] =  Ifcca41d795dde8a35d1654b9520c92e7['h017b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bda] =  Ifcca41d795dde8a35d1654b9520c92e7['h017b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bdb] =  Ifcca41d795dde8a35d1654b9520c92e7['h017b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bdc] =  Ifcca41d795dde8a35d1654b9520c92e7['h017b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bdd] =  Ifcca41d795dde8a35d1654b9520c92e7['h017ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bde] =  Ifcca41d795dde8a35d1654b9520c92e7['h017bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bdf] =  Ifcca41d795dde8a35d1654b9520c92e7['h017be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be0] =  Ifcca41d795dde8a35d1654b9520c92e7['h017c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be1] =  Ifcca41d795dde8a35d1654b9520c92e7['h017c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be2] =  Ifcca41d795dde8a35d1654b9520c92e7['h017c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be3] =  Ifcca41d795dde8a35d1654b9520c92e7['h017c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be4] =  Ifcca41d795dde8a35d1654b9520c92e7['h017c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be5] =  Ifcca41d795dde8a35d1654b9520c92e7['h017ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be6] =  Ifcca41d795dde8a35d1654b9520c92e7['h017cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be7] =  Ifcca41d795dde8a35d1654b9520c92e7['h017ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be8] =  Ifcca41d795dde8a35d1654b9520c92e7['h017d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00be9] =  Ifcca41d795dde8a35d1654b9520c92e7['h017d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bea] =  Ifcca41d795dde8a35d1654b9520c92e7['h017d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00beb] =  Ifcca41d795dde8a35d1654b9520c92e7['h017d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bec] =  Ifcca41d795dde8a35d1654b9520c92e7['h017d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bed] =  Ifcca41d795dde8a35d1654b9520c92e7['h017da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bee] =  Ifcca41d795dde8a35d1654b9520c92e7['h017dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bef] =  Ifcca41d795dde8a35d1654b9520c92e7['h017de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf0] =  Ifcca41d795dde8a35d1654b9520c92e7['h017e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf1] =  Ifcca41d795dde8a35d1654b9520c92e7['h017e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf2] =  Ifcca41d795dde8a35d1654b9520c92e7['h017e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf3] =  Ifcca41d795dde8a35d1654b9520c92e7['h017e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf4] =  Ifcca41d795dde8a35d1654b9520c92e7['h017e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf5] =  Ifcca41d795dde8a35d1654b9520c92e7['h017ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf6] =  Ifcca41d795dde8a35d1654b9520c92e7['h017ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf7] =  Ifcca41d795dde8a35d1654b9520c92e7['h017ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf8] =  Ifcca41d795dde8a35d1654b9520c92e7['h017f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bf9] =  Ifcca41d795dde8a35d1654b9520c92e7['h017f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bfa] =  Ifcca41d795dde8a35d1654b9520c92e7['h017f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bfb] =  Ifcca41d795dde8a35d1654b9520c92e7['h017f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bfc] =  Ifcca41d795dde8a35d1654b9520c92e7['h017f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bfd] =  Ifcca41d795dde8a35d1654b9520c92e7['h017fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bfe] =  Ifcca41d795dde8a35d1654b9520c92e7['h017fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00bff] =  Ifcca41d795dde8a35d1654b9520c92e7['h017fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c00] =  Ifcca41d795dde8a35d1654b9520c92e7['h01800] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c01] =  Ifcca41d795dde8a35d1654b9520c92e7['h01802] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c02] =  Ifcca41d795dde8a35d1654b9520c92e7['h01804] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c03] =  Ifcca41d795dde8a35d1654b9520c92e7['h01806] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c04] =  Ifcca41d795dde8a35d1654b9520c92e7['h01808] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c05] =  Ifcca41d795dde8a35d1654b9520c92e7['h0180a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c06] =  Ifcca41d795dde8a35d1654b9520c92e7['h0180c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c07] =  Ifcca41d795dde8a35d1654b9520c92e7['h0180e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c08] =  Ifcca41d795dde8a35d1654b9520c92e7['h01810] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c09] =  Ifcca41d795dde8a35d1654b9520c92e7['h01812] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01814] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01816] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01818] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0181a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0181c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c0f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0181e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c10] =  Ifcca41d795dde8a35d1654b9520c92e7['h01820] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c11] =  Ifcca41d795dde8a35d1654b9520c92e7['h01822] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c12] =  Ifcca41d795dde8a35d1654b9520c92e7['h01824] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c13] =  Ifcca41d795dde8a35d1654b9520c92e7['h01826] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c14] =  Ifcca41d795dde8a35d1654b9520c92e7['h01828] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c15] =  Ifcca41d795dde8a35d1654b9520c92e7['h0182a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c16] =  Ifcca41d795dde8a35d1654b9520c92e7['h0182c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c17] =  Ifcca41d795dde8a35d1654b9520c92e7['h0182e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c18] =  Ifcca41d795dde8a35d1654b9520c92e7['h01830] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c19] =  Ifcca41d795dde8a35d1654b9520c92e7['h01832] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01834] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01836] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01838] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0183a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0183c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c1f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0183e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c20] =  Ifcca41d795dde8a35d1654b9520c92e7['h01840] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c21] =  Ifcca41d795dde8a35d1654b9520c92e7['h01842] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c22] =  Ifcca41d795dde8a35d1654b9520c92e7['h01844] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c23] =  Ifcca41d795dde8a35d1654b9520c92e7['h01846] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c24] =  Ifcca41d795dde8a35d1654b9520c92e7['h01848] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c25] =  Ifcca41d795dde8a35d1654b9520c92e7['h0184a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c26] =  Ifcca41d795dde8a35d1654b9520c92e7['h0184c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c27] =  Ifcca41d795dde8a35d1654b9520c92e7['h0184e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c28] =  Ifcca41d795dde8a35d1654b9520c92e7['h01850] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c29] =  Ifcca41d795dde8a35d1654b9520c92e7['h01852] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01854] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01856] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01858] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0185a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0185c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c2f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0185e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c30] =  Ifcca41d795dde8a35d1654b9520c92e7['h01860] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c31] =  Ifcca41d795dde8a35d1654b9520c92e7['h01862] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c32] =  Ifcca41d795dde8a35d1654b9520c92e7['h01864] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c33] =  Ifcca41d795dde8a35d1654b9520c92e7['h01866] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c34] =  Ifcca41d795dde8a35d1654b9520c92e7['h01868] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c35] =  Ifcca41d795dde8a35d1654b9520c92e7['h0186a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c36] =  Ifcca41d795dde8a35d1654b9520c92e7['h0186c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c37] =  Ifcca41d795dde8a35d1654b9520c92e7['h0186e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c38] =  Ifcca41d795dde8a35d1654b9520c92e7['h01870] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c39] =  Ifcca41d795dde8a35d1654b9520c92e7['h01872] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01874] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01876] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01878] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0187a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0187c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c3f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0187e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c40] =  Ifcca41d795dde8a35d1654b9520c92e7['h01880] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c41] =  Ifcca41d795dde8a35d1654b9520c92e7['h01882] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c42] =  Ifcca41d795dde8a35d1654b9520c92e7['h01884] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c43] =  Ifcca41d795dde8a35d1654b9520c92e7['h01886] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c44] =  Ifcca41d795dde8a35d1654b9520c92e7['h01888] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c45] =  Ifcca41d795dde8a35d1654b9520c92e7['h0188a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c46] =  Ifcca41d795dde8a35d1654b9520c92e7['h0188c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c47] =  Ifcca41d795dde8a35d1654b9520c92e7['h0188e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c48] =  Ifcca41d795dde8a35d1654b9520c92e7['h01890] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c49] =  Ifcca41d795dde8a35d1654b9520c92e7['h01892] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01894] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01896] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01898] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0189a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0189c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c4f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0189e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c50] =  Ifcca41d795dde8a35d1654b9520c92e7['h018a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c51] =  Ifcca41d795dde8a35d1654b9520c92e7['h018a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c52] =  Ifcca41d795dde8a35d1654b9520c92e7['h018a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c53] =  Ifcca41d795dde8a35d1654b9520c92e7['h018a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c54] =  Ifcca41d795dde8a35d1654b9520c92e7['h018a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c55] =  Ifcca41d795dde8a35d1654b9520c92e7['h018aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c56] =  Ifcca41d795dde8a35d1654b9520c92e7['h018ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c57] =  Ifcca41d795dde8a35d1654b9520c92e7['h018ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c58] =  Ifcca41d795dde8a35d1654b9520c92e7['h018b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c59] =  Ifcca41d795dde8a35d1654b9520c92e7['h018b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5a] =  Ifcca41d795dde8a35d1654b9520c92e7['h018b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5b] =  Ifcca41d795dde8a35d1654b9520c92e7['h018b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5c] =  Ifcca41d795dde8a35d1654b9520c92e7['h018b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5d] =  Ifcca41d795dde8a35d1654b9520c92e7['h018ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5e] =  Ifcca41d795dde8a35d1654b9520c92e7['h018bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c5f] =  Ifcca41d795dde8a35d1654b9520c92e7['h018be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c60] =  Ifcca41d795dde8a35d1654b9520c92e7['h018c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c61] =  Ifcca41d795dde8a35d1654b9520c92e7['h018c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c62] =  Ifcca41d795dde8a35d1654b9520c92e7['h018c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c63] =  Ifcca41d795dde8a35d1654b9520c92e7['h018c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c64] =  Ifcca41d795dde8a35d1654b9520c92e7['h018c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c65] =  Ifcca41d795dde8a35d1654b9520c92e7['h018ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c66] =  Ifcca41d795dde8a35d1654b9520c92e7['h018cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c67] =  Ifcca41d795dde8a35d1654b9520c92e7['h018ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c68] =  Ifcca41d795dde8a35d1654b9520c92e7['h018d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c69] =  Ifcca41d795dde8a35d1654b9520c92e7['h018d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6a] =  Ifcca41d795dde8a35d1654b9520c92e7['h018d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6b] =  Ifcca41d795dde8a35d1654b9520c92e7['h018d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6c] =  Ifcca41d795dde8a35d1654b9520c92e7['h018d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6d] =  Ifcca41d795dde8a35d1654b9520c92e7['h018da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6e] =  Ifcca41d795dde8a35d1654b9520c92e7['h018dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c6f] =  Ifcca41d795dde8a35d1654b9520c92e7['h018de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c70] =  Ifcca41d795dde8a35d1654b9520c92e7['h018e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c71] =  Ifcca41d795dde8a35d1654b9520c92e7['h018e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c72] =  Ifcca41d795dde8a35d1654b9520c92e7['h018e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c73] =  Ifcca41d795dde8a35d1654b9520c92e7['h018e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c74] =  Ifcca41d795dde8a35d1654b9520c92e7['h018e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c75] =  Ifcca41d795dde8a35d1654b9520c92e7['h018ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c76] =  Ifcca41d795dde8a35d1654b9520c92e7['h018ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c77] =  Ifcca41d795dde8a35d1654b9520c92e7['h018ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c78] =  Ifcca41d795dde8a35d1654b9520c92e7['h018f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c79] =  Ifcca41d795dde8a35d1654b9520c92e7['h018f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7a] =  Ifcca41d795dde8a35d1654b9520c92e7['h018f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7b] =  Ifcca41d795dde8a35d1654b9520c92e7['h018f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7c] =  Ifcca41d795dde8a35d1654b9520c92e7['h018f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7d] =  Ifcca41d795dde8a35d1654b9520c92e7['h018fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7e] =  Ifcca41d795dde8a35d1654b9520c92e7['h018fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c7f] =  Ifcca41d795dde8a35d1654b9520c92e7['h018fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c80] =  Ifcca41d795dde8a35d1654b9520c92e7['h01900] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c81] =  Ifcca41d795dde8a35d1654b9520c92e7['h01902] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c82] =  Ifcca41d795dde8a35d1654b9520c92e7['h01904] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c83] =  Ifcca41d795dde8a35d1654b9520c92e7['h01906] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c84] =  Ifcca41d795dde8a35d1654b9520c92e7['h01908] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c85] =  Ifcca41d795dde8a35d1654b9520c92e7['h0190a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c86] =  Ifcca41d795dde8a35d1654b9520c92e7['h0190c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c87] =  Ifcca41d795dde8a35d1654b9520c92e7['h0190e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c88] =  Ifcca41d795dde8a35d1654b9520c92e7['h01910] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c89] =  Ifcca41d795dde8a35d1654b9520c92e7['h01912] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01914] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01916] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01918] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0191a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0191c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c8f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0191e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c90] =  Ifcca41d795dde8a35d1654b9520c92e7['h01920] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c91] =  Ifcca41d795dde8a35d1654b9520c92e7['h01922] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c92] =  Ifcca41d795dde8a35d1654b9520c92e7['h01924] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c93] =  Ifcca41d795dde8a35d1654b9520c92e7['h01926] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c94] =  Ifcca41d795dde8a35d1654b9520c92e7['h01928] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c95] =  Ifcca41d795dde8a35d1654b9520c92e7['h0192a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c96] =  Ifcca41d795dde8a35d1654b9520c92e7['h0192c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c97] =  Ifcca41d795dde8a35d1654b9520c92e7['h0192e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c98] =  Ifcca41d795dde8a35d1654b9520c92e7['h01930] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c99] =  Ifcca41d795dde8a35d1654b9520c92e7['h01932] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01934] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01936] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01938] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9d] =  Ifcca41d795dde8a35d1654b9520c92e7['h0193a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9e] =  Ifcca41d795dde8a35d1654b9520c92e7['h0193c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00c9f] =  Ifcca41d795dde8a35d1654b9520c92e7['h0193e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01940] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01942] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01944] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01946] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01948] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0194a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0194c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0194e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01950] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ca9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01952] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00caa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01954] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cab] =  Ifcca41d795dde8a35d1654b9520c92e7['h01956] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cac] =  Ifcca41d795dde8a35d1654b9520c92e7['h01958] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cad] =  Ifcca41d795dde8a35d1654b9520c92e7['h0195a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cae] =  Ifcca41d795dde8a35d1654b9520c92e7['h0195c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00caf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0195e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01960] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01962] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01964] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01966] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01968] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0196a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0196c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0196e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01970] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cb9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01972] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cba] =  Ifcca41d795dde8a35d1654b9520c92e7['h01974] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cbb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01976] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cbc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01978] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cbd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0197a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cbe] =  Ifcca41d795dde8a35d1654b9520c92e7['h0197c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cbf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0197e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01980] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01982] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01984] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01986] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01988] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc5] =  Ifcca41d795dde8a35d1654b9520c92e7['h0198a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc6] =  Ifcca41d795dde8a35d1654b9520c92e7['h0198c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc7] =  Ifcca41d795dde8a35d1654b9520c92e7['h0198e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01990] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cc9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01992] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cca] =  Ifcca41d795dde8a35d1654b9520c92e7['h01994] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ccb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01996] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ccc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01998] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ccd] =  Ifcca41d795dde8a35d1654b9520c92e7['h0199a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cce] =  Ifcca41d795dde8a35d1654b9520c92e7['h0199c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ccf] =  Ifcca41d795dde8a35d1654b9520c92e7['h0199e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd0] =  Ifcca41d795dde8a35d1654b9520c92e7['h019a0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd1] =  Ifcca41d795dde8a35d1654b9520c92e7['h019a2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd2] =  Ifcca41d795dde8a35d1654b9520c92e7['h019a4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd3] =  Ifcca41d795dde8a35d1654b9520c92e7['h019a6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd4] =  Ifcca41d795dde8a35d1654b9520c92e7['h019a8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd5] =  Ifcca41d795dde8a35d1654b9520c92e7['h019aa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd6] =  Ifcca41d795dde8a35d1654b9520c92e7['h019ac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd7] =  Ifcca41d795dde8a35d1654b9520c92e7['h019ae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd8] =  Ifcca41d795dde8a35d1654b9520c92e7['h019b0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cd9] =  Ifcca41d795dde8a35d1654b9520c92e7['h019b2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cda] =  Ifcca41d795dde8a35d1654b9520c92e7['h019b4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cdb] =  Ifcca41d795dde8a35d1654b9520c92e7['h019b6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cdc] =  Ifcca41d795dde8a35d1654b9520c92e7['h019b8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cdd] =  Ifcca41d795dde8a35d1654b9520c92e7['h019ba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cde] =  Ifcca41d795dde8a35d1654b9520c92e7['h019bc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cdf] =  Ifcca41d795dde8a35d1654b9520c92e7['h019be] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce0] =  Ifcca41d795dde8a35d1654b9520c92e7['h019c0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce1] =  Ifcca41d795dde8a35d1654b9520c92e7['h019c2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce2] =  Ifcca41d795dde8a35d1654b9520c92e7['h019c4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce3] =  Ifcca41d795dde8a35d1654b9520c92e7['h019c6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce4] =  Ifcca41d795dde8a35d1654b9520c92e7['h019c8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce5] =  Ifcca41d795dde8a35d1654b9520c92e7['h019ca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce6] =  Ifcca41d795dde8a35d1654b9520c92e7['h019cc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce7] =  Ifcca41d795dde8a35d1654b9520c92e7['h019ce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce8] =  Ifcca41d795dde8a35d1654b9520c92e7['h019d0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ce9] =  Ifcca41d795dde8a35d1654b9520c92e7['h019d2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cea] =  Ifcca41d795dde8a35d1654b9520c92e7['h019d4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ceb] =  Ifcca41d795dde8a35d1654b9520c92e7['h019d6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cec] =  Ifcca41d795dde8a35d1654b9520c92e7['h019d8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ced] =  Ifcca41d795dde8a35d1654b9520c92e7['h019da] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cee] =  Ifcca41d795dde8a35d1654b9520c92e7['h019dc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cef] =  Ifcca41d795dde8a35d1654b9520c92e7['h019de] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf0] =  Ifcca41d795dde8a35d1654b9520c92e7['h019e0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf1] =  Ifcca41d795dde8a35d1654b9520c92e7['h019e2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf2] =  Ifcca41d795dde8a35d1654b9520c92e7['h019e4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf3] =  Ifcca41d795dde8a35d1654b9520c92e7['h019e6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf4] =  Ifcca41d795dde8a35d1654b9520c92e7['h019e8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf5] =  Ifcca41d795dde8a35d1654b9520c92e7['h019ea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf6] =  Ifcca41d795dde8a35d1654b9520c92e7['h019ec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf7] =  Ifcca41d795dde8a35d1654b9520c92e7['h019ee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf8] =  Ifcca41d795dde8a35d1654b9520c92e7['h019f0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cf9] =  Ifcca41d795dde8a35d1654b9520c92e7['h019f2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cfa] =  Ifcca41d795dde8a35d1654b9520c92e7['h019f4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cfb] =  Ifcca41d795dde8a35d1654b9520c92e7['h019f6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cfc] =  Ifcca41d795dde8a35d1654b9520c92e7['h019f8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cfd] =  Ifcca41d795dde8a35d1654b9520c92e7['h019fa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cfe] =  Ifcca41d795dde8a35d1654b9520c92e7['h019fc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00cff] =  Ifcca41d795dde8a35d1654b9520c92e7['h019fe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d00] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d01] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d02] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d03] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d04] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d05] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d06] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d07] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d08] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d09] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d0f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d10] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d11] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d12] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d13] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d14] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d15] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d16] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d17] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d18] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d19] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d1f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d20] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d21] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d22] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d23] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d24] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d25] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d26] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d27] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d28] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d29] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d2f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d30] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d31] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d32] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d33] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d34] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d35] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d36] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d37] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d38] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d39] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d3f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d40] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d41] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d42] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d43] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d44] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d45] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d46] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d47] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d48] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d49] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d4f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01a9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d50] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aa0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d51] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aa2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d52] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aa4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d53] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aa6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d54] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aa8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d55] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aaa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d56] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d57] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d58] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ab0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d59] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ab2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ab4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ab6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ab8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01abc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d5f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01abe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d60] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ac0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d61] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ac2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d62] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ac4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d63] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ac6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d64] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ac8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d65] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d66] =  Ifcca41d795dde8a35d1654b9520c92e7['h01acc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d67] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ace] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d68] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ad0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d69] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ad2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ad4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ad6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ad8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ada] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01adc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d6f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ade] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d70] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ae0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d71] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ae2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d72] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ae4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d73] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ae6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d74] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ae8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d75] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d76] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d77] =  Ifcca41d795dde8a35d1654b9520c92e7['h01aee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d78] =  Ifcca41d795dde8a35d1654b9520c92e7['h01af0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d79] =  Ifcca41d795dde8a35d1654b9520c92e7['h01af2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01af4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01af6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01af8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01afa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01afc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d7f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01afe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d80] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d81] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d82] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d83] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d84] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d85] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d86] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d87] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d88] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d89] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d8f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d90] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d91] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d92] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d93] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d94] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d95] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d96] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d97] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d98] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d99] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00d9f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00da9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00daa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dab] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dac] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dad] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dae] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00daf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00db9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dba] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dbb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dbc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dbd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dbe] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dbf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dc9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dca] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dcb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dcc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dcd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dce] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dcf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01b9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ba0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ba2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ba4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ba6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ba8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01baa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bb0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dd9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bb2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dda] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bb4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ddb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bb6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ddc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bb8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ddd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dde] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bbc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ddf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bbe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bc0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bc2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bc4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bc6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bc8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bcc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bd0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00de9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bd2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dea] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bd4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00deb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bd6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dec] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bd8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ded] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dee] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bdc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00def] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bde] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01be0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01be2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01be4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01be6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01be8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bf0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00df9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bf2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dfa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bf4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dfb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bf6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dfc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bf8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dfd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bfa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dfe] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bfc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00dff] =  Ifcca41d795dde8a35d1654b9520c92e7['h01bfe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e00] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e01] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e02] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e03] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e04] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e05] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e06] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e07] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e08] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e09] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e0f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e10] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e11] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e12] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e13] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e14] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e15] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e16] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e17] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e18] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e19] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e1f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e20] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e21] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e22] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e23] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e24] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e25] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e26] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e27] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e28] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e29] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e2f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e30] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e31] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e32] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e33] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e34] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e35] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e36] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e37] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e38] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e39] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e3f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e40] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e41] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e42] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e43] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e44] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e45] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e46] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e47] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e48] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e49] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e4f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01c9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e50] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ca0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e51] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ca2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e52] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ca4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e53] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ca6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e54] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ca8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e55] =  Ifcca41d795dde8a35d1654b9520c92e7['h01caa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e56] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e57] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e58] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cb0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e59] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cb2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cb4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cb6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cb8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cbc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e5f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cbe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e60] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cc0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e61] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cc2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e62] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cc4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e63] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cc6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e64] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cc8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e65] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e66] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ccc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e67] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e68] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cd0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e69] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cd2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cd4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cd6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cd8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cdc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e6f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cde] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e70] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ce0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e71] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ce2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e72] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ce4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e73] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ce6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e74] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ce8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e75] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e76] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e77] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e78] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cf0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e79] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cf2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cf4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cf6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cf8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cfa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cfc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e7f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01cfe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e80] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e81] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e82] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e83] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e84] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e85] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e86] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e87] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e88] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e89] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e8f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e90] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e91] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e92] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e93] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e94] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e95] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e96] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e97] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e98] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e99] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00e9f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ea9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eaa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eab] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eac] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ead] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eae] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eaf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eb9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eba] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ebb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ebc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ebd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ebe] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ebf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ec9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eca] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ecb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ecc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ecd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ece] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ecf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01d9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01da0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01da2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01da4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01da6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01da8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01daa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01db0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ed9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01db2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eda] =  Ifcca41d795dde8a35d1654b9520c92e7['h01db4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00edb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01db6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00edc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01db8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00edd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ede] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dbc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00edf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dbe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dc0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dc2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dc4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dc6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dc8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dcc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dd0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ee9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dd2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eea] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dd4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eeb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dd6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eec] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dd8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eed] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eee] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ddc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eef] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dde] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01de0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01de2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01de4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01de6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01de8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01df0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ef9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01df2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00efa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01df4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00efb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01df6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00efc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01df8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00efd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dfa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00efe] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dfc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00eff] =  Ifcca41d795dde8a35d1654b9520c92e7['h01dfe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f00] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f01] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f02] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f03] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f04] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f05] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f06] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f07] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f08] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f09] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f0f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f10] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f11] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f12] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f13] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f14] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f15] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f16] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f17] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f18] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f19] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f1f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f20] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f21] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f22] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f23] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f24] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f25] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f26] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f27] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f28] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f29] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f2f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f30] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f31] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f32] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f33] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f34] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f35] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f36] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f37] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f38] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f39] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f3f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f40] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f41] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f42] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f43] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f44] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f45] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f46] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f47] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f48] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f49] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f4f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01e9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f50] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ea0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f51] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ea2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f52] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ea4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f53] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ea6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f54] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ea8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f55] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eaa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f56] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f57] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f58] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eb0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f59] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eb2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eb4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eb6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eb8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ebc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f5f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ebe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f60] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ec0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f61] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ec2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f62] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ec4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f63] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ec6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f64] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ec8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f65] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f66] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ecc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f67] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ece] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f68] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ed0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f69] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ed2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ed4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ed6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ed8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01edc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f6f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ede] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f70] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ee0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f71] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ee2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f72] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ee4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f73] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ee6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f74] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ee8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f75] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f76] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f77] =  Ifcca41d795dde8a35d1654b9520c92e7['h01eee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f78] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ef0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f79] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ef2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ef4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ef6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ef8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01efa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01efc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f7f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01efe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f80] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f00] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f81] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f02] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f82] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f04] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f83] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f06] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f84] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f08] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f85] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f0a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f86] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f0c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f87] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f0e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f88] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f10] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f89] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f12] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f14] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f16] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f18] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f1a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f1c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f8f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f1e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f90] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f20] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f91] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f22] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f92] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f24] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f93] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f26] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f94] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f28] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f95] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f2a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f96] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f2c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f97] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f2e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f98] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f30] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f99] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f32] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9a] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f34] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9b] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f36] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9c] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f38] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9d] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f3a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9e] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f3c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00f9f] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f3e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f40] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f42] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f44] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f46] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f48] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f4a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f4c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f4e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f50] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fa9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f52] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00faa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f54] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fab] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f56] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fac] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f58] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fad] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f5a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fae] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f5c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00faf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f5e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f60] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f62] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f64] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f66] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f68] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f6a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f6c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f6e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f70] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fb9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f72] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fba] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f74] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fbb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f76] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fbc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f78] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fbd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f7a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fbe] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f7c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fbf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f7e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f80] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f82] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f84] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f86] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f88] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f8a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f8c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f8e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f90] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fc9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f92] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fca] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f94] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fcb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f96] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fcc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f98] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fcd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f9a] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fce] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f9c] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fcf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01f9e] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fa0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fa2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fa4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fa6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fa8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01faa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fac] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fae] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fb0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fd9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fb2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fda] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fb4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fdb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fb6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fdc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fb8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fdd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fba] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fde] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fbc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fdf] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fbe] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fc0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fc2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fc4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fc6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fc8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fca] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fcc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fce] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fd0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fe9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fd2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fea] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fd4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00feb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fd6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fec] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fd8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fed] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fda] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fee] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fdc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fef] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fde] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff0] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fe0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff1] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fe2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff2] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fe4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff3] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fe6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff4] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fe8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff5] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fea] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff6] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fec] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff7] =  Ifcca41d795dde8a35d1654b9520c92e7['h01fee] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff8] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ff0] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ff9] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ff2] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ffa] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ff4] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ffb] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ff6] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ffc] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ff8] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ffd] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ffa] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00ffe] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ffc] ;
//end
//always_comb begin // 
               I1b23c494e0c04cc5a8a3ff99b6cdf26d['h00fff] =  Ifcca41d795dde8a35d1654b9520c92e7['h01ffe] ;
//end
