 reg  ['h7ff:0] [$clog2('h7000+1)-1:0] I38e438ab568822a1c40149a2acc5d876 ;
