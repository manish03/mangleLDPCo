 reg  ['h3f:0] [$clog2('h7000+1)-1:0] Ia2f891646e6ab8d9fb9ea77d93148790 ;
