 reg  ['h0:0] [$clog2('h7000+1)-1:0] I6be0bfc1327465230710d1b067b706d4 ;
