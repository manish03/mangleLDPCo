//#;; Ic23fa9996925b610710d93e28c59a3e2 I10df3d67626099df882920ba6552f16d I93762d802eed04b3e1c59d1d46b35248 Ic9f869114804f0a61ce9b03def9d71f5 I9fc5887c030f7a3e19821ebec457e719
/*I816842ff6f8526885b6ad2d49236bc84*/
////////////////////////////////////////////////////////////////////////////////
//# Copyright (c) 2018 Secantec
//# No Permission to modify and distribute this program
//# even if this copyright message remains unaltered.
//#
//# Author: Secantec 27 April, 2018
//# $Id: $//#
//# Revision History
//#       MM      17  April, 2018    Initial release
//#
////////////////////////////////////////////////////////////////////////////////

// /Ic1111bd512b29e821b120b86446026b8/Id67f249b90615ca158b1258712c3a9fc -Ibea2f3fe6ec7414cdf0bf233abba7ef0 *I66986ae1d2ec0253762b97e22f881595* *If4ed727b4ff4652b44f0b32f7198402e* ; If83a0aa1f9ca0f7dd5994445ba7d9e80 I21f66e7dd81ae29064c26b66d9b3e967.I288404204e3d452229308317344a285d -If83a0aa1f9ca0f7dd5994445ba7d9e80 Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.sv > Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv ; Id6bfe3ce1bf5714887f4ffbb7b94feab -I958fb7ed1fb6d4960d15ffd3254be634 -Ie1e1d3d40573127e9ee0480caf1283d6 -Ia823f97963868b5794f5a36e4dbe5dec Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv -I2db95e8e1a9267b7a1188556b2013b33 Ic4c7fcc09295dba6fc1fd0469d7e92e1.1.I21f66e7dd81ae29064c26b66d9b3e967.sv.Idc1d71bbb5c4d2a5e936db79ef10c19f

 /*I816842ff6f8526885b6ad2d49236bc84*/

/* I0c35fcd8aa6b70a1e6a2f67174222bd1 Ifaf61c215f3a90fcc150ac387f759daf I54a78636e8c6bd0efb73150b779d5eb5 */

module  sntc_ldpc_decoder#(
// NR_2_0_4/I58d53a433022417c56e36facb426c2b8.sv
parameter MM   = 'h 000a8 ,
// parameter MM =  'h  000a8  , 
parameter NN   = 'h 000d0 ,
// parameter NN =  'h  000d0  , 
parameter cmax = 'h 00017 ,
// parameter cmax =  'h  00017  , 
parameter rmax = 'h 0000a ,
// parameter rmax =  'h  0000a  , 






parameter SUM_NN         = $clog2(NN+1), // 8 : I307afb7f348272492f3cca58ef2f95d8
parameter SUM_MM         = $clog2(MM+1), // 8 : If78618843e4df2223e60ec190987c019
parameter LEN            = MM,
parameter SUM_NN_WDTH    = $clog2(SUM_NN+2),
parameter SUM_MM_WDTH    = $clog2(SUM_MM+2),
`include "NR_2_0_4/sntc_LDPC_dec_param.sv"
`include "NR_2_0_4/flogtanh/GF2_LDPC_flogtanh_param_inc.sv"
  ,
`include "NR_2_0_4/fgallag/GF2_LDPC_fgallag_param_inc.sv"
 ,
parameter MAX_SUM_WDTH_L = 24, //MAX_SUM_WDTH + 3,  // +1 for I04b29480233f4def5c875875b6bdc3b1 bit for I352655f17375a62637cdddfd1b812987
parameter SGN_MAX_SUM_WDTH = MAX_SUM_WDTH_L - 1, //Ie86b28b55eaf8feb03e24730be892314 I04b29480233f4def5c875875b6bdc3b1 bit
parameter MAX_SUM_WDTH_L_P1 = 24, //MAX_SUM_WDTH + 3,  // +1 for I04b29480233f4def5c875875b6bdc3b1 bit for I352655f17375a62637cdddfd1b812987
parameter SGN_MAX_SUM_WDTH_P1 = MAX_SUM_WDTH_L_P1 - 1, //Ie86b28b55eaf8feb03e24730be892314 I04b29480233f4def5c875875b6bdc3b1 bit
parameter SUM_LEN= $clog2(NN+1)
) (

input wire [NN-1:0]                  q0_0,
input wire [NN-1:0]                  q0_1,
output wire [NN-1:0]                 final_y_nr_dec,

input wire [MM-1:0]                  exp_syn,
input wire [31:0]                    percent_probability_int,


input wire  [SUM_LEN-1:0]            HamDist_sum_mm,
input wire  [SUM_LEN-1:0]            HamDist_loop,
input wire  [SUM_LEN-1:0]            HamDist_loop_max,
input wire  [SUM_LEN-1:0]            HamDist_loop_percentage,

output reg                           converged_loops_ended,
output reg                           converged_pass_fail,

output reg                           HamDist_cntr_inc_converged_valid,

input wire  [SUM_LEN-1:0]            HamDist_iir1,
input wire  [SUM_LEN-1:0]            HamDist_iir2,
input wire  [SUM_LEN-1:0]            HamDist_iir3,

input wire                           start_dec,
input wire                           iter_start_int,
/* I0c35fcd8aa6b70a1e6a2f67174222bd1 Ifaf61c215f3a90fcc150ac387f759daf I3bc180bd00be2c60a3a5a68e0dd49503 */
input wire                           clr,
/* I0c35fcd8aa6b70a1e6a2f67174222bd1 I18c0d99dcef0c6b3cc1cadd623fdbf9f I3bc180bd00be2c60a3a5a68e0dd49503 */
input wire                           rstn,
input wire                           clk

);

`ifdef ENCRYPT
`endif

reg [NN-1:0]                     tmp_bit;
reg [12-1:0]                     I112f8303dd783640746b7cebaf5bc327;
reg [12-1:0]                     I8ff243fdce9dce8c86b33239c193d9bb;
reg [12-1:0]                     If41bc339aeff21a33c6cb7e4ad526a2d;


wire [MAX_SUM_WDTH_L-1:0]        I43864225be03ea8e9379eb28dfa6c599;
wire [MAX_SUM_WDTH_L-1:0]        I31cb0c699cffcd2fedfbed0e1b86490e;
wire [MAX_SUM_WDTH_L-1:0]        Ibed5004d869a01005768ba694c2234d6;
wire [MAX_SUM_WDTH_L-1:0]        Ia4b2db3d48f946b0bfd0be0e32d7518d;
wire [MAX_SUM_WDTH_L-1:0]        I4d908bbe633c193cd9fc93dd33c60bd2;
wire [MAX_SUM_WDTH_L-1:0]        Ib14733d3585dbf7f196cfc068e9508f0;
wire [MAX_SUM_WDTH_L-1:0]        Idfcf7f3240d92bfc87d44833bc00ff9d;
wire [MAX_SUM_WDTH_L-1:0]        I1cff7306aaf303bb3342ea3d72048908;
wire [MAX_SUM_WDTH_L-1:0]        I26bdcc44692db066911c8d5b0a1aae0c;
wire [MAX_SUM_WDTH_L-1:0]        Id144785da9b171f1e2d0e9182d693e31;
wire [MAX_SUM_WDTH_L-1:0]        I6b7a8ba12de5b44817ec99faebe54617;
wire [MAX_SUM_WDTH_L-1:0]        I4a403449a9ba75243369032e1cca1a0d;
wire [MAX_SUM_WDTH_L-1:0]        If85d9a95c1c02ce2da1dc3486b53eb81;
wire [MAX_SUM_WDTH_L-1:0]        I8e470b68bf35c647af42b6e46201e570;
wire [MAX_SUM_WDTH_L-1:0]        I484ec87270fcc959a486ebce40a9a03c;
wire [MAX_SUM_WDTH_L-1:0]        I079932780612fbce79cbe9b58bb6c2b5;
wire [MAX_SUM_WDTH_L-1:0]        Ibb157b97546cb19fa7c1c0a7c79b1d38;
wire [MAX_SUM_WDTH_L-1:0]        I45cb51c25c426c296f97a5d23a08c063;
wire [MAX_SUM_WDTH_L-1:0]        Iff1d4b06901796098f91e87a3c30f7a5;
wire [MAX_SUM_WDTH_L-1:0]        I16db9cab1981451a02dab21e2ca221b4;
wire [MAX_SUM_WDTH_L-1:0]        I72756ea6a4997bc4afd4bfde1dfb2d26;
wire [MAX_SUM_WDTH_L-1:0]        I2882ae2eb6d79a5b96d1ed937dcfd8bf;
wire [MAX_SUM_WDTH_L-1:0]        I1a632a3e06ad738d5865acc77e204f48;
wire [MAX_SUM_WDTH_L-1:0]        I4d4ec5540257040d10182ed478a71918;
wire [MAX_SUM_WDTH_L-1:0]        I8da7e01f56dc9a70eb6b3f110dc005c2;
wire [MAX_SUM_WDTH_L-1:0]        Icc5d7bcbd7fcdb5092e6d8e18f6de6ec;
wire [MAX_SUM_WDTH_L-1:0]        I83cec264bd378f1dc23f87e439e7310e;
wire [MAX_SUM_WDTH_L-1:0]        Ied7e494fb288f78d110ed06662f1926a;
wire [MAX_SUM_WDTH_L-1:0]        Idd5b362dab4f93bba0c39af78c4c5981;
wire [MAX_SUM_WDTH_L-1:0]        Id033e7adfcfb0420cc592a1fb6c297b6;
wire [MAX_SUM_WDTH_L-1:0]        Iaee91a5e94c3f174682f72a1ebfd0021;
wire [MAX_SUM_WDTH_L-1:0]        I0cd8a6e719305ee3fbe8228081993957;
wire [MAX_SUM_WDTH_L-1:0]        I9b8cfdb69b76453a3ac687a1e098417f;
wire [MAX_SUM_WDTH_L-1:0]        Ic2159627df2efa5e677fa6f4498bdd31;
wire [MAX_SUM_WDTH_L-1:0]        I59fba74472ded0a985cb237104ac127f;
wire [MAX_SUM_WDTH_L-1:0]        Ia526539cc0f844b802d412b7a17cb6a6;
wire [MAX_SUM_WDTH_L-1:0]        I5d80b7c7d102d2c2bfa73a68c73376be;
wire [MAX_SUM_WDTH_L-1:0]        Ia92defa0ca87c7c30fbe901da40a575e;
wire [MAX_SUM_WDTH_L-1:0]        I8fb1602dcdcd2912ea8aec42e2b7848f;
wire [MAX_SUM_WDTH_L-1:0]        I0cedca0e2c589104d6f3318505910594;
wire [MAX_SUM_WDTH_L-1:0]        I54c260db5c1b2c76527c8fc1cee229fe;
wire [MAX_SUM_WDTH_L-1:0]        I3d700e050cb7f22b0e381f3c72a20124;
wire [MAX_SUM_WDTH_L-1:0]        I63c0c8bef1dea4e499a16ce01e781951;
wire [MAX_SUM_WDTH_L-1:0]        Ia8abcb8cf8d9ecc17c27ff015aa0b71f;
wire [MAX_SUM_WDTH_L-1:0]        I3f59174b3764a0b0741462024be9fb92;
wire [MAX_SUM_WDTH_L-1:0]        If0c2d002c315b21e11ae776bb48c9338;
wire [MAX_SUM_WDTH_L-1:0]        I18e548b082364c75686f2b7ad2ef46ab;
wire [MAX_SUM_WDTH_L-1:0]        I5e0d6b44474a226ab2ce916a6d46072a;
wire [MAX_SUM_WDTH_L-1:0]        I0c53d8d6a5b92960e29fc31cf456c23b;
wire [MAX_SUM_WDTH_L-1:0]        Ib16c6096ce80e2f15a5ccea145e28510;
wire [MAX_SUM_WDTH_L-1:0]        I0e7ca2d6470b9bfc6a1ca6143b468507;
wire [MAX_SUM_WDTH_L-1:0]        I4ba05e74c2f63e2f4c59268775d549aa;
wire [MAX_SUM_WDTH_L-1:0]        Iaed26e1c4a2578d16b111d15d31339d2;
wire [MAX_SUM_WDTH_L-1:0]        Ic566fe27ccaf2220101cbc49fc187a6b;
wire [MAX_SUM_WDTH_L-1:0]        Ibf9f6d7baed9e761b69fb41442761ac6;
wire [MAX_SUM_WDTH_L-1:0]        Id5b4ee69444e5b499476c05a7f1d6e60;
wire [MAX_SUM_WDTH_L-1:0]        Id6105518ade80c89d4f20222a2382efb;
wire [MAX_SUM_WDTH_L-1:0]        I26cf25e680483bf4e556d74efec35ee7;
wire [MAX_SUM_WDTH_L-1:0]        I8636f5c91b567780d3324e4b8a320fc2;
wire [MAX_SUM_WDTH_L-1:0]        I914bef0326cf82d350344317eb1359be;
wire [MAX_SUM_WDTH_L-1:0]        I7de222bc26e38b8b6543819701740302;
wire [MAX_SUM_WDTH_L-1:0]        Ie3361a270ebc41698ef4651bb3548a49;
wire [MAX_SUM_WDTH_L-1:0]        I1240c9410b897a4d0504affca5ba139e;
wire [MAX_SUM_WDTH_L-1:0]        If17b4f86674bc5fb212a1f7751fb043a;
wire [MAX_SUM_WDTH_L-1:0]        I275f6334127640b2de3f0f87f54fd74c;
wire [MAX_SUM_WDTH_L-1:0]        Iec844d10736440b96f9d6c651e604efd;
wire [MAX_SUM_WDTH_L-1:0]        Ie04ce30f26a4ef1ee5b34474368dbac7;
wire [MAX_SUM_WDTH_L-1:0]        Ibfee0b4ad5cdf16e88fcf469c5e031e9;
wire [MAX_SUM_WDTH_L-1:0]        I3a4a965f22487553dec2a3e8e7836264;
wire [MAX_SUM_WDTH_L-1:0]        I2a2d014f94d7a3b9fb3024a3e9107a73;
wire [MAX_SUM_WDTH_L-1:0]        I5bab5ae46114c487f67b8e779d7461df;
wire [MAX_SUM_WDTH_L-1:0]        I45373bff54eccf8137da2931d841934e;
wire [MAX_SUM_WDTH_L-1:0]        Ib9322ec1d3866ba3cb42e96b5ff5cfb2;
wire [MAX_SUM_WDTH_L-1:0]        I0a9cb91319cc0d0c1c4d0020cce321d7;
wire [MAX_SUM_WDTH_L-1:0]        I299b37fd45c6ee2031fb2c74caac73be;
wire [MAX_SUM_WDTH_L-1:0]        Ic2f450f7ab60ba57dfc1406c92c0f077;
wire [MAX_SUM_WDTH_L-1:0]        Ieca5b21b91e150c9d509964bdcea500d;
wire [MAX_SUM_WDTH_L-1:0]        I48b39ee498563e23c3a4be079b6100d8;
wire [MAX_SUM_WDTH_L-1:0]        Iac8cb32c2d86b975f51a2ed605002e51;
wire [MAX_SUM_WDTH_L-1:0]        Ic989dc794ce4356856b3916ab1889589;
wire [MAX_SUM_WDTH_L-1:0]        Ie380b37a78242e6d45b659d568887457;
wire [MAX_SUM_WDTH_L-1:0]        Ie43a7f8082f91c2955076a6373028b55;
wire [MAX_SUM_WDTH_L-1:0]        Iea765ae5e9c65b3186445b15c56f69e5;
wire [MAX_SUM_WDTH_L-1:0]        I74b55d2f94073ba8f948e4b02386867c;
wire [MAX_SUM_WDTH_L-1:0]        I015630502f5cb4eb27b2a673e810f1dc;
wire [MAX_SUM_WDTH_L-1:0]        I5085f161323433d8d38be2e4511b0c46;
wire [MAX_SUM_WDTH_L-1:0]        Ie9fd8f7dc0c3849c0437a2a3d8607b4c;
wire [MAX_SUM_WDTH_L-1:0]        I9306d9ef7934ffe5902306b9783c351e;
wire [MAX_SUM_WDTH_L-1:0]        I70e68beb262fbdeba621b3794adf9f84;
wire [MAX_SUM_WDTH_L-1:0]        Ie7bf11bab3d601fd0a6e3eb415e263c8;
wire [MAX_SUM_WDTH_L-1:0]        Ica3d4ebff001fb6ee69a66eb898eb5bd;
wire [MAX_SUM_WDTH_L-1:0]        I27951ef3d612004abdc639662807426b;
wire [MAX_SUM_WDTH_L-1:0]        Ice4f4ba8bb3381c8846941d5d5fe4534;
wire [MAX_SUM_WDTH_L-1:0]        I223151b6414d9979d71023053dd3f5e2;
wire [MAX_SUM_WDTH_L-1:0]        I73d2731c1b1ae5ef73ce0eb9c8995912;
wire [MAX_SUM_WDTH_L-1:0]        I5ca15c7da1f49580ddedd9ff8ba822c0;
wire [MAX_SUM_WDTH_L-1:0]        I8289bfc08a5d8979ec26825bcb6e3d18;
wire [MAX_SUM_WDTH_L-1:0]        Ie3c88bc240576aa220f0f110b13bfdd3;
wire [MAX_SUM_WDTH_L-1:0]        I583c6d23506c7d7b84403bfe977ec1ec;
wire [MAX_SUM_WDTH_L-1:0]        I768afe193d9d79b136736abc6846d945;
wire [MAX_SUM_WDTH_L-1:0]        I277d7065150714e33d8ba64875d18190;
wire [MAX_SUM_WDTH_L-1:0]        Ia5c77c9be26d62b026f24ee5a5e25fb8;
wire [MAX_SUM_WDTH_L-1:0]        I88a325547ccfe4eabf90792abd60e356;
wire [MAX_SUM_WDTH_L-1:0]        I21842d06e25948ef461d1fd03485f86c;
wire [MAX_SUM_WDTH_L-1:0]        Id65f22fa8fc9c47bfd00c796b63c9fa4;
wire [MAX_SUM_WDTH_L-1:0]        I288ff69a7395e74f7de8da5a6a7f9062;
wire [MAX_SUM_WDTH_L-1:0]        I2ba94ef71f97b9ba731b306d4a5fd02c;
wire [MAX_SUM_WDTH_L-1:0]        I26ae9e570a101c6f8237d7941285b924;
wire [MAX_SUM_WDTH_L-1:0]        Icb92c7c10f0bfc5d287228f98d8a235c;
wire [MAX_SUM_WDTH_L-1:0]        Iba4972a3b71a3101ab23190ed905dc17;
wire [MAX_SUM_WDTH_L-1:0]        I33703f538ec70268e6c00ad6eef6c4e0;
wire [MAX_SUM_WDTH_L-1:0]        I71b93abe4b20e6a17ff17e0f33ac2ca5;
wire [MAX_SUM_WDTH_L-1:0]        I91c2f3cdd7cc98a60090ec6e46d52ae7;
wire [MAX_SUM_WDTH_L-1:0]        I4254f2987cd014ed703ae18e9963e585;
wire [MAX_SUM_WDTH_L-1:0]        I9068cca0de6ecff56ca542d0998fcab2;
wire [MAX_SUM_WDTH_L-1:0]        Ib3ec015a3d43d46e0b7142b21a81cfee;
wire [MAX_SUM_WDTH_L-1:0]        I8cb171677016e4309034dc5d83981a48;
wire [MAX_SUM_WDTH_L-1:0]        I2a4b3573ae7c3b38ec34591f20c1d076;
wire [MAX_SUM_WDTH_L-1:0]        I276c2ce5d3a1b7551c2790971071b094;
wire [MAX_SUM_WDTH_L-1:0]        I9dff504e40aaddefedbb7b0f822c844a;
wire [MAX_SUM_WDTH_L-1:0]        I4ed5da534afbfe9ecbc10ef4cc649a55;
wire [MAX_SUM_WDTH_L-1:0]        I618363a8ac413dd0ee52eb658940eaed;
wire [MAX_SUM_WDTH_L-1:0]        I54166b387c02e12374d6febc425bfb7a;
wire [MAX_SUM_WDTH_L-1:0]        I0b6cdfa1dbfa774fc9a12d856e61cddb;
wire [MAX_SUM_WDTH_L-1:0]        Ic4af6c9097257c9b22a57ce4b79b40fe;
wire [MAX_SUM_WDTH_L-1:0]        Iae21bdea20a6266d3f69aa680b6b2817;
wire [MAX_SUM_WDTH_L-1:0]        I37e360420c7dd061de93a6647513676d;
wire [MAX_SUM_WDTH_L-1:0]        Ia81c31ea4f4786136b539c9766987596;
wire [MAX_SUM_WDTH_L-1:0]        I5a4f0749acdc34fd0786e4b3d062f88b;
wire [MAX_SUM_WDTH_L-1:0]        I5529d6db17b6184c45cc4487e5a2c24a;
wire [MAX_SUM_WDTH_L-1:0]        Iabe5aea929c668c9b9728d073ffb00c8;
wire [MAX_SUM_WDTH_L-1:0]        I4fb3fe065daa2708e55c812e57c19fb6;
wire [MAX_SUM_WDTH_L-1:0]        I4bd98e902e805426fdd4606fcb5a5214;
wire [MAX_SUM_WDTH_L-1:0]        Ia5e26c2417aba1005971749f4ab2f367;
wire [MAX_SUM_WDTH_L-1:0]        I0e112f1d4e9c934a118f79f3856744a9;
wire [MAX_SUM_WDTH_L-1:0]        I005e8b590924f9486cb23191d35c9797;
wire [MAX_SUM_WDTH_L-1:0]        I8c5f98353b5b082dc3cf056469945a08;
wire [MAX_SUM_WDTH_L-1:0]        I9aa11f30712f1779339b985212a7979c;
wire [MAX_SUM_WDTH_L-1:0]        I65928407b1d5447dbc815cd2d2e7b37d;
wire [MAX_SUM_WDTH_L-1:0]        If5b3850da967f6f3d7a71d680341ad1c;
wire [MAX_SUM_WDTH_L-1:0]        I0aa5522190c741b7df4c4d7d34e46987;
wire [MAX_SUM_WDTH_L-1:0]        Iff777b2c4a3939e330c4cbb36cbe1ac5;
wire [MAX_SUM_WDTH_L-1:0]        I2d839c10960739097d449efab58b9fd4;
wire [MAX_SUM_WDTH_L-1:0]        Ice8765807beffd3acf59fa137ee0baac;
wire [MAX_SUM_WDTH_L-1:0]        I529eaa7e5eeb6d0a1aba78df5d5a2fa0;
wire [MAX_SUM_WDTH_L-1:0]        Icb2805685607d5fedd0300c9d800f863;
wire [MAX_SUM_WDTH_L-1:0]        Idadf072247b351cf51d718f797c3b375;
wire [MAX_SUM_WDTH_L-1:0]        I6fcb3b133a6a654b69f41468a713d922;
wire [MAX_SUM_WDTH_L-1:0]        I77e1f5f504a794edbb89c66cf1ffcf66;
wire [MAX_SUM_WDTH_L-1:0]        I185085cbf8da6df921ba32442b28bcca;
wire [MAX_SUM_WDTH_L-1:0]        Ibcb80df5bed66f8498561e3f3ffa4ec4;
wire [MAX_SUM_WDTH_L-1:0]        I2cf5304a672431888916e08b3c15f0c7;
wire [MAX_SUM_WDTH_L-1:0]        Icf266f710358631b7119ef526acb301c;
wire [MAX_SUM_WDTH_L-1:0]        Ia209e5b03deaf4fcb8ae12b731a49e0a;
wire [MAX_SUM_WDTH_L-1:0]        Iffb7fe9c74dfc01a43e99a099c4e7e04;
wire [MAX_SUM_WDTH_L-1:0]        I43f52bcba1bd2e8ee5fac03320e4f19f;
wire [MAX_SUM_WDTH_L-1:0]        I9fdfe73e77c384d33196c0f2d2a2fde2;
wire [MAX_SUM_WDTH_L-1:0]        I546657528d591e8bb44c32fed7707af5;
wire [MAX_SUM_WDTH_L-1:0]        I6e4ae763dc4e8aa8afc4599de96c75d3;
wire [MAX_SUM_WDTH_L-1:0]        Id8c36004ae8e550569a491f6b514945a;
wire [MAX_SUM_WDTH_L-1:0]        I111ac0aadbdd3e4479ca0786491a7b08;
wire [MAX_SUM_WDTH_L-1:0]        Ib83242b57ab050b0e5f9bdf91fa118fb;
wire [MAX_SUM_WDTH_L-1:0]        I7be8b2f8a9fe8e13001c2a1fce4a8a3f;
wire [MAX_SUM_WDTH_L-1:0]        If4d030e5858f325debc6f37abf4a7d6c;
wire [MAX_SUM_WDTH_L-1:0]        I627e4bdc8061c69e3fcac17535b9f1e0;
wire [MAX_SUM_WDTH_L-1:0]        Ia443284a35e0873de59b3ae55b7f809d;
wire [MAX_SUM_WDTH_L-1:0]        Ibafedcf9f2990ed9c1efa973a0b1d81d;
wire [MAX_SUM_WDTH_L-1:0]        I439c7c302b535bfd7db655c3c607d71f;
wire [MAX_SUM_WDTH_L-1:0]        I2133d362ba45ceb3dceaa84e95ace1e6;
wire [MAX_SUM_WDTH_L-1:0]        I67534b68fee8f76ac0c5e64cd02aba42;
wire [MAX_SUM_WDTH_L-1:0]        I8613cac4ccd4f956e8a0ae7b627f5be2;
wire [MAX_SUM_WDTH_L-1:0]        I8493e2dac01f009db1d2d5504b49d135;
wire [MAX_SUM_WDTH_L-1:0]        I5c278aad08b7c4b0237d68f88fcb3f3a;
wire [MAX_SUM_WDTH_L-1:0]        Iba75ff0f3b67c7e28cf627706733d528;
wire [MAX_SUM_WDTH_L-1:0]        I9164fa2a9a33da6612ea692cf3fa7d2f;
wire [MAX_SUM_WDTH_L-1:0]        I0f3c4fb63ef1e88168b4d28175a0b68c;
wire [MAX_SUM_WDTH_L-1:0]        I99d236d41be79090ca7ba1fb6faaec4c;
wire [MAX_SUM_WDTH_L-1:0]        I487b9b236d118786e475ccc5e4e56a6d;
wire [MAX_SUM_WDTH_L-1:0]        I6cb09ac924c3b3b44443263e08c3315c;
wire [MAX_SUM_WDTH_L-1:0]        Id924dafd31fd0af0b28c7e6b7e95ec37;
wire [MAX_SUM_WDTH_L-1:0]        I9184110e3e9b8614460fc0abe5fff2d9;
wire [MAX_SUM_WDTH_L-1:0]        If8865fee7dbf593b34ea54692d947f10;
wire [MAX_SUM_WDTH_L-1:0]        I4854ff71aa885da3d07acaaa24740d7c;
wire [MAX_SUM_WDTH_L-1:0]        Ie8befb003fe83e774e8d1d01d4e2f4ad;
wire [MAX_SUM_WDTH_L-1:0]        Ie7e196fbb66ba6bee51ef0064ca519c2;
wire [MAX_SUM_WDTH_L-1:0]        I685699f60c76b00df87c9c53e9a8e448;
wire [MAX_SUM_WDTH_L-1:0]        Ib6c0e635e659f54724737f0cffd1b0fc;
wire [MAX_SUM_WDTH_L-1:0]        I3a8bcfdab631a268d21c87b98e9d1c49;
wire [MAX_SUM_WDTH_L-1:0]        I3faeba79f7af7a006ab5cd256352e2db;
wire [MAX_SUM_WDTH_L-1:0]        I02e672436ade3ee620c72c0d9ceee664;
wire [MAX_SUM_WDTH_L-1:0]        I65708fb59e90bb79b8107da619fe63eb;
wire [MAX_SUM_WDTH_L-1:0]        I840a1a7c0bf49f4f42499b33f32fa02d;
wire [MAX_SUM_WDTH_L-1:0]        If7543e2f5a158b1f3f3a4078ec54cab5;
wire [MAX_SUM_WDTH_L-1:0]        I98a2aa729628adde0b6047869bd12743;
wire [MAX_SUM_WDTH_L-1:0]        Ibfb57f2b507c27759a3556759f23977b;
wire [MAX_SUM_WDTH_L-1:0]        Ib20dec1346f227042c749ec1abfa4d39;
wire [MAX_SUM_WDTH_L-1:0]        Ifba318d4faf308168c5eac8fe92395b4;
wire [MAX_SUM_WDTH_L-1:0]        I95b923444062b4a98918c685c65996d0;
wire [MAX_SUM_WDTH_L-1:0]        I45a6ef43e6e42594444adcbda26700ab;
wire [MAX_SUM_WDTH_L-1:0]        I508cea40d87bec2672f980d145c89b55;
wire [MAX_SUM_WDTH_L-1:0]        I0ace1d51fdee91f8f3826a945c4e66a4;
wire [MAX_SUM_WDTH_L-1:0]        I99ff3922e018c409dc8ce5f3503e3c56;
wire [MAX_SUM_WDTH_L-1:0]        I6a3824a6598bbaa138e1e763ad85f5f7;
wire [MAX_SUM_WDTH_L-1:0]        I283107989a436e2c720123b8d9e335c2;
wire [MAX_SUM_WDTH_L-1:0]        I7b12345fe53174cadef6811fb8869b42;
wire [MAX_SUM_WDTH_L-1:0]        Iac6fcccf3a0cfe04edc0d998b60c2681;
wire [MAX_SUM_WDTH_L-1:0]        Ic9678deca4bf44a7b99f853334f6a05c;
wire [MAX_SUM_WDTH_L-1:0]        Ie40c90fdb38b3e4046ba89295ed77d7c;
wire [MAX_SUM_WDTH_L-1:0]        Iea4a7766d3b9d5d030ade1739859ef0d;
wire [MAX_SUM_WDTH_L-1:0]        I844b9a89ffb7a5e48979fdea546e244a;
wire [MAX_SUM_WDTH_L-1:0]        I656852be6f5b3542862e0f68d48be518;
wire [MAX_SUM_WDTH_L-1:0]        Id6551b6b053952162b90792ab73a1a49;
wire [MAX_SUM_WDTH_L-1:0]        Ib7fde6a2ec1ff0a3af10bccf3012e63f;
wire [MAX_SUM_WDTH_L-1:0]        I989091b3586964ab598f166a89279d16;
wire [MAX_SUM_WDTH_L-1:0]        I9785922874bba479ce4a9bf1759e2933;
wire [MAX_SUM_WDTH_L-1:0]        Ifbaae8b3da03911a4c96d4efdb9283c5;
wire [MAX_SUM_WDTH_L-1:0]        I77a54091bc2c3d9006ecb3471b94d8c8;
wire [MAX_SUM_WDTH_L-1:0]        I9859b94cda465ceaaa5674eb19e94824;
wire [MAX_SUM_WDTH_L-1:0]        I5a7746e9fbb8c009f83ae57423296cdf;
wire [MAX_SUM_WDTH_L-1:0]        Ibddcc2e26fba20dfe2a2d399be2bc45b;
wire [MAX_SUM_WDTH_L-1:0]        I8dbe6497a8deabcc60783bfe7548d0fb;
wire [MAX_SUM_WDTH_L-1:0]        Ifef870b405335975988b58b2273d4e1a;
wire [MAX_SUM_WDTH_L-1:0]        Ic1f6842b4f246d624d91daa6ada10ca9;
wire [MAX_SUM_WDTH_L-1:0]        Ibc8679379ddc43ee4bc508a1f577eb2c;
wire [MAX_SUM_WDTH_L-1:0]        Ibdd9957b7f1a319b797c021933ff75d7;
wire [MAX_SUM_WDTH_L-1:0]        I041f9455435bfa375395eb330a34993d;
wire [MAX_SUM_WDTH_L-1:0]        Ifbe29365e7035c78af9f42902b0d303e;
wire [MAX_SUM_WDTH_L-1:0]        Ic8759e2f58848b33082bd1b02acc9c0b;
wire [MAX_SUM_WDTH_L-1:0]        Ie2e3d64640c339dc51512979dbd6a173;
wire [MAX_SUM_WDTH_L-1:0]        Ib2c327648cce481482eaf0467e9227d4;
wire [MAX_SUM_WDTH_L-1:0]        I535cad8c919a4330257eb5b4bed61b3a;
wire [MAX_SUM_WDTH_L-1:0]        Ib2afdf9534deaae465d99b7e377788bb;
wire [MAX_SUM_WDTH_L-1:0]        I6eaffd980e4d77fdbda5e63bad9489d7;
wire [MAX_SUM_WDTH_L-1:0]        I6e4786234b286b12c83e06e93c628534;
wire [MAX_SUM_WDTH_L-1:0]        Idcc745602c4b7b34df9c3d68f9a9d76d;
wire [MAX_SUM_WDTH_L-1:0]        I0fc42ce9cc31d781ea3013318c25a571;
wire [MAX_SUM_WDTH_L-1:0]        I4363ca6b3d9ca9863f70958aa7c23777;
wire [MAX_SUM_WDTH_L-1:0]        Ic902e09b33db1b919c102f7971cdef7b;
wire [MAX_SUM_WDTH_L-1:0]        Icf4405d4a4063448a2be8ad0354ab1a8;
wire [MAX_SUM_WDTH_L-1:0]        I72108531a608f6d5e51a481c68d7b271;
wire [MAX_SUM_WDTH_L-1:0]        I6922b510e432e06d209095bcc6297e7e;
wire [MAX_SUM_WDTH_L-1:0]        Ief90f8a8efca2b06eff0d4cba1cbb342;
wire [MAX_SUM_WDTH_L-1:0]        Ib5334df42ee8f1574e41cb30b903fae9;
wire [MAX_SUM_WDTH_L-1:0]        I535b29f7177b4fc009ee998f1f4f7d7f;
wire [MAX_SUM_WDTH_L-1:0]        Id0842da8068ee88d99af7acea50e7b77;
wire [MAX_SUM_WDTH_L-1:0]        Ib6cdbbb765694d822639b7c8fbfc50c4;
wire [MAX_SUM_WDTH_L-1:0]        Ibdaa6d215d34aa0cc27d5234da6fd991;
wire [MAX_SUM_WDTH_L-1:0]        Id769d4a92f5f6da262ce0521e5509368;
wire [MAX_SUM_WDTH_L-1:0]        Iaf3a0b5ea5d9eda47fcced9260922bc6;
wire [MAX_SUM_WDTH_L-1:0]        I03a8a458ee0942c35001cbfe8e589222;
wire [MAX_SUM_WDTH_L-1:0]        I25eb943ea517a4827efb1e797bfdc4f5;
wire [MAX_SUM_WDTH_L-1:0]        Iac4b8906947fc90bfe76cee2f1d4c4ab;
wire [MAX_SUM_WDTH_L-1:0]        I58a490344f87b4d5bb319e3e85ba9278;
wire [MAX_SUM_WDTH_L-1:0]        I9222c4c0eb2b110fd80547d46ba17036;
wire [MAX_SUM_WDTH_L-1:0]        Ic1af7410a9d11c5324f3ee5b2e0e9dac;
wire [MAX_SUM_WDTH_L-1:0]        I9e0a36d0be66b4c02b03e5b75b686226;
wire [MAX_SUM_WDTH_L-1:0]        I1eef40a71c8d1e2da9802929a5347e90;
wire [MAX_SUM_WDTH_L-1:0]        Ied41909cd443432dafadba42672151c1;
wire [MAX_SUM_WDTH_L-1:0]        Ib2c1636a66f6479d6123a038cbc668d5;
wire [MAX_SUM_WDTH_L-1:0]        Ica02d19b129c8b1d491ea4747a55113e;
wire [MAX_SUM_WDTH_L-1:0]        I31bf4597a3b776962f5c820378254065;
wire [MAX_SUM_WDTH_L-1:0]        I58361fb97f1b5aff0a2751d35c8da672;
wire [MAX_SUM_WDTH_L-1:0]        I8ab7efc436a0f2cc3efbc299a0ddf914;
wire [MAX_SUM_WDTH_L-1:0]        I3934ed7170967ff3852944cc39ba1de9;
wire [MAX_SUM_WDTH_L-1:0]        Ic690477b1672dea4905a5e1c92b47366;
wire [MAX_SUM_WDTH_L-1:0]        I5eaa11e26f19b94dcb7eaee7f09d24b4;
wire [MAX_SUM_WDTH_L-1:0]        Iaf1d3be13e6441a7a9ab3f286a7dc21b;
wire [MAX_SUM_WDTH_L-1:0]        I61f5ebea2bbe443b644c95ee559c2234;
wire [MAX_SUM_WDTH_L-1:0]        I1fbcaf2f6be01b129ebc24dee8a65396;
wire [MAX_SUM_WDTH_L-1:0]        I1c0df8c2c64b688ae417a238263f33db;
wire [MAX_SUM_WDTH_L-1:0]        I4f169c2c8c0768f2725ed655a03acfc2;
wire [MAX_SUM_WDTH_L-1:0]        I96f65790e2cacf7b529ce5b88598da00;
wire [MAX_SUM_WDTH_L-1:0]        I6b5720d71a0b4cd10ea34affa6631a25;
wire [MAX_SUM_WDTH_L-1:0]        Ifc7eec6765af08463751db128f8818b3;
wire [MAX_SUM_WDTH_L-1:0]        I8dddcade21ad3bb330c1c25970c32b73;
wire [MAX_SUM_WDTH_L-1:0]        I74a7b85ddacad06ab1c6b0db9b084bd3;
wire [MAX_SUM_WDTH_L-1:0]        I2b0b168ce4fe8aa4a2e7cb69fe532aa3;
wire [MAX_SUM_WDTH_L-1:0]        I3e8d26ea83937cae01aadf1092c59bdf;
wire [MAX_SUM_WDTH_L-1:0]        I90a4190941651d885d04deb86a163365;
wire [MAX_SUM_WDTH_L-1:0]        I7d85b73e85379bf3a480e954c05516f3;
wire [MAX_SUM_WDTH_L-1:0]        Id5c9a9b9c34c8f9d56df0aa8d780c9d3;
wire [MAX_SUM_WDTH_L-1:0]        I21255a0ad20a9668c958faf68d53b2bc;
wire [MAX_SUM_WDTH_L-1:0]        Ifba1584d599da13b98a3b76b4db10974;
wire [MAX_SUM_WDTH_L-1:0]        Iad0f4602ec545dc6ef12aa34add00ed3;
wire [MAX_SUM_WDTH_L-1:0]        I8bb46c3eb9f54c5d1b28dc6aa0154358;
wire [MAX_SUM_WDTH_L-1:0]        Ic09b4671e867144fe9f54a09e74c5519;
wire [MAX_SUM_WDTH_L-1:0]        I391a2f354262558ff17d7d80b8c39e8c;
wire [MAX_SUM_WDTH_L-1:0]        If6b40a030cb120fe017bf9d39e1a35d1;
wire [MAX_SUM_WDTH_L-1:0]        I490996026af34eba5bcd8d553af818eb;
wire [MAX_SUM_WDTH_L-1:0]        Icbc12ab47f586b12402ae5d4361c967d;
wire [MAX_SUM_WDTH_L-1:0]        Iee0e45914c52a357e1e32922299d6937;
wire [MAX_SUM_WDTH_L-1:0]        Iefe423653d454e21324a6857b52f98ac;
wire [MAX_SUM_WDTH_L-1:0]        I6d6a242cdfadfc97fe656510bef73adc;
wire [MAX_SUM_WDTH_L-1:0]        Ib5c8d91204a2d313c9c23110a53cd0cf;
wire [MAX_SUM_WDTH_L-1:0]        Ic9740baafb1c92e3a25f0a1e7bc46486;
wire [MAX_SUM_WDTH_L-1:0]        I6f69796a6fe6da57066319ec8210c1a3;
wire [MAX_SUM_WDTH_L-1:0]        Idb862697f62a6c678072de760e176096;
wire [MAX_SUM_WDTH_L-1:0]        I06e05a1ed002175a75d02b8b76f52c50;
wire [MAX_SUM_WDTH_L-1:0]        I1e110e27162231650875dd1152d96e64;
wire [MAX_SUM_WDTH_L-1:0]        Ic46357bb77f6183329946f7e28294365;
wire [MAX_SUM_WDTH_L-1:0]        I8741c5cc763512d16cb1186fa3323f45;
wire [MAX_SUM_WDTH_L-1:0]        I30b5c7aadb5312ce96e833704bb3a320;
wire [MAX_SUM_WDTH_L-1:0]        If404a00ab81d6ebbc0dbdf4aecdce389;
wire [MAX_SUM_WDTH_L-1:0]        I19875f52f79482b477f1febaa7e97090;
wire [MAX_SUM_WDTH_L-1:0]        Ic7855ca956651bd368cbdde7ec93ba6d;
wire [MAX_SUM_WDTH_L-1:0]        Ic57a2627a194099105a2908a41feddfb;
wire [MAX_SUM_WDTH_L-1:0]        I4d1ba6ee8fb9505ba3b58b2b7553245b;
wire [MAX_SUM_WDTH_L-1:0]        Ieb7b388ff89e352dd239e0ccbe7b9ecc;
wire [MAX_SUM_WDTH_L-1:0]        Ib1461f456ebc14f449eee77e386a4c69;
wire [MAX_SUM_WDTH_L-1:0]        I8786eb767f02164cdc32f14f41b5d0e1;
wire [MAX_SUM_WDTH_L-1:0]        Id6fa8ec5d1062fc3e09bdac65ff79f45;
wire [MAX_SUM_WDTH_L-1:0]        I83b77ad1a40dc102f28153f692516eb4;
wire [MAX_SUM_WDTH_L-1:0]        I55e54359961ef6e5a63f1c2eb0ad4aa1;
wire [MAX_SUM_WDTH_L-1:0]        I90001da8c360ccff128f637cd672ad42;
wire [MAX_SUM_WDTH_L-1:0]        Ib38a46dc131d635b81fb7c196110fc4b;
wire [MAX_SUM_WDTH_L-1:0]        I926c049036f53f0a0a6ad369de116c57;
wire [MAX_SUM_WDTH_L-1:0]        Iac48d2ccf6c6e0c555e874ae77123f2e;
wire [MAX_SUM_WDTH_L-1:0]        Ic6f40833f5f6284c9015304fd3fc00f0;
wire [MAX_SUM_WDTH_L-1:0]        I3f2507530dd648814af0964f7da11d35;
wire [MAX_SUM_WDTH_L-1:0]        Id9edc6ac95a260bf5af3de25f00e9e9c;
wire [MAX_SUM_WDTH_L-1:0]        I28fa295ebd90c2b7255d48ca9ffcfcf3;
wire [MAX_SUM_WDTH_L-1:0]        Ia308e09137af1cb50167562efb5da628;
wire [MAX_SUM_WDTH_L-1:0]        I5aa85d9503b0e4ff46bbd63e873053ca;
wire [MAX_SUM_WDTH_L-1:0]        I7ea8fe50c45e213f3257060e2813240b;
wire [MAX_SUM_WDTH_L-1:0]        Ic3e6e38a2986c7f14fd0db2246367a1c;
wire [MAX_SUM_WDTH_L-1:0]        I581eb136fdd08302e02c1fafb5d5c90b;
wire [MAX_SUM_WDTH_L-1:0]        I080832c25509f7003ed50d71210bc7f7;
wire [MAX_SUM_WDTH_L-1:0]        Ib43383830037df764b48c637a28ab6b5;
wire [MAX_SUM_WDTH_L-1:0]        Iddf65ccb4396288264a400ba37cbb655;
wire [MAX_SUM_WDTH_L-1:0]        Ia7673d73f0535906a99d6cb467892104;
wire [MAX_SUM_WDTH_L-1:0]        I8bc3210e86a523accdbeefe7e72ee4fc;
wire [MAX_SUM_WDTH_L-1:0]        Ib63574478126e6ee30a388d9648cb548;
wire [MAX_SUM_WDTH_L-1:0]        Ic4501a8a1fb34c30a97e18a0ab189e3a;
wire [MAX_SUM_WDTH_L-1:0]        I2b807c16cfc6d65cb2a7f28ffa837974;
wire [MAX_SUM_WDTH_L-1:0]        I0aa93075086164fdbab3814d60633141;
wire [MAX_SUM_WDTH_L-1:0]        I886750aaf8d2040c3f12ff113294f658;
wire [MAX_SUM_WDTH_L-1:0]        I103ec7cf279f527fc6e3648a19a12a8a;
wire [MAX_SUM_WDTH_L-1:0]        I9a57f2f03cf8a154c3a7d48ec089306d;
wire [MAX_SUM_WDTH_L-1:0]        I9d8f8c1792427975a9e7024041f59be9;
wire [MAX_SUM_WDTH_L-1:0]        Ie8644d7edbadf19937c399cf275946e5;
wire [MAX_SUM_WDTH_L-1:0]        I2b32537c9178028493af165398a60875;
wire [MAX_SUM_WDTH_L-1:0]        If06a1563b9d7348de03a98d31bd85b06;
wire [MAX_SUM_WDTH_L-1:0]        I58a7c7b05b84d292cd06d68e96ecb9f8;
wire [MAX_SUM_WDTH_L-1:0]        I3fdec80112b3fc543b217d1c253406da;
wire [MAX_SUM_WDTH_L-1:0]        Ia1aedd38250e76763aaee3de2f832b3c;
wire [MAX_SUM_WDTH_L-1:0]        I2087576fbc15119bf5d9e8afa2603b69;
wire [MAX_SUM_WDTH_L-1:0]        I7a6ab9e700bd94208ab6528af413f3a9;
wire [MAX_SUM_WDTH_L-1:0]        I4481555c402ba99bee05658ba6017984;
wire [MAX_SUM_WDTH_L-1:0]        Ib849494e5087777f646ee0947b4f634a;
wire [MAX_SUM_WDTH_L-1:0]        I18d0dd7a10d6533f721a2392d4ad2d02;
wire [MAX_SUM_WDTH_L-1:0]        Ib8603cb82ceb97c2f35bf8209306a457;
wire [MAX_SUM_WDTH_L-1:0]        I2418ae211f327ed45cc70c42078180dc;
wire [MAX_SUM_WDTH_L-1:0]        I6521c9167261db6eb37f50b66159ddb7;
wire [MAX_SUM_WDTH_L-1:0]        I920f95bb52cdc9b07f93afc3a6b5c009;
wire [MAX_SUM_WDTH_L-1:0]        Iad0ecc5208263d239e4a62c5563f52ab;
wire [MAX_SUM_WDTH_L-1:0]        I0c0be3347a7df9cc39997208b013f17b;
wire [MAX_SUM_WDTH_L-1:0]        I70dc03a46e1ac0da826388abd3bdc503;
wire [MAX_SUM_WDTH_L-1:0]        I452ba61d5fb5c7ead1824dade4bd7801;
wire [MAX_SUM_WDTH_L-1:0]        I8b5d10c412daccdcb07645bf239d61bd;
wire [MAX_SUM_WDTH_L-1:0]        I9b1390839ee2b9ba591e3873e967c8e2;
wire [MAX_SUM_WDTH_L-1:0]        I17e818b67440efaba9a5d19e7467bf85;
wire [MAX_SUM_WDTH_L-1:0]        Ifa67d343acc6f3ec50c2b01fc26b4374;
wire [MAX_SUM_WDTH_L-1:0]        If0676ef300628c4097565b13ef2d8854;
wire [MAX_SUM_WDTH_L-1:0]        I8d26e73fafa909f1e26e329828cf4888;
wire [MAX_SUM_WDTH_L-1:0]        If29fcea810adbdb1c4d8a4ace1d8081b;
wire [MAX_SUM_WDTH_L-1:0]        I0e3286fca6cd040758950259ab663df7;
wire [MAX_SUM_WDTH_L-1:0]        I696db0b98e27dcc4657dc7feb23a881b;
wire [MAX_SUM_WDTH_L-1:0]        I06c0921675f464807a63c7965796f0d0;
wire [MAX_SUM_WDTH_L-1:0]        If36016df78d833c80e1355151c038225;
wire [MAX_SUM_WDTH_L-1:0]        I0dbf900b4f430b4c1106aa86b640bb37;
wire [MAX_SUM_WDTH_L-1:0]        Ib8664a2abe9d6326d6e45bb2a7ad59d0;
wire [MAX_SUM_WDTH_L-1:0]        I91893028c4409cfeceeb7976815b2d31;
wire [MAX_SUM_WDTH_L-1:0]        I2e14fb1e667e967ab4c116e0c7438aec;
wire [MAX_SUM_WDTH_L-1:0]        I0fb60c4f56f6d7b4007cf0dae39f4573;
wire [MAX_SUM_WDTH_L-1:0]        I24b4c998d19ae97f7178e37f75c77d06;
wire [MAX_SUM_WDTH_L-1:0]        Idb73eba1bd4ce25a6109e296f51e7dc4;
wire [MAX_SUM_WDTH_L-1:0]        Ibc1a16427d8dfa5ee20dac15327a53ea;
wire [MAX_SUM_WDTH_L-1:0]        I0e52c25aa840402d944cbd81f73c1ffe;
wire [MAX_SUM_WDTH_L-1:0]        Id7619819e1297844d92c8bf3a1d61926;
wire [MAX_SUM_WDTH_L-1:0]        Idfa432a87877e1ce103e56891745b62a;
wire [MAX_SUM_WDTH_L-1:0]        I13b9e098622d90a1074f636d8f351aca;
wire [MAX_SUM_WDTH_L-1:0]        I78e1205de9119fac3ae8f43c72ac71f4;
wire [MAX_SUM_WDTH_L-1:0]        I5bbbc4eedb7c61516769f429a8498ea7;
wire [MAX_SUM_WDTH_L-1:0]        Ia1d9dee7a9821283498d17de0cfacb32;
wire [MAX_SUM_WDTH_L-1:0]        Idd8643af2515f65fd9a1dfe66494ccf2;
wire [MAX_SUM_WDTH_L-1:0]        I1684820afb9d9cec38cfdfcd6ca8b36a;
wire [MAX_SUM_WDTH_L-1:0]        Ice8a82bdd966719098a8d5f2a826f73d;
wire [MAX_SUM_WDTH_L-1:0]        I338400586daa58006c0a3dcd82ea8f4a;
wire [MAX_SUM_WDTH_L-1:0]        Ie467c5fde1d123da4e9587b5a56748a0;
wire [MAX_SUM_WDTH_L-1:0]        Ifc52604a4f9f9de392a35f2f9fe885b8;
wire [MAX_SUM_WDTH_L-1:0]        I20c4e393929b875521e5316f4d8e2d42;
wire [MAX_SUM_WDTH_L-1:0]        I064499f0315fbeec7b6cb50583388a07;
wire [MAX_SUM_WDTH_L-1:0]        I894ef04bfa1b7b39ef51b7c82f7686eb;
wire [MAX_SUM_WDTH_L-1:0]        I8d6927b0bcbbb318cf52987c121a07b5;
wire [MAX_SUM_WDTH_L-1:0]        Ie0ce2826fd13b0e0b23c91e97787691f;
wire [MAX_SUM_WDTH_L-1:0]        I7dbd1aeba00bb8b257990b7bb294211f;
wire [MAX_SUM_WDTH_L-1:0]        Id5ddf5331aba567aaf5b7eb88b31a52e;
wire [MAX_SUM_WDTH_L-1:0]        I0f46a17f14ab18e6338aa3d06678b0a5;
wire [MAX_SUM_WDTH_L-1:0]        If1ec4241fd12255369f72b3f3310b6e7;
wire [MAX_SUM_WDTH_L-1:0]        Iedf37dac8b3a5331277ae4f0176968aa;
wire [MAX_SUM_WDTH_L-1:0]        Ia422fbdf8f318ff3ddc049d1374e7939;
wire [MAX_SUM_WDTH_L-1:0]        I9cbe73d708c561d43d05945552d32dde;
wire [MAX_SUM_WDTH_L-1:0]        I7e36dcae438a712fca2320117b7e3356;
wire [MAX_SUM_WDTH_L-1:0]        I0f9bc36c9d40290f83489aac3d674924;
wire [MAX_SUM_WDTH_L-1:0]        I3a09554ca009781e28ef1b3ea70d39ad;
wire [MAX_SUM_WDTH_L-1:0]        I28ea268c5b51ac1d9249e96599bb6b0d;
wire [MAX_SUM_WDTH_L-1:0]        I1d648ed8f07f0743a6d616584270c513;
wire [MAX_SUM_WDTH_L-1:0]        I82a225237aeb1ceb31e8cd18b1e45c6f;
wire [MAX_SUM_WDTH_L-1:0]        I36ed1a0d0d618f90443fbea17b7c97ec;
wire [MAX_SUM_WDTH_L-1:0]        I612a41511db375f10f3c2b10d13edb24;
wire [MAX_SUM_WDTH_L-1:0]        I19032091a26dfdfffff60818041ec79e;
wire [MAX_SUM_WDTH_L-1:0]        I6aba8ca0e4b20a6355b43a70f19d9d8c;
wire [MAX_SUM_WDTH_L-1:0]        I839895c8614ff28df83314c44824900b;
wire [MAX_SUM_WDTH_L-1:0]        I8cbafa797ef136d7e50c909dc160deb1;
wire [MAX_SUM_WDTH_L-1:0]        Ibac0851ce1a3c23f18b072d263afff36;
wire [MAX_SUM_WDTH_L-1:0]        Id58474582f209a3859f65a447fe99191;
wire [MAX_SUM_WDTH_L-1:0]        Ic9e06a355beabfacc053ec48f17f49de;
wire [MAX_SUM_WDTH_L-1:0]        I77fd8001d879fc9e9117464fba27902d;
wire [MAX_SUM_WDTH_L-1:0]        I2a0dc4ed573a544cb13544e049514903;
wire [MAX_SUM_WDTH_L-1:0]        I71bc7271cc432bb3c5d0b7a416cdfc60;
wire [MAX_SUM_WDTH_L-1:0]        Ib76e892d1a1271844338042381b5690b;
wire [MAX_SUM_WDTH_L-1:0]        Icb158c031d434cb419c15e0510511231;
wire [MAX_SUM_WDTH_L-1:0]        I563802213afb6abe2f6e8c6f4d1e5b08;
wire [MAX_SUM_WDTH_L-1:0]        Ia5b779ef95333736b08f63770900e275;
wire [MAX_SUM_WDTH_L-1:0]        Ic1120eb027841908cd64fe5c7274da14;
wire [MAX_SUM_WDTH_L-1:0]        I5160de2c5ce4782d8f8be10dc740694b;
wire [MAX_SUM_WDTH_L-1:0]        I5f7b6e6a30348ae86057f7e56f625846;
wire [MAX_SUM_WDTH_L-1:0]        I9de41d0b279b84366640880dbd18c502;
wire [MAX_SUM_WDTH_L-1:0]        Ifec9abca21cf476b70e0befa3926b46a;
wire [MAX_SUM_WDTH_L-1:0]        Ifc527b6af9486df7f52d7eb9637c671f;
wire [MAX_SUM_WDTH_L-1:0]        I31d94aae2e3721045fe850d84dd2225a;
wire [MAX_SUM_WDTH_L-1:0]        If3bdbb4c20efca0c5af78614b4271ed1;
wire [MAX_SUM_WDTH_L-1:0]        I4037f1b207aa101f354e59eddd7c9eb4;
wire [MAX_SUM_WDTH_L-1:0]        If4d63635a5f99c4dc9e5b57712830c20;
wire [MAX_SUM_WDTH_L-1:0]        I1f1f2fefd3381ee48ab0ec9c9301754b;
wire [MAX_SUM_WDTH_L-1:0]        Iba52b84e6e215842e0ca8e72c42ebce7;
wire [MAX_SUM_WDTH_L-1:0]        I597c3f5c14e235f90dc8c796bc3e931d;
wire [MAX_SUM_WDTH_L-1:0]        I397a69dab323c7148b620dd6fe0b0c51;
wire [MAX_SUM_WDTH_L-1:0]        I401ab1ad994f5018061a3f57d3a51ad1;
wire [MAX_SUM_WDTH_L-1:0]        I3a47540f34ce47bcfa1da66cc4e6e088;
wire [MAX_SUM_WDTH_L-1:0]        I18916d0023ca275d84c52af07dcc5ca2;
wire [MAX_SUM_WDTH_L-1:0]        Ic79072d9e42dbc9974231f1d642b3f12;
wire [MAX_SUM_WDTH_L-1:0]        I1140fa91b5e22ba0c094c03295781e5a;
wire [MAX_SUM_WDTH_L-1:0]        Id2989aaee3930698cd374e6c9feedf82;
wire [MAX_SUM_WDTH_L-1:0]        Icda9a86a25dbe516a93b46fe487029e3;
wire [MAX_SUM_WDTH_L-1:0]        I53971b75cbd7ebc74b579776a6ea4778;
wire [MAX_SUM_WDTH_L-1:0]        I37e5c3118e8536e37bd797aeaa92476c;
wire [MAX_SUM_WDTH_L-1:0]        I9c68bfa3b888b6a6d41e38e674578284;
wire [MAX_SUM_WDTH_L-1:0]        I2c72d6c5fa6968dffa6517cf81219875;
wire [MAX_SUM_WDTH_L-1:0]        I9bb4d58b1fe80549451b00c4ed2b3885;
wire [MAX_SUM_WDTH_L-1:0]        Ic488e78b5c73251b673301e84c4b5b0b;
wire [MAX_SUM_WDTH_L-1:0]        I8d07beccef519ab4ce4024d911ac2346;
wire [MAX_SUM_WDTH_L-1:0]        I7c191c2c2be09886d0f31e4368797afd;
wire [MAX_SUM_WDTH_L-1:0]        Ia3bfd86e26efbef2cf6bb72be7ac1453;
wire [MAX_SUM_WDTH_L-1:0]        I4ae59dd2f57bda295e11b077e8668f1a;
wire [MAX_SUM_WDTH_L-1:0]        I3f6fad8bb0fba790fcdb1612b6fa7712;
wire [MAX_SUM_WDTH_L-1:0]        I58416287b268462d28f55c6c2705e613;
wire [MAX_SUM_WDTH_L-1:0]        I106d0e71b7378d110b0a624e5cbf0d6e;
wire [MAX_SUM_WDTH_L-1:0]        I59adad4fd84c1fc233dc58f70a12779d;
wire [MAX_SUM_WDTH_L-1:0]        I8e01532a1ab9534b8de0474549d41a2e;
wire [MAX_SUM_WDTH_L-1:0]        I80af3dcb716f3474a7257700aef89b81;
wire [MAX_SUM_WDTH_L-1:0]        I07d68462362d8453e83570cc793c55db;
wire [MAX_SUM_WDTH_L-1:0]        I9a2bba3f62de5f750dc8161a488dc331;
wire [MAX_SUM_WDTH_L-1:0]        I71da7e172b2b967040b6e6d02ef9949e;
wire [MAX_SUM_WDTH_L-1:0]        Ib97b2670a6cd88b2327f07f62d887900;
wire [MAX_SUM_WDTH_L-1:0]        Ib2963b82260024e1853d297798d88d3c;
wire [MAX_SUM_WDTH_L-1:0]        I0722ec4e9d400f8eaeacd060e42de79c;
wire [MAX_SUM_WDTH_L-1:0]        I1972375d51767f0cffa5395a354b3493;
wire [MAX_SUM_WDTH_L-1:0]        Ifb19d75cfa0051107b5fba57bfc002b5;
wire [MAX_SUM_WDTH_L-1:0]        I9d05dc0e39e85c23b62f343a8de12e64;
wire [MAX_SUM_WDTH_L-1:0]        I64ae3cd6f36b8bde29cd3e1fcba7bade;
wire [MAX_SUM_WDTH_L-1:0]        Ia6a78664c080829664158f53ba330312;
wire [MAX_SUM_WDTH_L-1:0]        I2ba16a10a82c20d54c776a9804ee50e4;
wire [MAX_SUM_WDTH_L-1:0]        Ie9a316de516ec4fb828a614c67e38b2a;
wire [MAX_SUM_WDTH_L-1:0]        Ie945349d77442536992d9ad52ce84218;
wire [MAX_SUM_WDTH_L-1:0]        Ic6a7a82d16e6106071934ba79d3698cd;
wire [MAX_SUM_WDTH_L-1:0]        Ide40b1bf9c0b642c49a5685a62af1c93;
wire [MAX_SUM_WDTH_L-1:0]        I79280400a4c9bed015106e5d006de757;
wire [MAX_SUM_WDTH_L-1:0]        Ic6e3847f035738243f4c5f71f296da57;
wire [MAX_SUM_WDTH_L-1:0]        I45b64b2b963963d2d0a8318133941f1d;
wire [MAX_SUM_WDTH_L-1:0]        I1939152ddbede923cde577984e0aa743;
wire [MAX_SUM_WDTH_L-1:0]        Ifbcebda2bb0ce58a0e1764c392a816df;
wire [MAX_SUM_WDTH_L-1:0]        I6d0d098e6d47dea04d6d7be67b648a0d;
wire [MAX_SUM_WDTH_L-1:0]        Icaeb9a2ec8ec5822658fa85b88cca04b;
wire [MAX_SUM_WDTH_L-1:0]        I3cc30aaba3dcd3eda262a19e85e53117;
wire [MAX_SUM_WDTH_L-1:0]        Ic0b2f9717b8aacb34325fd5aaf03a366;
wire [MAX_SUM_WDTH_L-1:0]        I002869e450d79649d27441ce00bfb575;
wire [MAX_SUM_WDTH_L-1:0]        Ie4d20df6b1e7a42f0df9a3cc26b12ac1;
wire [MAX_SUM_WDTH_L-1:0]        Idd01d014f0469f893305057ae3f4cb2e;
wire [MAX_SUM_WDTH_L-1:0]        I79444eef1875b6ad1a0675b66392ff9d;
wire [MAX_SUM_WDTH_L-1:0]        I7caf8c7496dd96c1ed08e98b415f5775;
wire [MAX_SUM_WDTH_L-1:0]        I7fc6e2aecff5bd691872d1e10a39103b;
wire [MAX_SUM_WDTH_L-1:0]        I49321308413cb4dbe5e6c01ba5b9023c;
wire [MAX_SUM_WDTH_L-1:0]        Id27560fb44b4f2fda98d47e9f20d6898;
wire [MAX_SUM_WDTH_L-1:0]        I745187336b8a5ae4eac66e90539752cf;
wire [MAX_SUM_WDTH_L-1:0]        I772e844c41387e7079259875e0ba3fa0;
wire [MAX_SUM_WDTH_L-1:0]        I32c35da92922c5b477f8aba837fa6d92;
wire [MAX_SUM_WDTH_L-1:0]        I3bc01b072987a0c980615abbc2251e5f;
wire [MAX_SUM_WDTH_L-1:0]        If08adda7d796da7c7849e472a73282a3;
wire [MAX_SUM_WDTH_L-1:0]        Ife3bb8945e14d8746c82b66886293997;
wire [MAX_SUM_WDTH_L-1:0]        I45ef0ac486fe043f57e8a46aa91461a3;
wire [MAX_SUM_WDTH_L-1:0]        Ic0ae1191869e636f9e4391efe93309ae;
wire [MAX_SUM_WDTH_L-1:0]        Id92d779518ae724b5fef5221372f8f26;
wire [MAX_SUM_WDTH_L-1:0]        Id0762ac7710c93249bc11c6ce4ae51a0;
wire [MAX_SUM_WDTH_L-1:0]        Ife6be241bc50560a14f97650e5cc2959;
wire [MAX_SUM_WDTH_L-1:0]        I1062442edb2bff727ca6283c8270bf28;
wire [MAX_SUM_WDTH_L-1:0]        I6c9ae8b8191507f908c27bbde53bf2d5;
wire [MAX_SUM_WDTH_L-1:0]        Iec936eeebd1f8c95307bd8705e6def81;
wire [MAX_SUM_WDTH_L-1:0]        I6332af145d560e3f22a4a88106749f98;
wire [MAX_SUM_WDTH_L-1:0]        I0c121fa3e9e6e0e2e8291a594d6b4ceb;
wire [MAX_SUM_WDTH_L-1:0]        Ic3c59a5167cb83fd76ec6236572b1f3d;
wire [MAX_SUM_WDTH_L-1:0]        I3e8e280553edaa5c8555ace81ecc10e0;
wire [MAX_SUM_WDTH_L-1:0]        I3e466d40a4447a23953d96d2e6d61d47;
wire [MAX_SUM_WDTH_L-1:0]        I76e4c55148effeba62a4837cd19c5e51;
wire [MAX_SUM_WDTH_L-1:0]        Ie335e68643fd2b0a53351f4bd45c3475;
wire [MAX_SUM_WDTH_L-1:0]        I89f75107ea95f207b9e664a1f4f0746a;
wire [MAX_SUM_WDTH_L-1:0]        Ic8f0049e1298b14b4e039075dc0d5f74;
wire [MAX_SUM_WDTH_L-1:0]        I382153cec6f7d6258574e7c532186473;
wire [MAX_SUM_WDTH_L-1:0]        I351dc309e916f282cc1e19303eee4112;
wire [MAX_SUM_WDTH_L-1:0]        I9de5e90485b3f22e9003dc8a7b22a79b;
wire [MAX_SUM_WDTH_L-1:0]        Idc4171a40dd2470e852af37a461013c7;
wire [MAX_SUM_WDTH_L-1:0]        Ifae488cb68d95ea517376319eb11f1bf;
wire [MAX_SUM_WDTH_L-1:0]        I9cab38b69794ab661e12750cf69c822c;
wire [MAX_SUM_WDTH_L-1:0]        I24180fba17c21bacefa8a4514e4b685c;
wire [MAX_SUM_WDTH_L-1:0]        I83bbe6fa947f9f909e1a6785ab31901f;
wire [MAX_SUM_WDTH_L-1:0]        I202c385beeccee309104b66f8f096b2c;
wire [MAX_SUM_WDTH_L-1:0]        Idc549661d6694035874a3366704801c7;
wire [MAX_SUM_WDTH_L-1:0]        I778fbaea65beeb6de599490daf3b7e3c;
wire [MAX_SUM_WDTH_L-1:0]        I4fd45670f88265e5d7aa6582f3ad3ff8;
wire [MAX_SUM_WDTH_L-1:0]        I2d636a246d815a4d12c478794860dd40;
wire [MAX_SUM_WDTH_L-1:0]        I3319313fe1d2b4ec2626711b187b4a5a;
wire [MAX_SUM_WDTH_L-1:0]        I586aaa5c55efd37996b01febd3bc60a4;
wire [MAX_SUM_WDTH_L-1:0]        I95ccc219b5f5038641b38dff6db0b222;
wire [MAX_SUM_WDTH_L-1:0]        I5001118df37d08bd19d322aca8ff3996;
wire [MAX_SUM_WDTH_L-1:0]        I22c15857572603cc24d8a87cb47c33b0;
wire [MAX_SUM_WDTH_L-1:0]        Ifdcd91f925b63e0817798aa6e9200e50;
wire [MAX_SUM_WDTH_L-1:0]        I8435e69bc1ff06e7edfabbee7b9aa49e;
wire [MAX_SUM_WDTH_L-1:0]        Ibeff607ba15fd8ef504224a9c1d102fc;
wire [MAX_SUM_WDTH_L-1:0]        Id15c3bdce785df234c68432ccec8f959;
wire [MAX_SUM_WDTH_L-1:0]        I25888aa2135fc403ca9eac4df634549a;
wire [MAX_SUM_WDTH_L-1:0]        I632ffd09a9091335b3aa91ab2a8f1cce;
wire [MAX_SUM_WDTH_L-1:0]        I283331db80e6d0891b13dc55e6a7d76c;
wire [MAX_SUM_WDTH_L-1:0]        I134a734d93e62f6ac6635015fe3a2096;
wire [MAX_SUM_WDTH_L-1:0]        Id66798f8ea67e74a67f264fe6b4503a3;
wire [MAX_SUM_WDTH_L-1:0]        If2ce7b8d2573494564393f7d426fa47f;
wire [MAX_SUM_WDTH_L-1:0]        Id59cf860d9f4aff11b205b8970d93df3;
wire [MAX_SUM_WDTH_L-1:0]        I75aaeab4f372e28a8e51453540f9c6b2;
wire [MAX_SUM_WDTH_L-1:0]        I2266afbacf1ba750ce18f296aba1181d;
wire [MAX_SUM_WDTH_L-1:0]        I69c2b063e61e14f5d49b907095ece00f;
wire [MAX_SUM_WDTH_L-1:0]        If077c67a062095cfe69f2260cee82833;
wire [MAX_SUM_WDTH_L-1:0]        Ibc03a9b6115d0941ce9233df7ef2fa57;
wire [MAX_SUM_WDTH_L-1:0]        Ia18bdb8d2f02b50281f0acd4a45ac973;
wire [MAX_SUM_WDTH_L-1:0]        Ib88c884e54d6e6ecf5ac015bc304e4f3;
wire [MAX_SUM_WDTH_L-1:0]        If6f5efee5e1f9709d86bf28cfb741955;
wire [MAX_SUM_WDTH_L-1:0]        Ia0caf6693d441ac622f416a86b665166;
wire [MAX_SUM_WDTH_L-1:0]        I85dd6a9634284c22027b4241551ea628;
wire [MAX_SUM_WDTH_L-1:0]        Id5cedaa397ebfc2567efcc2f8a648db5;
wire [MAX_SUM_WDTH_L-1:0]        Ica0a119af1728ae253c16cc3eb93f802;
wire [MAX_SUM_WDTH_L-1:0]        Ie7274a7ffa053ced4f12a67986d3c81b;
wire [MAX_SUM_WDTH_L-1:0]        Ife7985db888089ea618413810611bfca;
wire [MAX_SUM_WDTH_L-1:0]        If49068db99aa9d09302eda27ab51fcb7;
wire [MAX_SUM_WDTH_L-1:0]        I2959f2dc554e599d675eb6912757e413;
wire [MAX_SUM_WDTH_L-1:0]        I898d1b59aab3d5d4adce8ec3c0e14a0d;
wire [MAX_SUM_WDTH_L-1:0]        Ibb6e54edb9d277242c06d386a9a75a26;
wire [MAX_SUM_WDTH_L-1:0]        I51b1cd475d0e389326b182cbe680a402;
wire [MAX_SUM_WDTH_L-1:0]        If12366160fdc899bd71cb0de5bcfd84d;
wire [MAX_SUM_WDTH_L-1:0]        I44e5ce0cdf812c5b73e6e638da36e414;
wire [MAX_SUM_WDTH_L-1:0]        I4f38c3d620b72f21cf6d54c7df4ba816;
wire [MAX_SUM_WDTH_L-1:0]        Ib66b897398ea0702b74bdd03774f3ae4;
wire [MAX_SUM_WDTH_L-1:0]        I0b3a936c3f7e0391111e696b2445803b;
wire [MAX_SUM_WDTH_L-1:0]        I10f045edf47784a91a5599494c2d3de2;
wire [MAX_SUM_WDTH_L-1:0]        I6a81b4485598387e4656c35e83866209;
wire [MAX_SUM_WDTH_L-1:0]        Icf7630b6002db2f9b59d5323d6cc8105;
wire [MAX_SUM_WDTH_L-1:0]        I3db0adb3457cb22c755f5d29a8fe7ed8;
wire [MAX_SUM_WDTH_L-1:0]        I887911fd9466f4d4fa7f50642d610d88;
wire [MAX_SUM_WDTH_L-1:0]        I9ae284c0089ae462a1bb9d168bde2fd0;
wire [MAX_SUM_WDTH_L-1:0]        I342a563de39175fe4a6eb7e3e1ccac9a;
wire [MAX_SUM_WDTH_L-1:0]        Idc758f8e6fabb6b31b0a7d9c0c590310;
wire [MAX_SUM_WDTH_L-1:0]        I72b4ef48363856af7faacc85eafbaf2f;
wire [MAX_SUM_WDTH_L-1:0]        I4ae2f2330a8ee7d5626499f2a030c7a5;
wire [MAX_SUM_WDTH_L-1:0]        I4aa98503fc71292d42dba1cab6db952f;
wire [MAX_SUM_WDTH_L-1:0]        Ic35d5ac4dac46d47b2796bbac6452161;
wire [MAX_SUM_WDTH_L-1:0]        I32679702c19eab37b46d13bb372967ea;
wire [MAX_SUM_WDTH_L-1:0]        I6a86b03402bd2e35208d3fc74601f9cf;
wire [MAX_SUM_WDTH_L-1:0]        If8a259e0c4f1839e852abec6e1b904ee;
wire [MAX_SUM_WDTH_L-1:0]        I938dd59e4cdf3434086f60d000113430;
wire [MAX_SUM_WDTH_L-1:0]        Idc198bd5732ca5760d1a700a25273ce3;
wire [MAX_SUM_WDTH_L-1:0]        I9dfdffbfdb83572cc3205f674e5db753;
wire [MAX_SUM_WDTH_L-1:0]        I60520c850a95b893528569c4069bd677;
wire [MAX_SUM_WDTH_L-1:0]        If525ac3dc97e3187e036d70e9984939d;
wire [MAX_SUM_WDTH_L-1:0]        I0c1e4d400520935c5c78b792a9d554ba;
wire [MAX_SUM_WDTH_L-1:0]        Ic7d5fe6c4b1dcb97d10ba3de2f95d1df;
wire [MAX_SUM_WDTH_L-1:0]        I8efad9622c05177563ab8a2747879044;
wire [MAX_SUM_WDTH_L-1:0]        Ied4ddedaf801fbd7238d8a55c17c8090;
wire [MAX_SUM_WDTH_L-1:0]        Ieb9720b6beb2363d651346ef0233cd49;
wire [MAX_SUM_WDTH_L-1:0]        I202aa0814e7e28a6bd21db116b652b4d;
wire [MAX_SUM_WDTH_L-1:0]        Id201f81bbd80a70006a10866b8efeeff;
wire [MAX_SUM_WDTH_L-1:0]        Ic227f42a20219c6638ee3343ca445acf;
wire [MAX_SUM_WDTH_L-1:0]        I507e9bd0265d9ca6cd21a46fa21ba084;
wire [MAX_SUM_WDTH_L-1:0]        Ie04e44d8e0756cdf34cf9ad53da76e47;
wire [MAX_SUM_WDTH_L-1:0]        Ic92ab3dac1a151d6ff0b4e0c21003eb0;
wire [MAX_SUM_WDTH_L-1:0]        I3da241c7f221413abfbf1b4384bfca5a;
wire [MAX_SUM_WDTH_L-1:0]        I0807a826e91f92ef279ccf0b6512a428;
wire [MAX_SUM_WDTH_L-1:0]        I05aabdf73200996b7bea8db700fa8930;
wire [MAX_SUM_WDTH_L-1:0]        I03038b940be8bd21bd26b150b28754a6;
wire [MAX_SUM_WDTH_L-1:0]        Ibf547f8a5e1059ffaabeb3f447904dcf;
wire [MAX_SUM_WDTH_L-1:0]        I2ea27544ba4cc14d0f7ccf7158a27a2f;
wire [MAX_SUM_WDTH_L-1:0]        Ib2f34922b0d5346500de093275bebc94;
wire [MAX_SUM_WDTH_L-1:0]        Id2e223005a932987b6f60663773187f8;
wire [MAX_SUM_WDTH_L-1:0]        I3188d354c2ba494ffe210dcd89c00620;
wire [MAX_SUM_WDTH_L-1:0]        I09faa07bf38acd96c4e29afd8a5167e8;
wire [MAX_SUM_WDTH_L-1:0]        I6d4867d03d9187e95e27e99f7aecddec;
wire [MAX_SUM_WDTH_L-1:0]        Ifb09b84f9681c7bc28ffd562b633ffd9;
wire [MAX_SUM_WDTH_L-1:0]        Ib55b0e4c45ebbdb605f0ba9d62bff21c;
wire [MAX_SUM_WDTH_L-1:0]        I4319fa23d59f4e690e31fb7e3a823d17;
wire [MAX_SUM_WDTH_L-1:0]        I4ee3f608cc8f8df27345949f1a3713a7;
wire [MAX_SUM_WDTH_L-1:0]        Iede5d56e52612e083407888da49470e5;
wire [MAX_SUM_WDTH_L-1:0]        I3b2739319710681986b9d3f8cd04f619;
wire [MAX_SUM_WDTH_L-1:0]        I850c257a0412bd9bd6001817bd9d0ee1;
wire [MAX_SUM_WDTH_L-1:0]        Ib7875bf9d30d071e62a474c50d88ba06;
wire [MAX_SUM_WDTH_L-1:0]        Ia92b76ee5b7d82a992a1b58147c0c0be;
wire [MAX_SUM_WDTH_L-1:0]        I2253b32e46200a23dba243819fce02f0;
wire [MAX_SUM_WDTH_L-1:0]        I1b01cadaac7d3d15007f0afe5c0ab0f2;
wire [MAX_SUM_WDTH_L-1:0]        Ie96877deef8b1676138f814c4a720800;
wire [MAX_SUM_WDTH_L-1:0]        I8ce945d9f70bb317064a8d2d4eafd2d3;
wire [MAX_SUM_WDTH_L-1:0]        Iaed105b99eae5b078521e3a94d8a79b7;
wire [MAX_SUM_WDTH_L-1:0]        I05a812cd935867d1e417c64c26ea0952;
wire [MAX_SUM_WDTH_L-1:0]        Ic0a580f94f3d03f72e3a487f84bf6612;
wire [MAX_SUM_WDTH_L-1:0]        I39d9044227c161f0163e58dd82aadc90;
wire [MAX_SUM_WDTH_L-1:0]        I5f607bdc9b276fdf07a17a11a20a6720;
wire [MAX_SUM_WDTH_L-1:0]        I12e8b8cf609c2fbdc72efce9bb5dabee;
wire [MAX_SUM_WDTH_L-1:0]        I6fdccefd034e8b4b86cfa997502512ae;
wire [MAX_SUM_WDTH_L-1:0]        Idcd5283cf7b42d403ee0e4404b5b311b;
wire [MAX_SUM_WDTH_L-1:0]        Ia020344403aad35e050765a4b0cc42b7;
wire [MAX_SUM_WDTH_L-1:0]        Id11fd3a31b70da0e64138e71840cfb83;
wire [MAX_SUM_WDTH_L-1:0]        Ie9c5e7c98281cd1deb6acc51590c9d9a;
wire [MAX_SUM_WDTH_L-1:0]        Ia0e77e9544481aa0f56dfdb6eb253137;
wire [MAX_SUM_WDTH_L-1:0]        Iec0d7ea31e0f1a75b15121090dcf1e11;
wire [MAX_SUM_WDTH_L-1:0]        Ia98bb3648ce3719b1c31ce0f41121c63;
wire [MAX_SUM_WDTH_L-1:0]        Id9c8055ef530f2cb8096cb7bb2af55a4;
wire [MAX_SUM_WDTH_L-1:0]        Ib9081d438413a627f5b16f68c2eabb80;
wire [MAX_SUM_WDTH_L-1:0]        I9c5bf5451736358f8c84e150004fa5a9;
wire [MAX_SUM_WDTH_L-1:0]        I377933518c3807edb71f648c65ad5c85;
wire [MAX_SUM_WDTH_L-1:0]        Icec98d794a64752081fadfa74308fad3;
wire [MAX_SUM_WDTH_L-1:0]        I7bbe4d0a7d61d3f7da346de71b9a3a5f;
wire [MAX_SUM_WDTH_L-1:0]        I197c05f74bf7fb8d44124d40bd7c6563;
wire [MAX_SUM_WDTH_L-1:0]        I92acc55d81ec6e02880337b0a451ae21;
wire [MAX_SUM_WDTH_L-1:0]        I35c0ca76b28cd2f9355276b5d2f29ad4;
wire [MAX_SUM_WDTH_L-1:0]        I29da0e5661f29bd8493c19885c998582;
wire [MAX_SUM_WDTH_L-1:0]        I9426c8c1b4d988d5cd7d89a7aed4f8fc;
wire [MAX_SUM_WDTH_L-1:0]        Ibd010f15e36194cbd2ce9f01c98a2b6f;
wire [MAX_SUM_WDTH_L-1:0]        I7e86ab53e6d9647b230a94e076831ba2;
wire [MAX_SUM_WDTH_L-1:0]        Ia0ecfaedbc1d546d484978fd50096d10;
wire [MAX_SUM_WDTH_L-1:0]        I27098cbe2d4fdd634385d771cc290c2b;
wire [MAX_SUM_WDTH_L-1:0]        I5d7a0739e447775e00115799c52b11dd;
wire [MAX_SUM_WDTH_L-1:0]        Ie95793e09085b6de1383a37cc7fc41ac;
wire [MAX_SUM_WDTH_L-1:0]        Ib24b68cb35da39a743e1d90bba3f0836;
wire [MAX_SUM_WDTH_L-1:0]        Id4cdd72193e90dddd211af73d7f3634a;
wire [MAX_SUM_WDTH_L-1:0]        Iccab4c19a9190689f90a42160e2379de;
wire [MAX_SUM_WDTH_L-1:0]        I275ea08a3dc0600d8ccb6300eb7f2a6b;
wire [MAX_SUM_WDTH_L-1:0]        I1b53098a7240d2b5dc1f5c5c3b4bcc11;
wire [MAX_SUM_WDTH_L-1:0]        I278659ca1a0b093fc883d01987989dc0;
wire [MAX_SUM_WDTH_L-1:0]        If92e66cba66732798dd19f968a5ef8ce;
wire [MAX_SUM_WDTH_L-1:0]        I784c4e9fb75c314f271477e0621aaf7c;
wire [MAX_SUM_WDTH_L-1:0]        I3d3aafdd4d9d3e9fdab1f487c48a0ea9;
wire [MAX_SUM_WDTH_L-1:0]        Idb4c722992139f39914af7085378c6cc;
wire [MAX_SUM_WDTH_L-1:0]        I63c9deb7e6a4b400e0aff6887a09e647;
wire [MAX_SUM_WDTH_L-1:0]        Ie6f67c6e4c5e2b8357c0a902979e8722;
wire [MAX_SUM_WDTH_L-1:0]        I1d7a4f99e3975fd01bfe5a9a1da84765;
wire [MAX_SUM_WDTH_L-1:0]        I059d847e09f5aa3f6a8147062f4b13bf;
wire [MAX_SUM_WDTH_L-1:0]        I48e5256ade4d061a3b5ba08a53252bc3;
wire [MAX_SUM_WDTH_L-1:0]        I635fb29c55e0fb5cff0b6f443c2e3de5;
wire [MAX_SUM_WDTH_L-1:0]        I088c5b971a2def57248769a33b7d2a2d;
wire [MAX_SUM_WDTH_L-1:0]        Ide22394fce1658f9e7002bdb30d03c2f;
wire [MAX_SUM_WDTH_L-1:0]        I9ff276a14d3205b98174a8a736f79774;
wire [MAX_SUM_WDTH_L-1:0]        I123255637493b9c7924e3a72d1b86ee9;
wire [MAX_SUM_WDTH_L-1:0]        I87e6ef84894cfc86b94e19c9d3065bc6;
wire [MAX_SUM_WDTH_L-1:0]        I4c32900878260a261bc5403e8abd6258;
wire [MAX_SUM_WDTH_L-1:0]        Ifc100357ae3f754fb0e3863334bcc764;
wire [MAX_SUM_WDTH_L-1:0]        Iefe9e5376010997c0ee52eeb28e57a25;
wire [MAX_SUM_WDTH_L-1:0]        Ie6060acdcb16b6fa6aeeb649ed621053;
wire [MAX_SUM_WDTH_L-1:0]        I46c2b923860b0d1c01b9475f4467f280;
wire [MAX_SUM_WDTH_L-1:0]        I38b4eceb159ecb0dda3920290a21a02a;
wire [MAX_SUM_WDTH_L-1:0]        Ic45561ffe1837c3d5bb42c695a377f82;
wire [MAX_SUM_WDTH_L-1:0]        I3e76abc721bf7ed186f4d0f8f4bbf4e3;
wire [MAX_SUM_WDTH_L-1:0]        I1afb4061458e9d2f5799afa1f2373bd2;
wire [MAX_SUM_WDTH_L-1:0]        I18bb9a781a4c314fe6bd990e4c275f67;
wire [MAX_SUM_WDTH_L-1:0]        I49d7342f105c4502377abd23db973752;
wire [MAX_SUM_WDTH_L-1:0]        Ieeb12d463444ca36af1ecf2e09504c06;
wire [MAX_SUM_WDTH_L-1:0]        I17525df1798fa2c1c4bbc4a1ddcdd0a5;
wire [MAX_SUM_WDTH_L-1:0]        I90c44c31fa7903a81826c1c568597362;
wire [MAX_SUM_WDTH_L-1:0]        I3997cf122743b612f49cd5dd125a9201;
wire [MAX_SUM_WDTH_L-1:0]        I1112c4267582ddb8148ee40d9529beee;
wire [MAX_SUM_WDTH_L-1:0]        I21c207af859b94634d3750482b42a2ca;
wire [MAX_SUM_WDTH_L-1:0]        I2ff2421bd86bf9ec110724460f1171e9;
wire [MAX_SUM_WDTH_L-1:0]        I6ba5c453b17e4b33c61caf5d70041c4a;
wire [MAX_SUM_WDTH_L-1:0]        I08318099725fbe033ab8d5427eb8b278;
wire [MAX_SUM_WDTH_L-1:0]        If36cb462cdf20b0b1758cd6417e524fa;
wire [MAX_SUM_WDTH_L-1:0]        I40e8463645b1122b7cb224770fa00447;
wire [MAX_SUM_WDTH_L-1:0]        Ide386e751e06dd5df0c042cd76f0f800;
wire [MAX_SUM_WDTH_L-1:0]        If63bb4681bf1116c0d1db3aa21bf52ac;
wire [MAX_SUM_WDTH_L-1:0]        I566c72342c69969892480fae41232c37;
wire [MAX_SUM_WDTH_L-1:0]        Ia0f7deea6b1ce1050dcf97fa99de9178;
wire [MAX_SUM_WDTH_L-1:0]        I992b9876530d53c1b62d98511bf41942;
wire [MAX_SUM_WDTH_L-1:0]        Ib8861f627f6273c0a031bf43e7812a5d;
wire [MAX_SUM_WDTH_L-1:0]        Ieb5bac4ef0f5e4e0b826cdc43ae71471;
wire [MAX_SUM_WDTH_L-1:0]        I3cd0883d9f0ba7475f474f1e318ef023;
wire [MAX_SUM_WDTH_L-1:0]        I5f8a41ab83a9257e534973e981e28e9b;
wire [MAX_SUM_WDTH_L-1:0]        I0e420136675d5f0d1aa027d589ee8741;
wire [MAX_SUM_WDTH_L-1:0]        I4aab6ff52e3fba90bb7417cb50766125;
wire [MAX_SUM_WDTH_L-1:0]        I1ba7f209cb735471073e8051026a148c;
wire [MAX_SUM_WDTH_L-1:0]        I711c5cf9fd8c5161bac36060b3443503;
wire [MAX_SUM_WDTH_L-1:0]        Ie3591b22e0e127f04658da68d4846be9;
wire [MAX_SUM_WDTH_L-1:0]        I409129c0bf5d361e9916b6dc98e69a7d;
wire [MAX_SUM_WDTH_L-1:0]        Ie4f4faa470f572da2081b63b6df6e392;
wire [MAX_SUM_WDTH_L-1:0]        I5011dfbbb0eccfebcff255e4a2c5e64c;
wire [MAX_SUM_WDTH_L-1:0]        Ie32ca6b91d1c55883be8f63acca78764;
wire [MAX_SUM_WDTH_L-1:0]        I6c7965d39dc839a9df56e628c77a5457;
wire [MAX_SUM_WDTH_L-1:0]        Ieac9cea5f36bd82f87105b530e8fb614;
wire [MAX_SUM_WDTH_L-1:0]        I79657595561eac53237215fb4110f09d;
wire [MAX_SUM_WDTH_L-1:0]        I9b46463a6c54c3668e76190d942b7b38;
wire [MAX_SUM_WDTH_L-1:0]        I3ff883ad434cd5153b67186b6b21418d;
wire [MAX_SUM_WDTH_L-1:0]        I92abaae6fb89206885616877cca1e25a;
wire [MAX_SUM_WDTH_L-1:0]        I33668b0ef7defef974b7a4c0f87689c0;
wire [MAX_SUM_WDTH_L-1:0]        I338daeacf82ad288b14c6b5bd4099870;
wire [MAX_SUM_WDTH_L-1:0]        Ibe085a39ecb07a8dca62002afa38df93;
wire [MAX_SUM_WDTH_L-1:0]        I1f88dddf05f255942e2749891a7733da;
wire [MAX_SUM_WDTH_L-1:0]        If1d0be4e9b995ec98c346e8392b9518a;
wire [MAX_SUM_WDTH_L-1:0]        I56a4443759b3d786bc9a34a0dc32abf0;
wire [MAX_SUM_WDTH_L-1:0]        Ic826d371f2cfc503f5d9e43dc17481e1;
wire [MAX_SUM_WDTH_L-1:0]        I5502f383dff392ef1be4cbbf9dbc3c2f;
wire [MAX_SUM_WDTH_L-1:0]        I96e6f1dc0cd451da6ac9170d5f83976d;
wire [MAX_SUM_WDTH_L-1:0]        I10cd840a369d3e25556a41beede2be27;
wire [MAX_SUM_WDTH_L-1:0]        Id85c2285fcc45211f0fa6963b74a663a;
wire [MAX_SUM_WDTH_L-1:0]        Ie0bdfac78159144aa65090028931a3bf;
wire [MAX_SUM_WDTH_L-1:0]        I28fa30cd1f3b476fa6a354863108cbcf;
wire [MAX_SUM_WDTH_L-1:0]        I7a927f4f266cc5253ec30f5c127bb17a;
wire [MAX_SUM_WDTH_L-1:0]        I7571c7c306861230de71a75fca79c5dc;
wire [MAX_SUM_WDTH_L-1:0]        Ic79811a48840357d0b6303e7b19413dc;
wire [MAX_SUM_WDTH_L-1:0]        I0f29300446f020dd23cf847d3e3d3530;
wire [MAX_SUM_WDTH_L-1:0]        I802bd5b13c183c37e842f7e9278f35a9;
wire [MAX_SUM_WDTH_L-1:0]        I0297905b35f06697625420b7fc2434f7;
wire [MAX_SUM_WDTH_L-1:0]        I8487a819dcb61016798cde56f9662fcf;
wire [MAX_SUM_WDTH_L-1:0]        Ia2904a5d5db43a209bd4b358ace68c6a;
wire [MAX_SUM_WDTH_L-1:0]        Ia8b29ca047a643f47bd3a0ffb50bf8cb;
wire [MAX_SUM_WDTH_L-1:0]        Ic45d0537b94bc30713c0a0ee07b1ec40;
wire [MAX_SUM_WDTH_L-1:0]        I337231f0dc7eb85f7d950262e0adb724;
wire [MAX_SUM_WDTH_L-1:0]        I530cf1f747d1df44b913f49eee90c079;
wire [MAX_SUM_WDTH_L-1:0]        Ief52461e4a5ddb128be5e439edf34862;
wire [MAX_SUM_WDTH_L-1:0]        I46d86bfa6de26f3cfef9d802549ef2ad;
wire [MAX_SUM_WDTH_L-1:0]        If6a3bd6f002d91e0773c4ab9caaaa01e;
wire [MAX_SUM_WDTH_L-1:0]        Ib33e1c6d57e5e6fc465dc9c9a7cf29fa;
wire [MAX_SUM_WDTH_L-1:0]        Id92a319da408be46970faf524513fdd8;
wire [MAX_SUM_WDTH_L-1:0]        Iae182ffae6cea89363f0ccc8b5679561;
wire [MAX_SUM_WDTH_L-1:0]        Idfe6aecb694385ce8c3c1544a4992a20;
wire [MAX_SUM_WDTH_L-1:0]        Idfbc5726963cfa31bb4324143ffd08c7;
wire [MAX_SUM_WDTH_L-1:0]        I205d5fdeae55fae7be2f06f11c949244;
wire [MAX_SUM_WDTH_L-1:0]        Ie667e1755ae1561a2eefae9b63845dec;
wire [MAX_SUM_WDTH_L-1:0]        If7348fdbe0400aab92e8fd6a7cf6c267;
wire [MAX_SUM_WDTH_L-1:0]        I143b91852fddcdcc30bf1041332c4ed7;
wire [MAX_SUM_WDTH_L-1:0]        Iee5e74945ba15220f0f707c9c1927ba1;
wire [MAX_SUM_WDTH_L-1:0]        I4d1c47569b0bc8c651c897ac8e88bd1f;
wire [MAX_SUM_WDTH_L-1:0]        Ib9d6c5be487a434fbafcda25ca9351dc;
wire [MAX_SUM_WDTH_L-1:0]        Ib0d033ba28e8c606ed92207049c76884;
wire [MAX_SUM_WDTH_L-1:0]        I300d9f403e33d860ff5dde9f91bae11b;
wire [MAX_SUM_WDTH_L-1:0]        Iebfe0fa45e4b34e142e82ddaa15243cf;
wire [MAX_SUM_WDTH_L-1:0]        Ieb778442bc855e93e11c9b13f1a7ae06;
wire [MAX_SUM_WDTH_L-1:0]        I57a393cc9cc9e1abc7962aa2cc840a7c;
wire [MAX_SUM_WDTH_L-1:0]        I0ffb8b65525af38861280645ac310e3d;
wire [MAX_SUM_WDTH_L-1:0]        I30fb41a57460a0b1f21065b4b97ddd42;
wire [MAX_SUM_WDTH_L-1:0]        Ie8298c5c8ff538a3e37af46798f6d753;
wire [MAX_SUM_WDTH_L-1:0]        Ie7dc322fee8ca0b6b9659e5183e0d6d6;
wire [MAX_SUM_WDTH_L-1:0]        I91bbec0523f77fc52a88ebcc49267e9c;
wire [MAX_SUM_WDTH_L-1:0]        I38ae79956762380fadc94f8126dc1c90;
wire [MAX_SUM_WDTH_L-1:0]        Id55a1ab9d158ea509e5f57286a3d1b67;
wire [MAX_SUM_WDTH_L-1:0]        Ice615e7e18356ae4c3f615dd997be943;
wire [MAX_SUM_WDTH_L-1:0]        I57b40c72004f2c3072cbdefbeef72b7c;
wire [MAX_SUM_WDTH_L-1:0]        Ie38351e19bdc4f2ce9caf75fc3937dd4;
wire [MAX_SUM_WDTH_L-1:0]        Ibba6269b560db9d4913e1e515ed8270d;
wire [MAX_SUM_WDTH_L-1:0]        Ie392719059587a201c0148138ba2a2d4;
wire [MAX_SUM_WDTH_L-1:0]        I4852d6bacfd82fef6fab4502d61e9a37;
wire [MAX_SUM_WDTH_L-1:0]        I9200526d94c38e638370e9a2d7fed75c;
wire [MAX_SUM_WDTH_L-1:0]        I15b8aa7d973edcf3b2365040f5570d82;
wire [MAX_SUM_WDTH_L-1:0]        Ic3f8e77259ee3eb5be80e11b607818bd;
wire [MAX_SUM_WDTH_L-1:0]        Iabf228f57ac154c417389f6711af1950;
wire [MAX_SUM_WDTH_L-1:0]        If37de611ce4fa330c4fc9dcb87d4d95c;
wire [MAX_SUM_WDTH_L-1:0]        If3c44eb85217da3b6bddb5aed97a9bb7;
wire [MAX_SUM_WDTH_L-1:0]        I8c36318c45dabe6bf540381373f09fe5;

wire [flogtanh_WDTH -1:0]        Ia67805b59c3011bc4fc5cb1d2996f90d;
wire [flogtanh_WDTH -1:0]        I5f68368511b59d2e365cc91b806b334e;
wire [flogtanh_WDTH -1:0]        I61fb47b07547e09c746b1fb5d7c8710d;
wire [flogtanh_WDTH -1:0]        I71e4d98dca37256fcc84248a26d703e2;
wire [flogtanh_WDTH -1:0]        Ib2220549c84e87683ccf85798b2bb22f;
wire [flogtanh_WDTH -1:0]        Ib8380902ac4082f834744ddef6d0cc6a;
wire [flogtanh_WDTH -1:0]        I12f063ad18938c2ca008e1165f9119e9;
wire [flogtanh_WDTH -1:0]        I9570f8498d95bee230bb3c5e720bb857;
wire [flogtanh_WDTH -1:0]        Iae6b4023f9f2641ca00636181f4fb028;
wire [flogtanh_WDTH -1:0]        I55c425102db0a6838012a165c0597680;
wire [flogtanh_WDTH -1:0]        Id11b7d1aeb413fd4920ef0e0097fc6c4;
wire [flogtanh_WDTH -1:0]        Ic970a88c435a85d21ed71c6060b8a8e4;
wire [flogtanh_WDTH -1:0]        I3af03d3e0bb7e0e73e034dceda70ff3a;
wire [flogtanh_WDTH -1:0]        Iec8dc328edd6cbaa2d697e05ed222746;
wire [flogtanh_WDTH -1:0]        Iba30a494dc1b66bd2862f82c16017a99;
wire [flogtanh_WDTH -1:0]        I16d2084ccfb102c3bafc701872f5ef2d;
wire [flogtanh_WDTH -1:0]        Iefa075dc743d616eca65f76d2c03371c;
wire [flogtanh_WDTH -1:0]        Id680a9affed622577164b3a8380494f5;
wire [flogtanh_WDTH -1:0]        Icc7a632da404a9cda7b8247706391f85;
wire [flogtanh_WDTH -1:0]        Ifcd68be4bea38622d2d57d3a4e6fc5bb;
wire [flogtanh_WDTH -1:0]        I708c5d8d6d8f7f16c2f348c3b97b906d;
wire [flogtanh_WDTH -1:0]        I16deb9107193a3536979e4b5e5654b9c;
wire [flogtanh_WDTH -1:0]        I51ba1e25e01c39a77559089626bafa09;
wire [flogtanh_WDTH -1:0]        I28cac65a4db3f708cc90a1b023bfe894;
wire [flogtanh_WDTH -1:0]        I2217e483aaf5124d9beb9baf5037326b;
wire [flogtanh_WDTH -1:0]        Ie763738b7faf253837e1c45de255cb5e;
wire [flogtanh_WDTH -1:0]        Ib47f8220e7a319e690649f9d6cc9f0cc;
wire [flogtanh_WDTH -1:0]        Icfef12499b53cd84f0aae067f30c17d0;
wire [flogtanh_WDTH -1:0]        Iffc502b536d88d080c59eb3aedd55bd1;
wire [flogtanh_WDTH -1:0]        I0982b8d7f99aceb8871c9c10448f54c5;
wire [flogtanh_WDTH -1:0]        Iaa823b6b13acb376f979dd52683a2231;
wire [flogtanh_WDTH -1:0]        I6c661048307c23c699d4b3636564de0f;
wire [flogtanh_WDTH -1:0]        Ic5f3f371b1ebfe733404b4165fe746dc;
wire [flogtanh_WDTH -1:0]        I786dfcaa131b99c254aaff15bd2c2b6d;
wire [flogtanh_WDTH -1:0]        I021d991730d154218106f00e74bf9d4c;
wire [flogtanh_WDTH -1:0]        I2b49d74cb130542f2ca99534e2c513b1;
wire [flogtanh_WDTH -1:0]        I688e5b6520508178afdf85bb2194186d;
wire [flogtanh_WDTH -1:0]        I0f6cb7a5a31d6f2f6178632c0c898bc6;
wire [flogtanh_WDTH -1:0]        I658630f3cf0e86ea86c5fb78b025b0a5;
wire [flogtanh_WDTH -1:0]        I03bea609a189246a2375b355df47cf81;
wire [flogtanh_WDTH -1:0]        I8b17f8bae259d829b52aba173bf10b4f;
wire [flogtanh_WDTH -1:0]        If56555b7cf539750706cf678030ccdb2;
wire [flogtanh_WDTH -1:0]        I944da8181119550916eaf431c7b04c50;
wire [flogtanh_WDTH -1:0]        I94e89b3a841f9760e3967c97e86d7160;
wire [flogtanh_WDTH -1:0]        I3aa615fa11ad382432ca658ec233f094;
wire [flogtanh_WDTH -1:0]        I8cab6f6faf0758f26d1a8851fae43896;
wire [flogtanh_WDTH -1:0]        Ib7c4f77c160ec436e93ca9de75b9fe42;
wire [flogtanh_WDTH -1:0]        I6ecf7249e6151477fe74a79d0b126b21;
wire [flogtanh_WDTH -1:0]        Ic1e06942b276ee0933dc8b85dec58756;
wire [flogtanh_WDTH -1:0]        I3753b2c4ba8f1bee70def390a96586b0;
wire [flogtanh_WDTH -1:0]        Idd96d8b4e7be386203ec3ed3a81391d9;
wire [flogtanh_WDTH -1:0]        I9b919f3d4ee3f33506b87bcdaf2d43a3;
wire [flogtanh_WDTH -1:0]        I7df43eec4d78baa1e0680be2715c4495;
wire [flogtanh_WDTH -1:0]        Ib3be128b6704cc04c61e0fc9814dcf20;
wire [flogtanh_WDTH -1:0]        Ief08536c38479e6bc7fe786cfaf9a10f;
wire [flogtanh_WDTH -1:0]        If365a3c3ef86dca7c7315b91298c2db8;
wire [flogtanh_WDTH -1:0]        I6ef440b2077563ebbe50dde593c3875a;
wire [flogtanh_WDTH -1:0]        I83560e8d0f8cd37815cca6336fb2208d;
wire [flogtanh_WDTH -1:0]        I20cfad172f0a614687d72d2337ef1003;
wire [flogtanh_WDTH -1:0]        I099441ae3d3dffe49b18bc578af54dc7;
wire [flogtanh_WDTH -1:0]        Icc6a92285959b25d53b452aed0718c8e;
wire [flogtanh_WDTH -1:0]        I58f89947eead94b5054a0fea3520ae33;
wire [flogtanh_WDTH -1:0]        I132c12f1eafbe34bca7b070354bd5f43;
wire [flogtanh_WDTH -1:0]        Ibf565bf1803ed43120fa54b80f6f1f29;
wire [flogtanh_WDTH -1:0]        I0f327225758bc82a67a65b8714949a91;
wire [flogtanh_WDTH -1:0]        I619957528c630e7f64924a25127c93fb;
wire [flogtanh_WDTH -1:0]        Ia90d4bc44d3687e912b59e4b6ca02718;
wire [flogtanh_WDTH -1:0]        If3cc31fd16469339470702045fc6d0da;
wire [flogtanh_WDTH -1:0]        I21c1757545cc2732445c7f978f7247c4;
wire [flogtanh_WDTH -1:0]        I338ccc17dc6158aec0129c8b0c02c429;
wire [flogtanh_WDTH -1:0]        I096fb1aff9431ed667e5d85a6f3726a4;
wire [flogtanh_WDTH -1:0]        I83d71a89f35eb73265ee3e54184e1277;
wire [flogtanh_WDTH -1:0]        Ia69d80cc1f2957ccd79cbd466dea987e;
wire [flogtanh_WDTH -1:0]        I7362f08ed4e4ae309dfbfda112c56ad6;
wire [flogtanh_WDTH -1:0]        I2243822bb5cdbca7f2ea942c7b720da8;
wire [flogtanh_WDTH -1:0]        I8be4be8471625db0749e6385f87d2dcc;
wire [flogtanh_WDTH -1:0]        Ia77953e90a0cb40984d138c2c209db01;
wire [flogtanh_WDTH -1:0]        I3d6a685a1913bd8be01fddbce1edec2e;
wire [flogtanh_WDTH -1:0]        Id0b03e6dafabbe570f2626f51c9b7121;
wire [flogtanh_WDTH -1:0]        Ifd77e040c5f82790b1d5636a42fca602;
wire [flogtanh_WDTH -1:0]        I5bfac7858439b218179c95c8d8669f17;
wire [flogtanh_WDTH -1:0]        Ifbe479e5cab3cba43444bec1e12e72a0;
wire [flogtanh_WDTH -1:0]        I52497c500164c2417f928196ddcdbf84;
wire [flogtanh_WDTH -1:0]        Ia784f35a5a46837b69eb048dabf84052;
wire [flogtanh_WDTH -1:0]        Ib499dd504da7e433bc1caa258d7e7101;
wire [flogtanh_WDTH -1:0]        I8d0f440df332ea96e2d56eec490fbd51;
wire [flogtanh_WDTH -1:0]        I7af88e2be096e488d7269479f935d185;
wire [flogtanh_WDTH -1:0]        I8d431a0524241fa54cf6dd1e79de4c74;
wire [flogtanh_WDTH -1:0]        Ief51cc849e0034a9a6b3ff061064ad64;
wire [flogtanh_WDTH -1:0]        If49f97cc0c42b23ce393b534015559a0;
wire [flogtanh_WDTH -1:0]        Ic5f096a42ae6fec933dcaf85faeeda49;
wire [flogtanh_WDTH -1:0]        Ie932a22a7f1fa37087cbc9e8d73efef4;
wire [flogtanh_WDTH -1:0]        Ic9c0a2ce51d641ba7896c2c6911d0f96;
wire [flogtanh_WDTH -1:0]        I2956687a5fc2fba7149889624ef85647;
wire [flogtanh_WDTH -1:0]        Ia96b3ea2e8395671b3ac674f5a956771;
wire [flogtanh_WDTH -1:0]        Iebf28886bd39c2540c90e808a9c20d3d;
wire [flogtanh_WDTH -1:0]        Ib81d241e073c97c8c8d1d0abd9a9a64f;
wire [flogtanh_WDTH -1:0]        I8d4f3e64c8e3b0710a4a6b30d27c8be8;
wire [flogtanh_WDTH -1:0]        I0fc5e49719d7132c7724ee0d406ff93e;
wire [flogtanh_WDTH -1:0]        I16e3f3a6802fd206654bb622fa1393fe;
wire [flogtanh_WDTH -1:0]        I4479a0c26d4fa67dee328ecae12d14a4;
wire [flogtanh_WDTH -1:0]        I4b5713aee09999592256c407d4b8a95a;
wire [flogtanh_WDTH -1:0]        If5693e079544d04478ec3da9a0ba28d7;
wire [flogtanh_WDTH -1:0]        Ieb1dbb98d5e5bda5b9ce803857f2ca26;
wire [flogtanh_WDTH -1:0]        I701a0ec899c88feef97aeb45fe19e639;
wire [flogtanh_WDTH -1:0]        Ife1c8d014675240a94f1133a78703ed5;
wire [flogtanh_WDTH -1:0]        I6e9d61b111a45e4ea92ff12d33801755;
wire [flogtanh_WDTH -1:0]        I94d9412a7b43fa0bd4b9a6d32d313fc7;
wire [flogtanh_WDTH -1:0]        Ief65b0dab6ce1c2fc23cd297a21ac8de;
wire [flogtanh_WDTH -1:0]        If13e359e530823319046ce20027445dd;
wire [flogtanh_WDTH -1:0]        Ibb843c4198a06c8e46bc954663c52a28;
wire [flogtanh_WDTH -1:0]        I221777352b48c4e228c6637410113854;
wire [flogtanh_WDTH -1:0]        I0c043ef5daa388e93fb3cf6465c217b5;
wire [flogtanh_WDTH -1:0]        I1ee46fec2b82cf8e5142f8e2ac5d9d8a;
wire [flogtanh_WDTH -1:0]        Ife3f07ad3ad5228f10da7020a01e7069;
wire [flogtanh_WDTH -1:0]        Ie45aaf966aa0a94803050b5f43d69e6c;
wire [flogtanh_WDTH -1:0]        I2dacd37cecd93c6e9134cb55ed917d78;
wire [flogtanh_WDTH -1:0]        I88aedd7f52399f5fd435c3415f2218ca;
wire [flogtanh_WDTH -1:0]        I2419bc316181acd41e29ad005241d812;
wire [flogtanh_WDTH -1:0]        I7651176b0a74846108fbaabc5cc4900a;
wire [flogtanh_WDTH -1:0]        I35faf0af91f4972ae843883993fc84f4;
wire [flogtanh_WDTH -1:0]        I57ac487adc18165136e9b3c7c50f95ad;
wire [flogtanh_WDTH -1:0]        I4dd2e7b6a685958d7aac77a38354e05f;
wire [flogtanh_WDTH -1:0]        Ic95668328a2121027436f682bac50b9c;
wire [flogtanh_WDTH -1:0]        Ib27460a2e2b13abc54f5ba37f32c8653;
wire [flogtanh_WDTH -1:0]        I118726375ca9381e45f001965fcefc5b;
wire [flogtanh_WDTH -1:0]        Ia3fa91387788798672eb6199a2eaa389;
wire [flogtanh_WDTH -1:0]        Ic8d47ff5d6c31601a57df868da78c2d4;
wire [flogtanh_WDTH -1:0]        Ieecd194ccc5698a2ba16efd969cfd621;
wire [flogtanh_WDTH -1:0]        I7cdc5ada6fc68ee31fd4062e2ff004d3;
wire [flogtanh_WDTH -1:0]        Ifb09fa1840c5a1ddbfc81cda21c11f1e;
wire [flogtanh_WDTH -1:0]        I59547aacdcfde31dc016ec2acbb2f4b4;
wire [flogtanh_WDTH -1:0]        I4ce505ae2025bab3abcf5a44e0ed5034;
wire [flogtanh_WDTH -1:0]        Ia7f53f0cd86055da72c13ac474f052a1;
wire [flogtanh_WDTH -1:0]        Id40a7ca1cde7a70cc13e752e19132808;
wire [flogtanh_WDTH -1:0]        I915054f2fbb8b93516d8748a3e3e29e2;
wire [flogtanh_WDTH -1:0]        If7274be2bcc8b2a235c3538db5506d90;
wire [flogtanh_WDTH -1:0]        If257757fa31c2f4cc9ec322e4ecccf83;
wire [flogtanh_WDTH -1:0]        I3e611982ec9ff6437f22e11b2552693a;
wire [flogtanh_WDTH -1:0]        If91268e2b84df18785cd6a53e53eb4e9;
wire [flogtanh_WDTH -1:0]        I8fcf0a468234f365c33059e26b9f5821;
wire [flogtanh_WDTH -1:0]        Ia072f1d679429d3c3180f8eb67fc7dd7;
wire [flogtanh_WDTH -1:0]        I3f80250ee19e8250898f2bcc055c2e5b;
wire [flogtanh_WDTH -1:0]        I91a8168d3b087ab3891cd6d479427b95;
wire [flogtanh_WDTH -1:0]        I06b3652935db14aaa057f0cf3cffef66;
wire [flogtanh_WDTH -1:0]        Id1dce8c1542f1279badb381aca3c9b51;
wire [flogtanh_WDTH -1:0]        Ib01d30e88a3a1fcb204246baafeb47c8;
wire [flogtanh_WDTH -1:0]        I8983f003c30a218543f39f5bbcd9a25c;
wire [flogtanh_WDTH -1:0]        I9f688c58878405d1d2865ddc40659c2b;
wire [flogtanh_WDTH -1:0]        Id1b5c33bc63f75561b7cce6fc0981c69;
wire [flogtanh_WDTH -1:0]        Ic9c77123914f831cee5bc4586b6a2a8b;
wire [flogtanh_WDTH -1:0]        I003f95fb8f2027efa41a1936e8b53986;
wire [flogtanh_WDTH -1:0]        Ifd42760504e0f106eb9061d9b9a2d18a;
wire [flogtanh_WDTH -1:0]        Ie16dc913f571ae73ce03d755077345a9;
wire [flogtanh_WDTH -1:0]        I452794105cca79653f5509dac3794327;
wire [flogtanh_WDTH -1:0]        I86e53eed5b857c439039238bb486067c;
wire [flogtanh_WDTH -1:0]        I33431ed9c549f5525adfa5d45fbc7653;
wire [flogtanh_WDTH -1:0]        I89433799cfa534afd66e8d6b9f1b62b9;
wire [flogtanh_WDTH -1:0]        I4b8b4fd334b176cb449ad0296ebff4c8;
wire [flogtanh_WDTH -1:0]        I80f2e8f6743e28e86e4d85b295e2f768;
wire [flogtanh_WDTH -1:0]        I66e7dacba9dbfb14e9a71b9d57229880;
wire [flogtanh_WDTH -1:0]        I1391018fb93372ccc2fcc08700e38b65;
wire [flogtanh_WDTH -1:0]        If3a842c52c8c0b2fd24ef265e8cfe330;
wire [flogtanh_WDTH -1:0]        I8fd26d47ecd4cdd08294cf6133468d17;
wire [flogtanh_WDTH -1:0]        I0f3aea4265966e7bc673d3a08ad1c2e4;
wire [flogtanh_WDTH -1:0]        I7097c9518bb3351818b96f31ed49c6d3;
wire [flogtanh_WDTH -1:0]        Ia9de78211d220e68835ff757eb75d919;
wire [flogtanh_WDTH -1:0]        Id683d693cd50645c3d6d657aa1c8bdb2;
wire [flogtanh_WDTH -1:0]        I2c1c31b8bda73b145cdf74b18bc46a4d;
wire [flogtanh_WDTH -1:0]        I88bd8012c93dd9e2ed52ea5e9b8b0004;
wire [flogtanh_WDTH -1:0]        I300a84deada851e18835d6af55c5e2a3;
wire [flogtanh_WDTH -1:0]        Ia8d3667adc34b2b50acf7edb970538d8;
wire [flogtanh_WDTH -1:0]        I1fc6745ba86be641dc9bdac044c19519;
wire [flogtanh_WDTH -1:0]        I3f0bba472e912f11dea8e788fbc1cb63;
wire [flogtanh_WDTH -1:0]        I2791cc5f69dd0e7f306760048c759af7;
wire [flogtanh_WDTH -1:0]        I6dc671e73b4e9c70cabfdeaac2e5c40b;
wire [flogtanh_WDTH -1:0]        Ie8157cde860052619820431f87e13c83;
wire [flogtanh_WDTH -1:0]        Ia6255a136d5f36ea6cba654bd5823850;
wire [flogtanh_WDTH -1:0]        I9059b74a8f3cf2e4905756cc9c71597f;
wire [flogtanh_WDTH -1:0]        I2b9584392ef9a7828ff57bd4c522a302;
wire [flogtanh_WDTH -1:0]        I99584eabd3cbd2546c85f474afa6fabb;
wire [flogtanh_WDTH -1:0]        I6c1235e88ae444a96ea64fd1bfd04d8f;
wire [flogtanh_WDTH -1:0]        I047abade6abf10a65a5b835ac725fa7c;
wire [flogtanh_WDTH -1:0]        Id09b8242c22851fb960d55222fe733d4;
wire [flogtanh_WDTH -1:0]        Icf7ab1d1113bc44358c56a56fca7caf9;
wire [flogtanh_WDTH -1:0]        Ie355fa27abbc41291eaf08f2cf9a6ff7;
wire [flogtanh_WDTH -1:0]        I4d24650be7a1088c2310d93000d6392a;
wire [flogtanh_WDTH -1:0]        I566224393f6bb27bfd8b0b0d6b8e53d6;
wire [flogtanh_WDTH -1:0]        Ic3aea8ebb8eab44a92e7d7d950e1a917;
wire [flogtanh_WDTH -1:0]        I8fcad6e7d5ffc9f79eaaf634f6fe8cda;
wire [flogtanh_WDTH -1:0]        I82af0956870500474eac2505bbf15e35;
wire [flogtanh_WDTH -1:0]        I6f0f74dcc830fdcb0af9df75a2b722f7;
wire [flogtanh_WDTH -1:0]        I2d8a8efaa0179340bf5d3ebbd4c11831;
wire [flogtanh_WDTH -1:0]        Idd95fd099dd2b53c46d02f09575b8032;
wire [flogtanh_WDTH -1:0]        I32ff895ff659ec448270067f76e97a90;
wire [flogtanh_WDTH -1:0]        I0f277bc88d46a4e6e9f1f2c410b503fd;
wire [flogtanh_WDTH -1:0]        I15a7fd79aeb5eed24b1c7be3d48296e0;
wire [flogtanh_WDTH -1:0]        I66b92f1de2cf408c3af53b161a6ffa60;
wire [flogtanh_WDTH -1:0]        I12f311f2311e26320a178d6fec95d9d0;
wire [flogtanh_WDTH -1:0]        Id28d9545e8d20ac080fbac5e345692da;
wire [flogtanh_WDTH -1:0]        I2b8ce30d1338ad506e4996d2dd1dc11a;
wire [flogtanh_WDTH -1:0]        I4a5cfd6ebd47cda4fa2e06ba9ad6e5b2;
wire [flogtanh_WDTH -1:0]        Ic2b65e7bd42e94f2ad8b6506a6fce7af;
wire [flogtanh_WDTH -1:0]        I62bda8dc70e0b5eb38abe094bbe92fc6;
wire [flogtanh_WDTH -1:0]        I0f54a697ea3e2bbf90354c9a6173fb80;
wire [flogtanh_WDTH -1:0]        I223b05d94c09b095d1988df121aa5e37;
wire [flogtanh_WDTH -1:0]        I6a6c0f8e4399c21285d66ddc0f1f70c0;
wire [flogtanh_WDTH -1:0]        I5f73e5faf1aca83ee0a415c9ac4a1b9a;
wire [flogtanh_WDTH -1:0]        Ibfcdfc01f09bcff031e359394947efef;
wire [flogtanh_WDTH -1:0]        I75f9d3a41019dca3044a1c2cf7069662;
wire [flogtanh_WDTH -1:0]        I8efd478f1ae2ea6090774e1ed3bd7b28;
wire [flogtanh_WDTH -1:0]        I820fa56328e3919970dd64adb1d4d8e7;
wire [flogtanh_WDTH -1:0]        I502d3210c60c82ca682d8e2168d54be0;
wire [flogtanh_WDTH -1:0]        I05eadf11cdc6c2f2b021e33f2438fa49;
wire [flogtanh_WDTH -1:0]        I337d74c3c773a358a936806f751c1117;
wire [flogtanh_WDTH -1:0]        I2c487770d606451440eecf358202db32;
wire [flogtanh_WDTH -1:0]        Ia494fdbd70bff11510eb685f3b5d0aae;
wire [flogtanh_WDTH -1:0]        I082aa8c413d7ef8f054b1c2857cbe39f;
wire [flogtanh_WDTH -1:0]        I547f7a4c3801c1caa4587c9aef397652;
wire [flogtanh_WDTH -1:0]        I420e2c5a8745133f6263a71b458f1e2f;
wire [flogtanh_WDTH -1:0]        I8009d84fd826dd21eb7091744792f4a7;
wire [flogtanh_WDTH -1:0]        I4b8d520ee88fd39d83a16432e962f731;
wire [flogtanh_WDTH -1:0]        If724b1c92350989910925d275353e544;
wire [flogtanh_WDTH -1:0]        Ia3f7f07ddb09ea33218afe14281ac3c6;
wire [flogtanh_WDTH -1:0]        I26f4a180e992f5de04bc047f539bcb48;
wire [flogtanh_WDTH -1:0]        I25aefb53f59a00abe88b9dcf6be6907a;
wire [flogtanh_WDTH -1:0]        I83ca10d71caf5ac98fef3d45d228be8e;
wire [flogtanh_WDTH -1:0]        I22c3140a8db02352d2e2a2a11eeba117;
wire [flogtanh_WDTH -1:0]        Ib8407faa17d1e96cd317c65459c4fa71;
wire [flogtanh_WDTH -1:0]        I954dd66f60316803a8f13a39c460a39a;
wire [flogtanh_WDTH -1:0]        I73829d98e5e2f368c4a2020e3d7814be;
wire [flogtanh_WDTH -1:0]        I37b3988d699a1ed42923e3fd1584ecc0;
wire [flogtanh_WDTH -1:0]        I9a120c441f8d9ccb617057e042587ba1;
wire [flogtanh_WDTH -1:0]        If79bc5a35cb55036a367efb88c7d5510;
wire [flogtanh_WDTH -1:0]        I8064df8bc33998ad58d460afae699e48;
wire [flogtanh_WDTH -1:0]        Ideab06dc2448a6950cd1a06a0c90c2c6;
wire [flogtanh_WDTH -1:0]        If016e079d3b453444558706ef9073233;
wire [flogtanh_WDTH -1:0]        I1d7d7a68fc53b8be89c4637ac8f29380;
wire [flogtanh_WDTH -1:0]        I51cc187d91ee3c480a759104aed41b1b;
wire [flogtanh_WDTH -1:0]        Ib34ad1d14978608d1440f59998a31672;
wire [flogtanh_WDTH -1:0]        I4b8068a6a866c2424439b2956245ac8d;
wire [flogtanh_WDTH -1:0]        Id081512cd113e4d09df0fb13e443d76b;
wire [flogtanh_WDTH -1:0]        I60513d924016bd300559b7a1bea7f521;
wire [flogtanh_WDTH -1:0]        I57a0f8c3710cf8e216d6dc2420f7621c;
wire [flogtanh_WDTH -1:0]        Iec98284ab12724bb63360f29d00f1ecb;
wire [flogtanh_WDTH -1:0]        Iaa164a078c8cdaad694a053c9c1e0313;
wire [flogtanh_WDTH -1:0]        I3e3eba8135eb797d0a5e8ac1feefce0c;
wire [flogtanh_WDTH -1:0]        I7eb76b3d17296fdae702d8f820f1428d;
wire [flogtanh_WDTH -1:0]        I6aa98bc7265b8b7c25181a06e75c24c0;
wire [flogtanh_WDTH -1:0]        I00ecb5e329390023b318a2ceba0df231;
wire [flogtanh_WDTH -1:0]        I47f9c7018999e1cea25feddbe399e6b7;
wire [flogtanh_WDTH -1:0]        Iea32ebc385c6cfc9212ff37973a0a05d;
wire [flogtanh_WDTH -1:0]        I7224803ba8f0a16a7b2e969fe727bfa1;
wire [flogtanh_WDTH -1:0]        If845af0d620024f04525244753ba5d18;
wire [flogtanh_WDTH -1:0]        I65bc4e0d837f94c4301cb2c87e24969c;
wire [flogtanh_WDTH -1:0]        I08e907b0619bec3ef2cf4cb3779e0794;
wire [flogtanh_WDTH -1:0]        I444f8e61602b8994f7a01f3ebd4ac6ab;
wire [flogtanh_WDTH -1:0]        I68e5b12792a86dda0576742831d3b728;
wire [flogtanh_WDTH -1:0]        I86c51ec7ff965132e195835d21c24881;
wire [flogtanh_WDTH -1:0]        I72db05084d30d7c59ba1cb06d3b09400;
wire [flogtanh_WDTH -1:0]        I07aa1b2db5dedc3230dff10534311a56;
wire [flogtanh_WDTH -1:0]        Ib1f1aef6c0a9291553b62fd555feb2e7;
wire [flogtanh_WDTH -1:0]        Ia8809cc89c377e8b4109cdc8976daa54;
wire [flogtanh_WDTH -1:0]        Ib504b808f724ca6032e7c746517cd4fd;
wire [flogtanh_WDTH -1:0]        I7402dc21bfbc0af749dd8fb03c516a50;
wire [flogtanh_WDTH -1:0]        Ia47f7fb27f2d965cfd2989569c257356;
wire [flogtanh_WDTH -1:0]        I8ca06f4250a69dde75889f7a6ba3f456;
wire [flogtanh_WDTH -1:0]        If2b17f9e9186542117f43d0dd342326e;
wire [flogtanh_WDTH -1:0]        Ibab00faeaa6a7be99fa6a239193b92cb;
wire [flogtanh_WDTH -1:0]        I6c4ba0863ab4c8d1a56324a4d89ccbeb;
wire [flogtanh_WDTH -1:0]        I8e44b109466e00487db9dfb7ae225f89;
wire [flogtanh_WDTH -1:0]        I4dbd1bb8f1641f15e3a4f1e309962811;
wire [flogtanh_WDTH -1:0]        Ib3e38e46bfa9e1bdc032918269223b32;
wire [flogtanh_WDTH -1:0]        I26781ef851ed43c6f88ff1215cddca6b;
wire [flogtanh_WDTH -1:0]        I659fb1602b9d248940523c14c628ce86;
wire [flogtanh_WDTH -1:0]        Ia349e1f7c10a63ddccb3f300c73b4572;
wire [flogtanh_WDTH -1:0]        I1a264a901911abed928628d819c162b2;
wire [flogtanh_WDTH -1:0]        I50c4e1d3a3f63b93bc36b5141226fb3c;
wire [flogtanh_WDTH -1:0]        I2a53bd293919bc846ab816144b42592a;
wire [flogtanh_WDTH -1:0]        I12334038c2be8634c47869f397503019;
wire [flogtanh_WDTH -1:0]        I35ce9e616a3213f2b4ce0597a47f998c;
wire [flogtanh_WDTH -1:0]        I64692d5168554dfd7ce1c7a046aecf72;
wire [flogtanh_WDTH -1:0]        Ic3f28aa77fc84cb8e2fe43bac7ede253;
wire [flogtanh_WDTH -1:0]        Ia4b438844530fff602ea04e72b07db8d;
wire [flogtanh_WDTH -1:0]        I7f91c0e606b4082c6aec2e1f111079c5;
wire [flogtanh_WDTH -1:0]        I9574759e112f27778f3645d5d49126b7;
wire [flogtanh_WDTH -1:0]        I8e0d66c2112193437146e0f503623559;
wire [flogtanh_WDTH -1:0]        I2ffb7c2ad09bac694ef13ec41e5de327;
wire [flogtanh_WDTH -1:0]        Iabe6bf045784762fb6b97be3587fd68d;
wire [flogtanh_WDTH -1:0]        Ib190f589f4d663dbc0a3c166a8dcf5fa;
wire [flogtanh_WDTH -1:0]        I11f0fd7033065e1695d846f08d11aed5;
wire [flogtanh_WDTH -1:0]        I459c59ac61179d74170db53bf45ba89e;
wire [flogtanh_WDTH -1:0]        Ife1589d99f0764e3757de2a7d8b43008;
wire [flogtanh_WDTH -1:0]        Ie5e432a991aff25577639f1b4ffd594f;
wire [flogtanh_WDTH -1:0]        I7cb3f1f2e7f997b861d6c63d55c0f4ca;
wire [flogtanh_WDTH -1:0]        I72064a6a84ff956d76a5aa590bbc05a9;
wire [flogtanh_WDTH -1:0]        Iae2f185d6338026f3e37696327f214df;
wire [flogtanh_WDTH -1:0]        Iea74ecbac92e1b8f2ec7ad68d10b8e7d;
wire [flogtanh_WDTH -1:0]        I4da8f5b31f5cf7c70bba0cf661d727d8;
wire [flogtanh_WDTH -1:0]        I4f72d0db9fcc358c6fbec9964fbe0bbb;
wire [flogtanh_WDTH -1:0]        I46dd3a6d37d3df901689403a6215b65d;
wire [flogtanh_WDTH -1:0]        Ifd958901d2ea2284f506e04a058012fa;
wire [flogtanh_WDTH -1:0]        I84f43bb1814bdd83a682f7a859cfd611;
wire [flogtanh_WDTH -1:0]        Ie317bbd70b9092b840c0f2713204fb9d;
wire [flogtanh_WDTH -1:0]        I476ea921894e07d3f1d2ff3e7c3b660a;
wire [flogtanh_WDTH -1:0]        I2f9e56d570e72714a06c59aa9e4334c0;
wire [flogtanh_WDTH -1:0]        I5cc52764eb8a9961469e1892559ed7ee;
wire [flogtanh_WDTH -1:0]        I5b53fd45210b92703cb10d583f471ab9;
wire [flogtanh_WDTH -1:0]        I76f68c50b69a7545c0077f5333bfa3e2;
wire [flogtanh_WDTH -1:0]        I8edbe77bacf1975e014faeee6b861980;
wire [flogtanh_WDTH -1:0]        Id0bd4407ef72994435b3794096636553;
wire [flogtanh_WDTH -1:0]        I174fcbc2ee01fc55edbc8238e5da7f0c;
wire [flogtanh_WDTH -1:0]        I0879a96ba0ef5eb523ae807c40c66a63;
wire [flogtanh_WDTH -1:0]        Id4dc304aef5f35f6ceb91796c278e716;
wire [flogtanh_WDTH -1:0]        I8304ab4dc851d69a7ad7db75ced3eb9e;
wire [flogtanh_WDTH -1:0]        I0cbdfae6f75a639eb591d9c0022f5838;
wire [flogtanh_WDTH -1:0]        I24d773b608ba1ee21855540ee84028da;
wire [flogtanh_WDTH -1:0]        I088898ee932a96c14f2f0f568f5455b6;
wire [flogtanh_WDTH -1:0]        I9458b9a213600ce0c8c1d54d31c8c5c2;
wire [flogtanh_WDTH -1:0]        Ide0abde3644a4fafb436aa59768d016e;
wire [flogtanh_WDTH -1:0]        Idb6b8e6f2df9b8d96efa93830df86a71;
wire [flogtanh_WDTH -1:0]        I08581dc8d42be712cfb36d744f2786e0;
wire [flogtanh_WDTH -1:0]        I0a8fb8a7a28b364bc8cf49b96fdc66a4;
wire [flogtanh_WDTH -1:0]        I29fb3830a5fc5922f1ec687a38941e97;
wire [flogtanh_WDTH -1:0]        I938f8896ddbf95751aea2b327f5d40f0;
wire [flogtanh_WDTH -1:0]        I715d59fb27e519a9b76bdd8b5139a619;
wire [flogtanh_WDTH -1:0]        Ib5b964583d3ef33b47643ca212bc0ada;
wire [flogtanh_WDTH -1:0]        Ibe6a876a041198a581c95457a7d1fcf8;
wire [flogtanh_WDTH -1:0]        I4bae2a264af742ffe7be73f9a1129efe;
wire [flogtanh_WDTH -1:0]        Iec078a95a69b081cfb5e987ba9c5a613;
wire [flogtanh_WDTH -1:0]        I041c1a7ef6128c7a1a8f8593d4401f1b;
wire [flogtanh_WDTH -1:0]        I0e8f3f56bce3be1ee4d5f780a2f2a9fe;
wire [flogtanh_WDTH -1:0]        I22c6d2c87ef183ef45805a7c99a7e473;
wire [flogtanh_WDTH -1:0]        Ia73cacadbf80c0701a5b5b430c0d5c98;
wire [flogtanh_WDTH -1:0]        I45fef5261954fc84be265f39eb8f9647;
wire [flogtanh_WDTH -1:0]        Ic634d26fc09589a29a160e4efb5613a8;
wire [flogtanh_WDTH -1:0]        I3b292cf842e3a7ca9e6d0c4ab345446f;
wire [flogtanh_WDTH -1:0]        Ie1374cac341cf353b1863dae9f544e8b;
wire [flogtanh_WDTH -1:0]        Ie7bff678d39738eb49b599772586210a;
wire [flogtanh_WDTH -1:0]        Ia07447985347e9a7f3739bd98867cdfb;
wire [flogtanh_WDTH -1:0]        Ib9d80aab3818d682b54122974fa3a424;
wire [flogtanh_WDTH -1:0]        I2121318f589878b4a9260625f97de518;
wire [flogtanh_WDTH -1:0]        Iaa05186a94ba0559ab57ced9202ccefb;
wire [flogtanh_WDTH -1:0]        Ibd8424c228f87f85df3da6204edff2b5;
wire [flogtanh_WDTH -1:0]        I506f39735c3743b3705980c73295c035;
wire [flogtanh_WDTH -1:0]        I8a7fb51566bf215af214cd2fb5209974;
wire [flogtanh_WDTH -1:0]        I8f16ead6735608b15b364b9af9b3a22a;
wire [flogtanh_WDTH -1:0]        I7c0f872988488ac69815d288885dfd2f;
wire [flogtanh_WDTH -1:0]        Id07af023803badc88c51b891cad1b7e5;
wire [flogtanh_WDTH -1:0]        I3521b10b97b0e74888ce385cfc772945;
wire [flogtanh_WDTH -1:0]        Iecb522fa10764b2c0c044be6c1ca807d;
wire [flogtanh_WDTH -1:0]        I58f0b81a46549cab8e74ecbc285df23a;
wire [flogtanh_WDTH -1:0]        I58b9a09be96353ba6c18f310e1987742;
wire [flogtanh_WDTH -1:0]        I7095040b38bf9d6b5229c11d2a0d7c57;
wire [flogtanh_WDTH -1:0]        I86ced95bff4327e4ab07338663f82029;
wire [flogtanh_WDTH -1:0]        I675ab6c4fb93b006f3fcafc985fbc405;
wire [flogtanh_WDTH -1:0]        Ia802328754db2d72d6ec8e12a79b2341;
wire [flogtanh_WDTH -1:0]        I239a992ebb62899120a74b1c9e6cc4b4;
wire [flogtanh_WDTH -1:0]        I5b5a9fa50a6e4c7e07017249e5dee137;
wire [flogtanh_WDTH -1:0]        I927c870d09285dcb47e6d399f319471e;
wire [flogtanh_WDTH -1:0]        I73ef262450353dfcfabe3051ab0006f9;
wire [flogtanh_WDTH -1:0]        Ie23ed3ee61f468f59f2baf661cb7f85d;
wire [flogtanh_WDTH -1:0]        I959c5d62629333d1d60766a6d935ae4a;
wire [flogtanh_WDTH -1:0]        I68e58664be09261e5a80d6f8ecdd1b60;
wire [flogtanh_WDTH -1:0]        I659d579ea5b5d24ef0ccbb8160dfe2ae;
wire [flogtanh_WDTH -1:0]        Id2808e0f40992c79ead4da7c734e5b79;
wire [flogtanh_WDTH -1:0]        Icae3ba8a84ee6ee051a3caf210f47b51;
wire [flogtanh_WDTH -1:0]        Icb2b390266bff241a688961136db0f51;
wire [flogtanh_WDTH -1:0]        I92a005abe2d27beb2949fe29c0d8bc65;
wire [flogtanh_WDTH -1:0]        I54cfd68212d97a2cc8241ef429429453;
wire [flogtanh_WDTH -1:0]        I28fb1164936618d653aa7bf06c03b38f;
wire [flogtanh_WDTH -1:0]        I8d4e3962525c424786ae822a6981a5e6;
wire [flogtanh_WDTH -1:0]        I8720bdf2c91f113b39aa5b6f82421feb;
wire [flogtanh_WDTH -1:0]        I1a5f22b4e326d1684c0a8c7a7e754ab4;
wire [flogtanh_WDTH -1:0]        I07320e5fb3beddb93ae325a98c5e3782;
wire [flogtanh_WDTH -1:0]        I8c2e0c83a8204d6b21e0e3e458d56f05;
wire [flogtanh_WDTH -1:0]        Ib8b29bc86ad9c07d7ae5b358f66cb9ba;
wire [flogtanh_WDTH -1:0]        Ie0622ff815747e4a9f368c74787026ec;
wire [flogtanh_WDTH -1:0]        I8e2ed2040f5bf8ea125e5b953cf89300;
wire [flogtanh_WDTH -1:0]        I5ffed139764d90825b9f2eddacd0eddc;
wire [flogtanh_WDTH -1:0]        I4ad3a5b591cd6b13de04897fbbd068ec;
wire [flogtanh_WDTH -1:0]        I5a3297f48e1045273db6522744582b05;
wire [flogtanh_WDTH -1:0]        If5208f94e99b0e7ff353c048b55ad7ba;
wire [flogtanh_WDTH -1:0]        I9858bb2a3cc458aca5bf7eb077ee55dd;
wire [flogtanh_WDTH -1:0]        I66106fad536bb49418e7d09e3f4221ac;
wire [flogtanh_WDTH -1:0]        I6e7e27bb176196e4493bf9c45ca19719;
wire [flogtanh_WDTH -1:0]        I6af88c096ca3af849bbedb15b2ac7153;
wire [flogtanh_WDTH -1:0]        I4cff1804df738cbf4f940c775236df9c;
wire [flogtanh_WDTH -1:0]        I15d6e1e431457b954b5f86cd4fb16a77;
wire [flogtanh_WDTH -1:0]        I0c1e22375d5e023c24519901b92eceb5;
wire [flogtanh_WDTH -1:0]        Ifd67d6dec292171610a805560d7cb9a0;
wire [flogtanh_WDTH -1:0]        Ida5b16851dc06534844a0b037d74feb3;
wire [flogtanh_WDTH -1:0]        I681c4ec303ff366746d35234fe5a1ff4;
wire [flogtanh_WDTH -1:0]        Iac3cb5b4481687fcf430c8bf52cfb74d;
wire [flogtanh_WDTH -1:0]        I5df2eac3ace0bcef9e48b0850d975cce;
wire [flogtanh_WDTH -1:0]        Ia1499972c4995268acd828c1289f353d;
wire [flogtanh_WDTH -1:0]        Icf6f5254160a82036c4ba0367e8f0404;
wire [flogtanh_WDTH -1:0]        Ie559401a3a913400dc5e3e5641297fa6;
wire [flogtanh_WDTH -1:0]        If1de12bbb90e49cc1b28eafc2aa551e5;
wire [flogtanh_WDTH -1:0]        Ie0667fbe76244eaec0b155d69dcc9447;
wire [flogtanh_WDTH -1:0]        Ibf9f7f1f6a759af21ac82d6e6ff7df43;
wire [flogtanh_WDTH -1:0]        I1d0f031e8ae9c0335d501d1565118220;
wire [flogtanh_WDTH -1:0]        Ie44bc9632854c4c2077bcec5f46d29ad;
wire [flogtanh_WDTH -1:0]        Ie2c801b2de066c3218d7312615b7bfda;
wire [flogtanh_WDTH -1:0]        I97ae894cd928e17cad4c4631aec2c7a0;
wire [flogtanh_WDTH -1:0]        I64c4bb0d40d80ec52aab61ce46954f43;
wire [flogtanh_WDTH -1:0]        I500a903104b4b532b3c07d1640e80b55;
wire [flogtanh_WDTH -1:0]        I512f57a40c7c8cb2f040bdde73e44ca3;
wire [flogtanh_WDTH -1:0]        I1d3ae54c8fa3d87a39e3a51018a20727;
wire [flogtanh_WDTH -1:0]        Id60cbf534604e5dba988050ef5abe625;
wire [flogtanh_WDTH -1:0]        I23d3b6da58b66185ddb3c5eae0f68dae;
wire [flogtanh_WDTH -1:0]        I37998a91d20db2248ebdd8e661d42f70;
wire [flogtanh_WDTH -1:0]        I88b1352db9aa35be019bc0f345c7131e;
wire [flogtanh_WDTH -1:0]        Ib65ff82aff398f6ff7ba711a36f41ee4;
wire [flogtanh_WDTH -1:0]        I1115071c073981f4db4917844fb12a73;
wire [flogtanh_WDTH -1:0]        I3d1dd8b9c7c6d3913f7ac369ad7e625c;
wire [flogtanh_WDTH -1:0]        Ia9e4e593fd82657c81aeea8fbcd1194b;
wire [flogtanh_WDTH -1:0]        I097722547450582dc5776bdaff914741;
wire [flogtanh_WDTH -1:0]        I22300986ed621a97a6dac1f3b4d59b8e;
wire [flogtanh_WDTH -1:0]        Id4a213e494f9c9be0fd1a307e87c756a;
wire [flogtanh_WDTH -1:0]        Icc08ab7c64b40e53278a93f4ae0f9209;
wire [flogtanh_WDTH -1:0]        I21594c8b0169efd7c2aa6cbc31f4a901;
wire [flogtanh_WDTH -1:0]        I8cc9f5531f2675b3058df110912551b6;
wire [flogtanh_WDTH -1:0]        I15022e1b349eee259d3567837283dbf6;
wire [flogtanh_WDTH -1:0]        Icdba6332ba9ea91ffefd690150fba09f;
wire [flogtanh_WDTH -1:0]        I1070940dc2ef6e8ee3d1227ec9ff3162;
wire [flogtanh_WDTH -1:0]        Idaef789d04cd5c6291dae88f616460e6;
wire [flogtanh_WDTH -1:0]        I8922cc37cde6ba132f632743113e42af;
wire [flogtanh_WDTH -1:0]        I016cb9c8307b28a7cabf9a91e8da03d6;
wire [flogtanh_WDTH -1:0]        Ia66c399023e500ed67197dcf236f5d42;
wire [flogtanh_WDTH -1:0]        I54517f62dd6f2e7de7d522dfc506383e;
wire [flogtanh_WDTH -1:0]        I1171dc208d5db1024dc3f09a90c78ca0;
wire [flogtanh_WDTH -1:0]        I6b0c1ef6f0a94adaf62425829edf28dd;
wire [flogtanh_WDTH -1:0]        Ic28b148967a5b3d05409976fa9001ac8;
wire [flogtanh_WDTH -1:0]        I067ce754b1084de762c33b295f2f47b2;
wire [flogtanh_WDTH -1:0]        I79fe46308b93fbb24245fe1c75edf4a5;
wire [flogtanh_WDTH -1:0]        Ib2fe88cfe23c363993dfcb7722c4fef0;
wire [flogtanh_WDTH -1:0]        I3bfcd63e92f1949234ab1d2701dbb499;
wire [flogtanh_WDTH -1:0]        I71f836227a1f7f81500a6c980c06f1f7;
wire [flogtanh_WDTH -1:0]        I5e2331edf6e881e9f3a8c47eebda0ac4;
wire [flogtanh_WDTH -1:0]        I6faf34757a61a0b64e61ba059aca33fa;
wire [flogtanh_WDTH -1:0]        I4b66c202450986ef0df05e979cc8bc7f;
wire [flogtanh_WDTH -1:0]        Ib1821b79b79aadf1486fe1e2df2f297c;
wire [flogtanh_WDTH -1:0]        I737daf208eccf95feb3192897586cdce;
wire [flogtanh_WDTH -1:0]        I84daf07d3f3790c691b9192f7e2018c1;
wire [flogtanh_WDTH -1:0]        I29c8133231cfda17668bbe7b692bdfe2;
wire [flogtanh_WDTH -1:0]        Ib4b3ed1f9d1dee96a3ec846424412e2f;
wire [flogtanh_WDTH -1:0]        Id9d56f09595e80d66c2ac300f7d1d972;
wire [flogtanh_WDTH -1:0]        Ibe73f00bb6f1494ede2e6f11f5e7d3f8;
wire [flogtanh_WDTH -1:0]        I97e89a2ee18d2688d7c1a640318a1e0d;
wire [flogtanh_WDTH -1:0]        I1542461b996a466d7d3d50bb48ebd690;
wire [flogtanh_WDTH -1:0]        Ife123bf57fe693dabe6aeaa236c4e058;
wire [flogtanh_WDTH -1:0]        If97a5a2c523f51c5881496c5dc8ad11e;
wire [flogtanh_WDTH -1:0]        I0c0d844fe3b7d35c1ed6bd7cc4e0dc24;
wire [flogtanh_WDTH -1:0]        Ie19ea558cf2a95ca0c8ae769a809d908;
wire [flogtanh_WDTH -1:0]        I2d9632ae6a0f3ba44c3da8f56ba3fedf;
wire [flogtanh_WDTH -1:0]        I6532e6299b8c1fdf7f61b3a44b61c35c;
wire [flogtanh_WDTH -1:0]        I38cc7b117c0bcd5e3060cd370d710d7e;
wire [flogtanh_WDTH -1:0]        Ic7102fb8b5df222fff6151e8794bec3c;
wire [flogtanh_WDTH -1:0]        I793ddbf6a5d026a57ab72984ca19deac;
wire [flogtanh_WDTH -1:0]        I1f97ea0e7bf46382824cbffc3e94e9df;
wire [flogtanh_WDTH -1:0]        I79458089b042e181e37cc44c06d08681;
wire [flogtanh_WDTH -1:0]        I801dfe17655932ad8fe9702cbaad270f;
wire [flogtanh_WDTH -1:0]        I42460fae0acff25fa2b829e39ddcc4fd;
wire [flogtanh_WDTH -1:0]        Idbd834f0c907b233a8eff58eaca28863;
wire [flogtanh_WDTH -1:0]        Id3670a6f05d40ab69624544de92b9c64;
wire [flogtanh_WDTH -1:0]        Ic69e0c34630bde15f4172714bc3d92be;
wire [flogtanh_WDTH -1:0]        I81800fb49855a4fd2737faa07ff15d29;
wire [flogtanh_WDTH -1:0]        I465a735c8e94ddbfdbaeb2a7652e481e;
wire [flogtanh_WDTH -1:0]        Ibfe325e48511372569e0d98d9c4e70e3;
wire [flogtanh_WDTH -1:0]        Id1c6a3f52dd7972f47cbd8103ace643f;
wire [flogtanh_WDTH -1:0]        I326660e98f61bb2ced4c23c7bcc9324a;
wire [flogtanh_WDTH -1:0]        I26b9e2d073b20376980662c249bf9d43;
wire [flogtanh_WDTH -1:0]        Ic6fa98631d742b27f252fe7c95caef55;
wire [flogtanh_WDTH -1:0]        Id4cc1b15055941d401ded6ff8b777461;
wire [flogtanh_WDTH -1:0]        Iab6d0f72579687407e029c630b107f7d;
wire [flogtanh_WDTH -1:0]        I064bd1f4b7fa40b2cae3ea361edf9167;
wire [flogtanh_WDTH -1:0]        I19eae741ef89baa1a64c403fb29f14f4;
wire [flogtanh_WDTH -1:0]        I4b5aadc25b0ed6811a665b33d6c4ae2a;
wire [flogtanh_WDTH -1:0]        I749b9c345f23aae03c595a2c76126ecb;
wire [flogtanh_WDTH -1:0]        Ic883bcc70572a237ba0e3d465337bc59;
wire [flogtanh_WDTH -1:0]        Idc77c7d5123717fc2596a51d904c6d82;
wire [flogtanh_WDTH -1:0]        I7181ab1d663b0cbe30861e29fc3f8532;
wire [flogtanh_WDTH -1:0]        I779da979707d9712c1626d6025f97599;
wire [flogtanh_WDTH -1:0]        Id3fbb6d083344684de89d99c040b2100;
wire [flogtanh_WDTH -1:0]        I97aede8502e443f98938487a5a5c072c;
wire [flogtanh_WDTH -1:0]        Iee8d139aa5a8ae046f5019abecdbc3c4;
wire [flogtanh_WDTH -1:0]        Ie7820d1a242bc28c19ec32d2c91e47b7;
wire [flogtanh_WDTH -1:0]        Idc0bfe36a3a9b3006a04d5dfc31b8107;
wire [flogtanh_WDTH -1:0]        I82a14e1ee4723e7d9a13c1f2b8b13691;
wire [flogtanh_WDTH -1:0]        Ia2462ec52aaccc97597d1dfc2e33b7e2;
wire [flogtanh_WDTH -1:0]        I77a94cd9186ca546ca9664942ea3537f;
wire [flogtanh_WDTH -1:0]        I8048bbe27b49b9d248fee919be6dc977;
wire [flogtanh_WDTH -1:0]        I3c0ddec25c53c166d30eb78d4518840e;
wire [flogtanh_WDTH -1:0]        I838d1cc5e9ca5058c25223ec53d9c34f;
wire [flogtanh_WDTH -1:0]        I98bbe3b75958f10195dee6460cf2aca6;
wire [flogtanh_WDTH -1:0]        Id9e5147e089e6e52ef2a687d76534f16;
wire [flogtanh_WDTH -1:0]        If6d436031f68ef587750c5c1dfcfffc2;
wire [flogtanh_WDTH -1:0]        Ia043941abbcf10c16f086fe8d61dd456;
wire [flogtanh_WDTH -1:0]        I461398638cb8280f1779915298540b00;
wire [flogtanh_WDTH -1:0]        I625ab32380498dfbf9d3290c2053bf3d;
wire [flogtanh_WDTH -1:0]        I20c65000bbc10299168af7390776a03c;
wire [flogtanh_WDTH -1:0]        I903f7844e55d1cd6969352490c275c8e;
wire [flogtanh_WDTH -1:0]        Ia840e19ca36795a50ab1a6e6a1729edb;
wire [flogtanh_WDTH -1:0]        Ie5951bc919195ba594fe87375ad41269;
wire [flogtanh_WDTH -1:0]        I7d98d1e5f07fccff5f20eaca6363c700;
wire [flogtanh_WDTH -1:0]        Ieeed8d4eebc0adea7ee0af6a5dbe045c;
wire [flogtanh_WDTH -1:0]        I97a75b8625ae2a143cf364790ae77753;
wire [flogtanh_WDTH -1:0]        I266cd5f0a56cd5171da8d59df0042d5d;
wire [flogtanh_WDTH -1:0]        Idbea892c8109117f90b453efe8ae25af;
wire [flogtanh_WDTH -1:0]        Ie5a57c603ad520441bc5819c81fb877f;
wire [flogtanh_WDTH -1:0]        Icfc1c6d96a3598af73e99a350c387d72;
wire [flogtanh_WDTH -1:0]        I17ac503f4f952f9e2fcdea3f955cc1a9;
wire [flogtanh_WDTH -1:0]        I523e9b6f828ec7f166750112f8a3f676;
wire [flogtanh_WDTH -1:0]        Id8b704aada09411d5f5153d088c1c613;
wire [flogtanh_WDTH -1:0]        I79259217f63b2f6263552c434d0e5c93;
wire [flogtanh_WDTH -1:0]        If64a200b2dac7049b77e5b6bb03b9cc3;
wire [flogtanh_WDTH -1:0]        Ice6db5ba70d3c7499df6723a2df56bfe;
wire [flogtanh_WDTH -1:0]        Iee1b48cae01fe51344b8d662ace9c6f1;
wire [flogtanh_WDTH -1:0]        I28aa517220bf597cf898660f698ef19d;
wire [flogtanh_WDTH -1:0]        Ic879cd355d61eb021250d62841115a52;
wire [flogtanh_WDTH -1:0]        I07048dc5cbe24ff72d24902d572face0;
wire [flogtanh_WDTH -1:0]        I46e2d889b9ba7eccad5529200852ca17;
wire [flogtanh_WDTH -1:0]        Iab3876e5107e3a56b1fafe41e16d9482;
wire [flogtanh_WDTH -1:0]        Ia4e080f13520998be95b64eb883f8e32;
wire [flogtanh_WDTH -1:0]        I511a55c2f4d6d3727dff5825597f55a9;
wire [flogtanh_WDTH -1:0]        I2ad2ede07f1ffac643211e88bf8ddbd6;
wire [flogtanh_WDTH -1:0]        I2493237a24acdcab8b5bda10e804a5cf;
wire [flogtanh_WDTH -1:0]        I5bc390dc300be5f8bc85f928cca1cd0b;
wire [flogtanh_WDTH -1:0]        I03829256e357ac17c7ca7cae2f980f41;
wire [flogtanh_WDTH -1:0]        I3e7efaed64fd3c276e882ab38109d538;
wire [flogtanh_WDTH -1:0]        Iae32c44b88fe7ddb5d4f19cf8fff3ba6;
wire [flogtanh_WDTH -1:0]        Ib4738fe629dbe40eefed821b40ab93c8;
wire [flogtanh_WDTH -1:0]        I3bdc5ba374f85dc61346e4868c41a6bf;
wire [flogtanh_WDTH -1:0]        I30268ed341753c3ab53b65ad43e94923;
wire [flogtanh_WDTH -1:0]        I557ef77ce931535467a07a8d70145f55;
wire [flogtanh_WDTH -1:0]        I2f10be9cbe2a935475077c0218031a5a;
wire [flogtanh_WDTH -1:0]        Ib4695d4389db72c5ac7e31809072c290;
wire [flogtanh_WDTH -1:0]        I41d598b80334ab12e5f53b2a6c721517;
wire [flogtanh_WDTH -1:0]        Ie81315a3a14a5ef879d8e3f405936365;
wire [flogtanh_WDTH -1:0]        I94b3d895ee69e3ab482ff1aa0798c92a;
wire [flogtanh_WDTH -1:0]        Ia7520053a7c4a94437c6a780b03a28a5;
wire [flogtanh_WDTH -1:0]        I24a25d4725db6bcb4732fa21bc861736;
wire [flogtanh_WDTH -1:0]        Ic308a5413f38b96d244cac3b0bc9462c;
wire [flogtanh_WDTH -1:0]        I1877b73e028c908de9dc734b93cbf8bb;
wire [flogtanh_WDTH -1:0]        I034fb3850485fae2d1358041a1c41888;
wire [flogtanh_WDTH -1:0]        Ic99b64430e5dfdabe3634fbddeb41b3c;
wire [flogtanh_WDTH -1:0]        I0e7079db66c15210046b997f319ece89;
wire [flogtanh_WDTH -1:0]        I3c0ddec6d702a344930fd04f923bb2f1;
wire [flogtanh_WDTH -1:0]        I9a5388f8aa6e9924a309aa8db4c1983b;
wire [flogtanh_WDTH -1:0]        I41829e511abe1ddf9b67f899143db19a;
wire [flogtanh_WDTH -1:0]        Ief76663994991118b1899ea4ddf4527d;
wire [flogtanh_WDTH -1:0]        I41961139f5b650e4f4ba5c2eadda6702;
wire [flogtanh_WDTH -1:0]        I6fb63ea54e492bdbc6d1145affc683e9;
wire [flogtanh_WDTH -1:0]        I8ef0ac3bf43f16d2edf5a5045b0eb498;
wire [flogtanh_WDTH -1:0]        If83ce1cbe3a73472419520c225b288a6;
wire [flogtanh_WDTH -1:0]        I4084e3c9ba635fc4a8d281015bdeb33a;
wire [flogtanh_WDTH -1:0]        Id1df78ab32daf524b77c0431c782f2bf;
wire [flogtanh_WDTH -1:0]        I199a14038a0ff6ac25dab60162f8c6c9;
wire [flogtanh_WDTH -1:0]        Iff142b88493149045fc0de355b767c16;
wire [flogtanh_WDTH -1:0]        Ic6859263f79d29d5f4896d85367be2bf;
wire [flogtanh_WDTH -1:0]        I28c3818247c7c6de11790f6692882b5a;
wire [flogtanh_WDTH -1:0]        If0af3259e321390fffe518318f0f2545;
wire [flogtanh_WDTH -1:0]        Ib451127b69a0a800332a712af77c6d29;
wire [flogtanh_WDTH -1:0]        Icafbf36da24f4db99e0ce4eeca6ca338;
wire [flogtanh_WDTH -1:0]        I3d601db540da359ae4d22f960d3d5af8;
wire [flogtanh_WDTH -1:0]        Ia614303d31afc0ef4f15ec5b43231cd8;
wire [flogtanh_WDTH -1:0]        I2c1f2476efe593829ade470fe8ec2526;
wire [flogtanh_WDTH -1:0]        I28ff2f86da2016b00bd0c21cbd1b4530;
wire [flogtanh_WDTH -1:0]        I7e685b06df8a8c2ac351fa9f9b76a81d;
wire [flogtanh_WDTH -1:0]        I2b8c969c11b4117c96470f4f6ed6963a;
wire [flogtanh_WDTH -1:0]        I1338d211b5d2d409bfe0df76d2ca2701;
wire [flogtanh_WDTH -1:0]        Iea563639beb7fcb0291b5dc1410951d1;
wire [flogtanh_WDTH -1:0]        Ia40dad546d9c852e2fa8942c62a1c1f8;
wire [flogtanh_WDTH -1:0]        Ic1b35046657e23f42199e39343a652a8;
wire [flogtanh_WDTH -1:0]        I0b0dd019d8bd24684403a29aed668b6d;
wire [flogtanh_WDTH -1:0]        Ie7b26120ee77b43574c1ca171d7ec15f;
wire [flogtanh_WDTH -1:0]        I66a304016a9adfd85a2abb6f8fd39afc;
wire [flogtanh_WDTH -1:0]        I2ed61ced1577d905da91d97592006ed5;
wire [flogtanh_WDTH -1:0]        I177be24718c59688752097fe2a4085c4;
wire [flogtanh_WDTH -1:0]        I332dc26a52194745d19c4d8468e42864;
wire [flogtanh_WDTH -1:0]        I7e66a42eb7cdb820cd1297c39f0625e8;
wire [flogtanh_WDTH -1:0]        Ibb4fefe05e94e055e86a743c40fb1c5e;
wire [flogtanh_WDTH -1:0]        If2021f0735c6c5649ebac0d230fda87c;
wire [flogtanh_WDTH -1:0]        Ia56a76a20d4f11b0e80cbe31820a6977;
wire [flogtanh_WDTH -1:0]        Ie1bf5d97b8f679095d2442bbf9f95608;
wire [flogtanh_WDTH -1:0]        I054ebc7f9e3da325ba0c6e329f2ee770;
wire [flogtanh_WDTH -1:0]        I632469889d6bb1c268b45fb805467ebd;
wire [flogtanh_WDTH -1:0]        I3361df26cc86ca8be1653d9376d0c8e0;
wire [flogtanh_WDTH -1:0]        Ie230ba3c73808e102eee9e5868595e7c;
wire [flogtanh_WDTH -1:0]        I586fbde80f0130c4a6ead49de11efdd9;
wire [flogtanh_WDTH -1:0]        Ie1e9326e4eee006ec07abb6bb7d269a5;
wire [flogtanh_WDTH -1:0]        Ifa087137c8a6028b13bfa95aba19fc34;
wire [flogtanh_WDTH -1:0]        Ica4ec1647bdb5a3aad6db6b447bd7995;
wire [flogtanh_WDTH -1:0]        I51a3a6c79c488c092394375891775be3;
wire [flogtanh_WDTH -1:0]        Ia17295aec0a40c2b46a595dacfede2d5;
wire [flogtanh_WDTH -1:0]        I01a7ebdc760227ee40b85828e28238a9;
wire [flogtanh_WDTH -1:0]        I4c6d3d6fc2d10066a744fdd9405a7902;
wire [flogtanh_WDTH -1:0]        Ib3f9e4c05e363069775e5de9d240b3dc;
wire [flogtanh_WDTH -1:0]        Ia9c043c5e8873fd13e39cf6bd8136c51;
wire [flogtanh_WDTH -1:0]        I18664482dcc1371fa4b915af96070539;
wire [flogtanh_WDTH -1:0]        I2e802c75c6ce34b05943b678ecbfacb1;
wire [flogtanh_WDTH -1:0]        I6a41c6cf78cb25ad1c47550756449002;
wire [flogtanh_WDTH -1:0]        Ieb3f28762410fb40a0c8a8556b4b3ca0;
wire [flogtanh_WDTH -1:0]        Iaf660a97d66e0d7f8e26f65229b7683f;
wire [flogtanh_WDTH -1:0]        Ie3e0c0e40c7a67ce7f957e74bd2a895d;
wire [flogtanh_WDTH -1:0]        I7ded197ff64af1bce0e0d85705900a42;
wire [flogtanh_WDTH -1:0]        I491f2373b2df19a4c22e1787ef034179;
wire [flogtanh_WDTH -1:0]        I7c06179d5424165f8a805754834fd98c;
wire [flogtanh_WDTH -1:0]        Ief96603d41b4f670d2bbfa3d3875c903;
wire [flogtanh_WDTH -1:0]        Id364f2a517a0f3109564a025ffd8eec3;
wire [flogtanh_WDTH -1:0]        I7a029c27d92754041eb6d605837238dd;
wire [flogtanh_WDTH -1:0]        Ie3ea12584ed3e255073776620d778f06;
wire [flogtanh_WDTH -1:0]        I00dad36628d2fa923120fdaa79bf0045;
wire [flogtanh_WDTH -1:0]        I38d885c58b4f7333c679b0b5783418df;
wire [flogtanh_WDTH -1:0]        I3707f68de059df0af5c652fc0478e543;
wire [flogtanh_WDTH -1:0]        I69251440f80eb2e177307aec4cb0111f;
wire [flogtanh_WDTH -1:0]        I94af4b6b9dc11935db54ba872889392d;
wire [flogtanh_WDTH -1:0]        I0a9bcd4a3b79b003b5df8afa0d6b6782;
wire [flogtanh_WDTH -1:0]        I38e2dbba093928b874d447362d89b291;
wire [flogtanh_WDTH -1:0]        I36569656996bf98bce33b2d7a4b79def;
wire [flogtanh_WDTH -1:0]        Ia48f0029e9e76386f3dd70aacd9adbfa;
wire [flogtanh_WDTH -1:0]        I7e408a50d0511909aeb57d5a00535e80;
wire [flogtanh_WDTH -1:0]        Ic2b20168744fafbe15037ed7fa83da72;
wire [flogtanh_WDTH -1:0]        Iacc6f48dd92dc515be06a681cc5b56e9;
wire [flogtanh_WDTH -1:0]        I62fdc8936121a2707d94cf3bd6e660ac;
wire [flogtanh_WDTH -1:0]        Icafa051878ad3421c31ed2550ea09945;
wire [flogtanh_WDTH -1:0]        Ia0932b3fd6a5ae6da2bacd2b86ba3a43;
wire [flogtanh_WDTH -1:0]        If4e4f2776b1467e4f03bf15ff5f43c04;
wire [flogtanh_WDTH -1:0]        I9fce6091885f1bb97d29fb1f543b1a38;
wire [flogtanh_WDTH -1:0]        I9387cd07e38260005bb3e41807d2d794;
wire [flogtanh_WDTH -1:0]        Ib402cdbfaa9900820b85bd625415c547;
wire [flogtanh_WDTH -1:0]        I8bede290f421e6a05e49244f0d1d3d9b;
wire [flogtanh_WDTH -1:0]        I518a2736384c14c02f27bfa3d8ea7aff;
wire [flogtanh_WDTH -1:0]        I6d8c2489fdeb42411f2e12bfa30752d2;
wire [flogtanh_WDTH -1:0]        I847cf7ff866f8a666872c12d6b67b1b1;
wire [flogtanh_WDTH -1:0]        I082715d1b8943faf11d464087542a83e;
wire [flogtanh_WDTH -1:0]        I9e45e3d7117ce48cdbfc5db8c0ccfcf4;
wire [flogtanh_WDTH -1:0]        I4de91d9613edc5c4d096b717d9df5de4;
wire [flogtanh_WDTH -1:0]        I380ff8528cdba4026fac3c4eda8b2c52;
wire [flogtanh_WDTH -1:0]        Ifb2a91a74b87c75592cb046b9bfd9c8b;
wire [flogtanh_WDTH -1:0]        Iee8f9b0654f6f6797f11cae0947e454e;
wire [flogtanh_WDTH -1:0]        Ie21cffaecd7fe37601dcaef49a0d6cc3;
wire [flogtanh_WDTH -1:0]        Ie3e54a4700d8d0f6478187e06cb6f85d;
wire [flogtanh_WDTH -1:0]        Ia648c9d395ad2727209229807b4224fb;
wire [flogtanh_WDTH -1:0]        I8c0069e8756bcff203ce21ae3170aa42;
wire [flogtanh_WDTH -1:0]        Ib415da845b88e5a8261beaf88b7ec804;
wire [flogtanh_WDTH -1:0]        I856eada207c5006beb8f83f01d5d74c9;
wire [flogtanh_WDTH -1:0]        I6dffcf934a74385aa716db9d7fa29ed1;
wire [flogtanh_WDTH -1:0]        I79a46279070c53678a5af54f661c5821;
wire [flogtanh_WDTH -1:0]        I13383df545ed8620a17a4fc2493cd770;
wire [flogtanh_WDTH -1:0]        Ica807adc510a2e32580ca77c18ea0b45;
wire [flogtanh_WDTH -1:0]        I87ea43bfae8fad4e4c26741fd2de5b41;
wire [flogtanh_WDTH -1:0]        Ia8094903aed8dd0ce8e9ff459a5287b0;
wire [flogtanh_WDTH -1:0]        I6d2022ba184980b8e5bc5edb4f4b0ff3;
wire [flogtanh_WDTH -1:0]        Ie018f3003c5f124bddd13c359257bf35;
wire [flogtanh_WDTH -1:0]        I68f98b68c9a3836d0c7dc152a2d441da;
wire [flogtanh_WDTH -1:0]        Ice18bceb10fec484ffc96155e14c4974;
wire [flogtanh_WDTH -1:0]        I2dc3cec85c37aa943f01df545f952e05;
wire [flogtanh_WDTH -1:0]        Ib484aa64b795f7e36198b800f302164f;
wire [flogtanh_WDTH -1:0]        Ieed49c262f87c86b30d94e9842525ab0;
wire [flogtanh_WDTH -1:0]        Icdb143a4ce96029c2441758bf2edd7b0;
wire [flogtanh_WDTH -1:0]        Ib9ab475010c98fc4e06df5c98944387a;
wire [flogtanh_WDTH -1:0]        I3a76f70ca3bfbcacc6f3342aa71f1912;
wire [flogtanh_WDTH -1:0]        If7c8bdd5bae4a1bffd4bd2c8015bb738;
wire [flogtanh_WDTH -1:0]        I9470c7ab9634c01bb832c9e4ff5496bf;
wire [flogtanh_WDTH -1:0]        I6463249144cd032e1c5af9e2987254b3;
wire [flogtanh_WDTH -1:0]        I218ee96418a4f5d734d3d71685bc09c7;
wire [flogtanh_WDTH -1:0]        I5f9e468fc1bc199574d719d866d52dfc;
wire [flogtanh_WDTH -1:0]        I924514226fdb5bac110a2650bcb2e85f;
wire [flogtanh_WDTH -1:0]        Ie69f792c606c3162052840dec732ef99;
wire [flogtanh_WDTH -1:0]        Idc57f37015a48393608e2b026bc7065c;
wire [flogtanh_WDTH -1:0]        If874254c3c6813ff0d5184b574cb613d;
wire [flogtanh_WDTH -1:0]        I41af7e4c97fc04154fe6de66b82499f5;
wire [flogtanh_WDTH -1:0]        I90969c917df8480d379afef834c1a253;
wire [flogtanh_WDTH -1:0]        I972bee4216f8e532e8fa4bd25fbb9c57;
wire [flogtanh_WDTH -1:0]        I07280ae3417855f994980fbb95696fc6;
wire [flogtanh_WDTH -1:0]        Ib303ea0240e7ab5f000dd10e975b2274;
wire [flogtanh_WDTH -1:0]        I852c62fffff0fd7bf06939d75fada3eb;
wire [flogtanh_WDTH -1:0]        I5971253546899e9a82f387d5eabcc7b3;
wire [flogtanh_WDTH -1:0]        I9e0a2da5a82f1b509bd502554f4760aa;
wire [flogtanh_WDTH -1:0]        I1fc36e6f738fab96df356979e1e3a612;
wire [flogtanh_WDTH -1:0]        I6293c2b405087f14b42b423336f6990c;
wire [flogtanh_WDTH -1:0]        Ie2d8c84d8c9a4c8f637068a2ae39fdde;
wire [flogtanh_WDTH -1:0]        I70e8d96970e69bc828a6aea5ade3bdd1;
wire [flogtanh_WDTH -1:0]        I114c595caa67a3f777f087a634130a6d;
wire [flogtanh_WDTH -1:0]        I0380003f741eedb994793c2cb7e6c5c3;
wire [flogtanh_WDTH -1:0]        Idad14b6383b9af54eb35e72ff3d10035;
wire [flogtanh_WDTH -1:0]        Ia884fcfa49cfe0b404bf49b99d7381aa;
wire [flogtanh_WDTH -1:0]        I46e9c76b19ed1ff21f102efe6ee5c732;
wire [flogtanh_WDTH -1:0]        Ie4ecd4c122ea5b478f3d7d2d632b8bf4;
wire [flogtanh_WDTH -1:0]        Ic75b8bbb1b80001ec188a0cd25623420;
wire [flogtanh_WDTH -1:0]        I82e534ecaabf5af6a9b6a567b862800a;
wire [flogtanh_WDTH -1:0]        Idc7df6877bdb7e7d392307d78183d31c;
wire [flogtanh_WDTH -1:0]        I1c9684b45467216a18a3a0d93b555b60;
wire [flogtanh_WDTH -1:0]        Ib8b95ece5da3877b261a06e6d0571921;
wire [flogtanh_WDTH -1:0]        Ice212c509101d6d41b52ea0cb85dacc0;
wire [flogtanh_WDTH -1:0]        Ic99654bf4833c9132912eeb4c0dc92fa;
wire [flogtanh_WDTH -1:0]        I37ee7a2fab22cf8e6452fb408b849595;
wire [flogtanh_WDTH -1:0]        I2461055ef9b1aa2ffca0f5cac3300e71;
wire [flogtanh_WDTH -1:0]        I0ec18ade132eede6849e0607af608726;
wire [flogtanh_WDTH -1:0]        I2bc3ffbe5b42b0833206437d3863278e;
wire [flogtanh_WDTH -1:0]        I4651eab27cb766a1792f9564bcb2764a;
wire [flogtanh_WDTH -1:0]        Id5e02d4c48fa6c3b0d45a9e66f09448f;
wire [flogtanh_WDTH -1:0]        Ibbdbc4e4fc2ee018a0e7a4da29e85b56;
wire [flogtanh_WDTH -1:0]        I40e99289d5762e77a3766eb8251eef00;
wire [flogtanh_WDTH -1:0]        Ic67b9e090d6815b2a745bdc4983f9c69;
wire [flogtanh_WDTH -1:0]        I20beb3fdbe91936f74a200cd8ec9817b;
wire [flogtanh_WDTH -1:0]        I8327267045af5da02c066a5eab25f13a;
wire [flogtanh_WDTH -1:0]        Id435b68afb53bef4afc7b70a9512e955;
wire [flogtanh_WDTH -1:0]        Id91ef7e27c689cdf5ce50d705017e40e;
wire [flogtanh_WDTH -1:0]        I0cf5cb4cd472502b84dbf6fe1af0be78;
wire [flogtanh_WDTH -1:0]        I60498760f3c03cf92ceeb99c5096fe54;
wire [flogtanh_WDTH -1:0]        Iacf6340a29a5592b61ea875304a2de48;
wire [flogtanh_WDTH -1:0]        I63169dbc533400e0db5e37a8ebeca1aa;
wire [flogtanh_WDTH -1:0]        I5dfc71255cba279420b7545df4d35c40;
wire [flogtanh_WDTH -1:0]        I150f11a565ad39c59d8f9e4c94d397e2;
wire [flogtanh_WDTH -1:0]        Ibadcb205c7e9a0f3345cac7eb41b5985;
wire [flogtanh_WDTH -1:0]        Icadb816a238ba165425e5a30bd0bb8e6;
wire [flogtanh_WDTH -1:0]        I762b2abb876381eff6de97cef0798405;
wire [flogtanh_WDTH -1:0]        I3b55785b9625ac53f6c00ba5a10a481b;
wire [flogtanh_WDTH -1:0]        Ib3e7633767b6e09e4ee54f6feaddd31e;
wire [flogtanh_WDTH -1:0]        If7317c81c9b6503386cab33fa812e80e;
wire [flogtanh_WDTH -1:0]        I3f193e9c265c1dfaeada63d59db5b79f;
wire [flogtanh_WDTH -1:0]        I095672e79ca3a6dd8589b7821f06cdb9;
wire [flogtanh_WDTH -1:0]        Ie72268e979cf069b88f6eadde789e5ab;
wire [flogtanh_WDTH -1:0]        Ibf2f43980e835dd7ae7535957e3ec131;
wire [flogtanh_WDTH -1:0]        I5732fdb805258fc13c8ba4aaf56574ca;
wire [flogtanh_WDTH -1:0]        Iaa980a50205025e3e1b09c6ce8ee53dd;
wire [flogtanh_WDTH -1:0]        I3afe987d8f2c93cc19534a3221d1939c;
wire [flogtanh_WDTH -1:0]        I829aa657f0dd13c3fb86baeda8a3b4c8;
wire [flogtanh_WDTH -1:0]        Ic66af6c3c0268cfb0e9f0776c4f4e961;
wire [flogtanh_WDTH -1:0]        I1ae4334c32094064c19df0dac77bd03d;
wire [flogtanh_WDTH -1:0]        Ia605d14205926b3edc6d1c2f69f70ac0;
wire [flogtanh_WDTH -1:0]        I78788f7e0845e4353145012efa04a48c;
wire [flogtanh_WDTH -1:0]        I0071f2168787bd42ab7f2370aed9d0f5;
wire [flogtanh_WDTH -1:0]        I359f3e3bb2a69349f8564466fa81a054;
wire [flogtanh_WDTH -1:0]        I4936f823841b0ffe32f801f5134c0211;
wire [flogtanh_WDTH -1:0]        I7b630e8ac26638fb858dd3b5d2d56385;
wire [flogtanh_WDTH -1:0]        I5975ef8f6cf53cf2132cdd9d707e7912;
wire [flogtanh_WDTH -1:0]        I859bef71501c2f2a994a0cdf8a94b2a7;
wire [flogtanh_WDTH -1:0]        I954ff0f9ee871a31774a3d786128fa13;
wire [flogtanh_WDTH -1:0]        Ib51b9e41161f4273f6469e8965acd7dd;
wire [flogtanh_WDTH -1:0]        I31f6bbfbbbd4c20d0c5c71663da1d4c1;
wire [flogtanh_WDTH -1:0]        I78bb23c008613c0f07f6f85172482296;
wire [flogtanh_WDTH -1:0]        I1898bc3cc6a8b6f71d65c758d1f08366;
wire [flogtanh_WDTH -1:0]        I8b883a5bc22b2cde03f4074357be7c88;
wire [flogtanh_WDTH -1:0]        If86532f849bd392dbf599eeb2fae0545;
wire [flogtanh_WDTH -1:0]        Ic2727e097ffbce70f07fc9f3d9395b54;
wire [flogtanh_WDTH -1:0]        Ia344734d285ac29b53cf401c08a0f987;
wire [flogtanh_WDTH -1:0]        I096397439036b0056c979054528ce1fd;
wire [flogtanh_WDTH -1:0]        I502a8e382aa0881dc86f3c13e0566ca3;
wire [flogtanh_WDTH -1:0]        Ifcc83d9007aafdf32acf04f062e008c8;
wire [flogtanh_WDTH -1:0]        Ic462cebbfc39190b22d20013259e39eb;
wire [flogtanh_WDTH -1:0]        I53c01c60f4061d970e4491564ddf88ae;
wire [flogtanh_WDTH -1:0]        I385d03def4cfb49f54867687ebd710ed;
wire [flogtanh_WDTH -1:0]        I0b4d34aa164c014f9315debd37fa534b;
wire [flogtanh_WDTH -1:0]        If8aa3ec1b5a4a3c122da82467be917da;
wire [flogtanh_WDTH -1:0]        Iac97aad4ca2c93e387ff0c1340143029;
wire [flogtanh_WDTH -1:0]        I8daf79a0a2ee1bac7f055af441539fa4;
wire [flogtanh_WDTH -1:0]        I8b4c2d8a5f2b796029575ecf3b89e2b9;
wire [flogtanh_WDTH -1:0]        I6261e0d339762cb2364421e6b87086cb;
wire [flogtanh_WDTH -1:0]        I06dd747316fa36a8dbdbb4ddf011230b;
wire [flogtanh_WDTH -1:0]        I0e2f746715b901feb69f6b3c94f3a828;
wire [flogtanh_WDTH -1:0]        I1594e7dfaedd9e7f5818dc4d639bb663;
wire [flogtanh_WDTH -1:0]        I7b8da162c08f8aa2ae90522ee1526cf6;
wire [flogtanh_WDTH -1:0]        Ic8111eb95e6b6ab35bcd8e2cafcd0c1e;
wire [flogtanh_WDTH -1:0]        I5e8ecdbb018402b2fbc0049ee44bae8c;
wire [flogtanh_WDTH -1:0]        I650b4641d233096a77ae15c8254a29b1;
wire [flogtanh_WDTH -1:0]        I06d859184884c07a14c83d2f06587ad5;
wire [flogtanh_WDTH -1:0]        Ia905d37c471bdf7258a547be95b85e4f;
wire [flogtanh_WDTH -1:0]        I79e3e49f57d47231c0fe6aaafdbc57f1;
wire [flogtanh_WDTH -1:0]        Icfc2b5de1aa36d81de3f163880d48a68;
wire [flogtanh_WDTH -1:0]        I12c07042202f66db926861c9ce7c2b25;
wire [flogtanh_WDTH -1:0]        I3c6893d360627cd954db1c20f3c9d319;
wire [flogtanh_WDTH -1:0]        I9d0fdb45b9e86bd409740e538a690320;
wire [flogtanh_WDTH -1:0]        Ibc971e0b7ade69365d2c23f30ba0c1ea;
wire [flogtanh_WDTH -1:0]        Id5fd6f25dc3df22a322434ae3c90dea6;
wire [flogtanh_WDTH -1:0]        I562d9a1676d27c7966d2920bb6be3b38;
wire [flogtanh_WDTH -1:0]        Id812a8ea2a3b4a912d151be582833fcf;
wire [flogtanh_WDTH -1:0]        I8aa258f382bea1eb300b006c3083bec1;
wire [flogtanh_WDTH -1:0]        Ifd3638d44e1ba2285891fac152dee327;
wire [flogtanh_WDTH -1:0]        Iec0e7232ec94c15d7d50866ad5eb85fb;
wire [flogtanh_WDTH -1:0]        Idd1b6014de2f053554ed09c29bf3e640;
wire [flogtanh_WDTH -1:0]        I0d252b23e06d25aee4afd84b4c5b4ba9;
wire [flogtanh_WDTH -1:0]        I0d96336eb4d5071d7e1d350e86513b25;
wire [flogtanh_WDTH -1:0]        I430703cef7ec173f9099c8391132e5c4;
wire [flogtanh_WDTH -1:0]        I31e5b2cdc3dc571eafa37510076bcc64;
wire [flogtanh_WDTH -1:0]        I5788d966ba8393f5d76dcfcb9294b52e;
wire [flogtanh_WDTH -1:0]        Ia8849f78971a45ed0daa2489e7d27dd7;
wire [flogtanh_WDTH -1:0]        Ied561890134d28b451f26da773ea5525;
wire [flogtanh_WDTH -1:0]        Ie4749f8e9ad2b370f9f9814b5a463c43;
wire [flogtanh_WDTH -1:0]        I52e018ad790a1e406777510a0f4b6c29;
wire [flogtanh_WDTH -1:0]        I3096d11098113da669ee0a94686e600d;
wire [flogtanh_WDTH -1:0]        I25eb66d8589cbb35b32cd25539a24f7f;
wire [flogtanh_WDTH -1:0]        I09a1d04c307fcb8a0e30925d86df3fe9;
wire [flogtanh_WDTH -1:0]        Icd4716d0d66d95a532544461c4872d11;
wire [flogtanh_WDTH -1:0]        Idb0a98cea3ee6cd4308bfc2414a003e1;
wire [flogtanh_WDTH -1:0]        I266ba4229056534d310d982253b5f9b9;
wire [flogtanh_WDTH -1:0]        Id4788855f9a503e8b506d012aaeea445;
wire [flogtanh_WDTH -1:0]        I86498c8c820d276ac12764b5df267252;
wire [flogtanh_WDTH -1:0]        I5b937934e7aae1f916c2848889f12685;
wire [flogtanh_WDTH -1:0]        I7bb9ad1a2cd32966746b05b7604a09b6;
wire [flogtanh_WDTH -1:0]        I9275bb36e58e0f17964e13ee7f027ab7;
wire [flogtanh_WDTH -1:0]        Id0998cc2848a6a72ed2701a8e720946e;
wire [flogtanh_WDTH -1:0]        I02330ade2eed926076cc071e45eed82c;
wire [flogtanh_WDTH -1:0]        If1ed051cd94d42e7836f82c10538b302;
wire [flogtanh_WDTH -1:0]        I296bc392d4223cbdd6f77be6523df819;
wire [flogtanh_WDTH -1:0]        I780afd116929565d1ff9b3833ba242d5;
wire [flogtanh_WDTH -1:0]        I31b0f2fe98cfddbc05dbd14be8be394b;
wire [flogtanh_WDTH -1:0]        I89ee99e699676bcec20031b6cad0e2ac;
wire [flogtanh_WDTH -1:0]        Ia71663e8f563041c27cd21a0c9c27a28;
wire [flogtanh_WDTH -1:0]        I862b467403c045e4694fb57d59e10064;
wire [flogtanh_WDTH -1:0]        Ib46b13498ec14ceaa56719f26f18febb;
wire [flogtanh_WDTH -1:0]        Ic3b554c66f652f027159dbc0fccc5ba3;
wire [flogtanh_WDTH -1:0]        I9bc2d5692474b8368c570d92835191b3;
wire [flogtanh_WDTH -1:0]        I04635713f6d70142b7ab3ecb5ffe6ac9;
wire [flogtanh_WDTH -1:0]        If8b0b96a659183e3651c691a2848b86b;
wire [flogtanh_WDTH -1:0]        I1917eae0dbcc0a941718c3248c7d4b11;
wire [flogtanh_WDTH -1:0]        I87d958c00fc6209d901147831b0c951c;
wire [flogtanh_WDTH -1:0]        Ifa60c3079164485f31442d9cf12bd2ad;
wire [flogtanh_WDTH -1:0]        Ie4e4eaf3e5d2f581210af8054df71c6c;
wire [flogtanh_WDTH -1:0]        I5616405acf49c3e8608ae4d2b544b0d6;
wire [flogtanh_WDTH -1:0]        I0b557cf102da41afd26936cbdb64b6e8;
wire [flogtanh_WDTH -1:0]        Ie6f9ae463fa1add4de23463435a23d25;
wire [flogtanh_WDTH -1:0]        I49eb064043f91112c854e31e4eb9b885;
wire [flogtanh_WDTH -1:0]        Ib16a67d67a4650e53547312e3af60363;
wire [flogtanh_WDTH -1:0]        I1039bc43e88eee527d2ed6adb8c7d1ba;
wire [flogtanh_WDTH -1:0]        I8fa4ad645ca2ef21dea8669d2e2afbe2;
wire [flogtanh_WDTH -1:0]        I9aab16e89f1b64117caece8ca8af5940;
wire [flogtanh_WDTH -1:0]        I41ea2e3d798ff8e0a95f04e4773c59b4;
wire [flogtanh_WDTH -1:0]        I343df614f97cf732e57cf2ad3f95dc9e;
wire [flogtanh_WDTH -1:0]        Id7f4c6208197cdbf48fecdb2a18b81fc;
wire [flogtanh_WDTH -1:0]        Ie02de90d8eb06b16314946d21299500c;
wire [flogtanh_WDTH -1:0]        I0adb66417482782dd71da1678c1f7412;
wire [flogtanh_WDTH -1:0]        I3353a7916b569f2c0ca122180608dccc;
wire [flogtanh_WDTH -1:0]        I2abe89a1366a1ad862266ad88101baa2;
wire [flogtanh_WDTH -1:0]        Ibfe760474fcac99f1e5ffa2e008fef99;
wire [flogtanh_WDTH -1:0]        I8d10f0c6dc026005f7882ca013283099;
wire [flogtanh_WDTH -1:0]        I3caf1211dcbcdc746a3e4c7fbbdae4a8;
wire [flogtanh_WDTH -1:0]        I4ef16908ce9b89771f94068eec1a983e;
wire [flogtanh_WDTH -1:0]        I2dcc0d17b9fcac35693bf32b5c5540fd;
wire [flogtanh_WDTH -1:0]        I4f6bcd6e0bcd77730248b69d2b93c904;
wire [flogtanh_WDTH -1:0]        Ie6764a631310e312ba5c2c1e601d828f;
wire [flogtanh_WDTH -1:0]        Iea1ae39e18f083fb8f855fd9ad3d4f8e;
wire [flogtanh_WDTH -1:0]        I220f8e45e5fe6e69f02cded87f12e1e5;
wire [flogtanh_WDTH -1:0]        I795ae30dec63ef2952917eb3355148a2;
wire [flogtanh_WDTH -1:0]        I896cd566a3d078b0f697a788efd223f2;
wire [flogtanh_WDTH -1:0]        I188813c5474bf304b59dbe07c78bef6f;
wire [flogtanh_WDTH -1:0]        I7caa41076a293edf18c7c4309fdcfc91;
wire [flogtanh_WDTH -1:0]        I1760a42d85513ea751e94a8b829b5f1a;
wire [flogtanh_WDTH -1:0]        I928a0e4951208aab170656596f456209;
wire [flogtanh_WDTH -1:0]        I8c652055cfcd230426887e171eaf2511;
wire [flogtanh_WDTH -1:0]        Ia3d129fd297905bee180293c0c39d9ef;
wire [flogtanh_WDTH -1:0]        I9a88a91b0fcc6dd1a7b4ed24e676d9e1;
wire [flogtanh_WDTH -1:0]        Id555c88cf7f0904db74d45cc75c8f5d6;
wire [flogtanh_WDTH -1:0]        I89f6566e2295d58668e63b9529d94df8;
wire [flogtanh_WDTH -1:0]        I1ddfd31bbf062aa5c3c71d61e492e3a2;
wire [flogtanh_WDTH -1:0]        I08295c218fd06a8900974edc9c2924f2;
wire [flogtanh_WDTH -1:0]        Iae9e023628eb6686708b2656f15616cc;
wire [flogtanh_WDTH -1:0]        I0a39fdea8b5bfac1862f199152e26ffe;
wire [flogtanh_WDTH -1:0]        If4b100d26126e460c41b8c1bc8fbbb96;
wire [flogtanh_WDTH -1:0]        Ib36a71ff310882325be0a2745e48f708;
wire [flogtanh_WDTH -1:0]        I85a7fede715578be0634d71e9c7951cd;
wire [flogtanh_WDTH -1:0]        I75e4d037cc2ed0b0f75fc1fe9cb21da3;
wire [flogtanh_WDTH -1:0]        I2d7715a3af03d9664729fa6df85034a2;
wire [flogtanh_WDTH -1:0]        Iee9e9849924642a9579a10655624fa17;
wire [flogtanh_WDTH -1:0]        I571ddcb0a10938e4c0816c965214b4a8;
wire [flogtanh_WDTH -1:0]        I0a267feb8313c9fa5c663a3fe68284dd;
wire [flogtanh_WDTH -1:0]        I8bf8b0cf27a2654a0e7fdf3255945b67;
wire [flogtanh_WDTH -1:0]        I0e0ff3511e65a1dda10ec944c89d09d7;
wire [flogtanh_WDTH -1:0]        I63f82f075d53205b5b556c0054f1a0b8;
wire [flogtanh_WDTH -1:0]        I4504a0a17633d26163a0afae21ad0f43;
wire [flogtanh_WDTH -1:0]        I3c6fb0df5846a19228a4e6cf9f9106ac;
wire [flogtanh_WDTH -1:0]        Ibd7b7f4ba86b6c61a0dd38f71c67ae05;
wire [flogtanh_WDTH -1:0]        I7168b0efdd2fae57292379c9d15c62eb;
wire [flogtanh_WDTH -1:0]        Icddd184270ffda26b803956883400ad0;
wire [flogtanh_WDTH -1:0]        Ibe502ebbb366f54a8f8fda4e361308e3;
wire [flogtanh_WDTH -1:0]        Id3da7061c05091ffc520d4480058e8e9;
wire [flogtanh_WDTH -1:0]        Ifce70fefde8f5ea4d2c1857236f66d65;
wire [flogtanh_WDTH -1:0]        Ie63d649228270b34d8ed25e7c4b09883;
wire [flogtanh_WDTH -1:0]        Ice2c390d296e09b117d60905343e9098;
wire [flogtanh_WDTH -1:0]        I8eed3f7b36c046fff1e41dd52a300d29;
wire [flogtanh_WDTH -1:0]        I4b94402a53d981e953c21ef316c709b7;
wire [flogtanh_WDTH -1:0]        Iefcebe38e0c2d6d570017e165d70d3b1;
wire [flogtanh_WDTH -1:0]        I450c0d6ad5d3b1f18bb28e3a432b5442;
wire [flogtanh_WDTH -1:0]        Ia153222350357443978d7426663c3eaa;
wire [flogtanh_WDTH -1:0]        I2587a5800a5a9ffeabc4dca503e3d964;
wire [flogtanh_WDTH -1:0]        I06f0fd2d9d46a2fdb4221217ee2496d1;
wire [flogtanh_WDTH -1:0]        I1182655739d7ab5bbe4a6546a5ca36fd;
wire [flogtanh_WDTH -1:0]        I9533ff0882ed01409795d7269329fd76;
wire [flogtanh_WDTH -1:0]        I8110a5a62607093b21b7cd088b1d9ee0;
wire [flogtanh_WDTH -1:0]        Ia9eb9821e7dc31c23d7e60839949c1ff;
wire [flogtanh_WDTH -1:0]        I8b611f7c12ddd81de403ba74e212857f;
wire [flogtanh_WDTH -1:0]        I3663fc86620d6244a850819bd3ebe72c;
wire [flogtanh_WDTH -1:0]        I84a62a133dbceb5a32a7c907f371663d;
wire [flogtanh_WDTH -1:0]        I11293e7cdeddf352011d46abd6c3bb72;
wire [flogtanh_WDTH -1:0]        Ia2fc8a1bbc3cb0dd7d89a7f05b04909c;
wire [flogtanh_WDTH -1:0]        Ic9339e415d0f756e34bcd930de63ad87;
wire [flogtanh_WDTH -1:0]        I2a3eb42a4402e873d081f94a14a99c20;
wire [flogtanh_WDTH -1:0]        Icf109f65e24d3a23ecad9e7d4cc54dc1;
wire [flogtanh_WDTH -1:0]        I58447d6ae49a6be2d043477a06f83df0;
wire [flogtanh_WDTH -1:0]        Idf7dd0ff83b2d56693e729a1a375fabb;
wire [flogtanh_WDTH -1:0]        I83292bcda4645233d8e8a1dfe8e5f60b;
wire [flogtanh_WDTH -1:0]        I312a248019372261c0959cdc9378ec93;
wire [flogtanh_WDTH -1:0]        Ic5e0a84cf1a2ef907b2456559ea26c75;
wire [flogtanh_WDTH -1:0]        I8e311b9891dda272762da2c640019e8c;
wire [flogtanh_WDTH -1:0]        I2cefbf897bb7f6f67ca500727e85c683;
wire [flogtanh_WDTH -1:0]        I1874dd9f7c0a93310873173561402912;
wire [flogtanh_WDTH -1:0]        If47be2ca4617a426258c51f8d977ba3f;
wire [flogtanh_WDTH -1:0]        I04adb3964e739a106098a6c4d2f49e94;
wire [flogtanh_WDTH -1:0]        I7c68e0ae30efc4ca4d68b6047119c6c3;
wire [flogtanh_WDTH -1:0]        I9135b709c3c802a42c7186087b5664cc;
wire [flogtanh_WDTH -1:0]        Iccca1936f4c1c9496205e77b588e9985;
wire [flogtanh_WDTH -1:0]        Ia236dfe34ff4938456d76f787d2db945;
wire [flogtanh_WDTH -1:0]        I59d4567d3355fdae5660a1364d1b8d00;
wire [flogtanh_WDTH -1:0]        I41c98bae5fbdb31bac0913930573e80c;
wire [flogtanh_WDTH -1:0]        I4600963866dcb9bbea2515c805f885cb;
wire [flogtanh_WDTH -1:0]        I226befd72285893998aca87fe34d9aaf;
wire [flogtanh_WDTH -1:0]        If26d90629e70c5a871e6f5b14471b8cf;
wire [flogtanh_WDTH -1:0]        I20ab7c6174af39aee99492f704b2748c;
wire [flogtanh_WDTH -1:0]        Iedb9bb14951bf67bc8865b0983490c14;
wire [flogtanh_WDTH -1:0]        I0a1c5724ffa14df653142a1f8bcf44a4;
wire [flogtanh_WDTH -1:0]        I6a3854ed571e8c262aa3ec377c247778;
wire [flogtanh_WDTH -1:0]        I481973954b81accf069dd80830fba3bc;
wire [flogtanh_WDTH -1:0]        I05028975b49ec0c089bd981696f85a8b;
wire [flogtanh_WDTH -1:0]        Ia6825c3edc9d2a6832db7a7d684faf98;
wire [flogtanh_WDTH -1:0]        Ife732309efcc740cfff5c747aab2e3d6;
wire [flogtanh_WDTH -1:0]        I5c964036207f47629302e282d56fef7b;
wire [flogtanh_WDTH -1:0]        Idcef10a0465614cf38e0d6f503b5174a;
wire [flogtanh_WDTH -1:0]        I00b74ed4d6730b37c6fbfd42dee42584;
wire [flogtanh_WDTH -1:0]        Ibd4aaf02982068ffbfd1b8b3795d9217;
wire [flogtanh_WDTH -1:0]        I0345fc4a507f9e3be3e1d46b71693de1;
wire [flogtanh_WDTH -1:0]        I788c64785b992c675fe348a1fa181525;
wire [flogtanh_WDTH -1:0]        I9f0735c1cf5d1af7c82a251ef4886f9c;
wire [flogtanh_WDTH -1:0]        Ib235af5b28d56f24372d3f0af816f2c2;
wire [flogtanh_WDTH -1:0]        I861cf5dffb18c84953013dc4026bd08a;
wire [flogtanh_WDTH -1:0]        I4c03a6569d1b954d088053e38827e811;
wire [flogtanh_WDTH -1:0]        I19722ceada71cc9cc06edde39142ff17;
wire [flogtanh_WDTH -1:0]        Idda26504e422367082caeafbb29871f9;
wire [flogtanh_WDTH -1:0]        Id8349128e2c391df008828494da928c6;
wire [flogtanh_WDTH -1:0]        I195c3a82123142d509886ee37dc6fc98;
wire [flogtanh_WDTH -1:0]        I27209805df490a07f1726875a7b69922;
wire [flogtanh_WDTH -1:0]        I1abb512ca0383c9e7104418e07281841;
wire [flogtanh_WDTH -1:0]        I7532c1f0624a2d5a94321c89c73e38df;
wire [flogtanh_WDTH -1:0]        I00ff1331b1900bb031ee81d2a58c1bd5;
wire [flogtanh_WDTH -1:0]        Ife892846e66e2522c06b170811a11ada;
wire [flogtanh_WDTH -1:0]        If65eb5e743a7b1878fb232ef2fe13cb0;
wire [flogtanh_WDTH -1:0]        Ib905ede2830f7e3c8cf993075f07345c;
wire [flogtanh_WDTH -1:0]        I24ae7de3549a84f4f88f561b6017b7a8;
wire [flogtanh_WDTH -1:0]        Ibf169f844d9e00eca8f3821ddc952ef0;
wire [flogtanh_WDTH -1:0]        I449c77140475475b138d839a74078337;
wire [flogtanh_WDTH -1:0]        I3137f75629e72f78abdac088e18608d5;
wire [flogtanh_WDTH -1:0]        Ia9e102d8679943c079f16c0228f0f0d1;
wire [flogtanh_WDTH -1:0]        I8fbcabc2f5c30fcf1c5b46de5dfe887d;
wire [flogtanh_WDTH -1:0]        Ibf1c9d86665f696d91c554db748ff42b;
wire [flogtanh_WDTH -1:0]        Ie7acfb624aa6242b558481350c85fda3;
wire [flogtanh_WDTH -1:0]        Ieb0336a1974a2aec0966f4f59f460802;
wire [flogtanh_WDTH -1:0]        I11e0b915338d5d649c800455b9a7695f;
wire [flogtanh_WDTH -1:0]        Ic0819ccefe784a6379716b3633ae0196;
wire [flogtanh_WDTH -1:0]        Ia9e4e68dcd3d0281decde939eed0c3bd;
wire [flogtanh_WDTH -1:0]        I0c4bbd1827b1859caabb067e864ce4b3;
wire [flogtanh_WDTH -1:0]        Id508f63a381fc565a28fe4e662b33efb;
wire [flogtanh_WDTH -1:0]        I004c98da87996b77b5761d366210f782;
wire [flogtanh_WDTH -1:0]        I33582dc83370e68b0ae7b22b553276b4;
wire [flogtanh_WDTH -1:0]        Ia457938da4efe847cb06f645f2a54a52;
wire [flogtanh_WDTH -1:0]        I8aeca996ad6820edcc6fcbaa8a0f15ce;
wire [flogtanh_WDTH -1:0]        I7e0474089ebc1c34747be1bc17a81d72;
wire [flogtanh_WDTH -1:0]        Ica86e8037319b868c8cb89f3cb02b136;
wire [flogtanh_WDTH -1:0]        Ib0b46b99e61d724ae664d9d1fec1e29f;
wire [flogtanh_WDTH -1:0]        Ia95013b19d9fc12d19ff9924007113d4;
wire [flogtanh_WDTH -1:0]        I56d1025271f1f7704a40dd7f0df02b0b;
wire [flogtanh_WDTH -1:0]        Ifcf979b713b014f22c1c8ce1d42132c2;
wire [flogtanh_WDTH -1:0]        I72c2256ba47cf03f95143df8f741fd83;
wire [flogtanh_WDTH -1:0]        I973b3306021532f286cf248084398c26;
wire [flogtanh_WDTH -1:0]        I733c3fa4d84e5680792b16a70bb1a51d;
wire [flogtanh_WDTH -1:0]        Iea7940bb396d1a436f56806fc533edee;
wire [flogtanh_WDTH -1:0]        If367d63311c96726517240de13bd2a4b;
wire [flogtanh_WDTH -1:0]        Ied55045b003302c294591a8d2a6a39fd;
wire [flogtanh_WDTH -1:0]        Icc6d895d943e14f2801c22e79ce190e8;
wire [flogtanh_WDTH -1:0]        Ib64e948413d5dce1d9309fe95c0919ab;
wire [flogtanh_WDTH -1:0]        Ieb664ac9be65fba2e25960141f7fb4b6;
wire [flogtanh_WDTH -1:0]        I682fe6c6c621db5dd867574e8573d8ed;
wire [flogtanh_WDTH -1:0]        I66071f20991b414140869a2e3b750471;
wire [flogtanh_WDTH -1:0]        I508b57f6ebc45eb70aa7b114096a7d12;
wire [flogtanh_WDTH -1:0]        Iffeefa89a2ba7d032db5db64cbf05e20;
wire [flogtanh_WDTH -1:0]        I8e82b8914260669ed1d88a690467a7b4;
wire [flogtanh_WDTH -1:0]        I9ab3cea6ee8d8473221da21bae06066b;
wire [flogtanh_WDTH -1:0]        I525feb94b558fb4bb8db8eead9f05afa;
wire [flogtanh_WDTH -1:0]        I3403ce6e697b523a9f441d8fd5e2d420;
wire [flogtanh_WDTH -1:0]        Ie5e4cf2b42054822a9091f5ef67cd968;
wire [flogtanh_WDTH -1:0]        Ia98a70144e466b356d2998948dc4b602;
wire [flogtanh_WDTH -1:0]        I0d08d26e31c8b69ed8c089cdcd055a50;
wire [flogtanh_WDTH -1:0]        Ie4ca0836695d951ee09622892ee35928;
wire [flogtanh_WDTH -1:0]        I877f44c880a781381bfa8a8f8471d697;
wire [flogtanh_WDTH -1:0]        I485a48b4ff4da08f977425fd10e6d392;
wire [flogtanh_WDTH -1:0]        I7fc78273dc765cf1c03b3c1a043b35f8;
wire [flogtanh_WDTH -1:0]        Ie8c79e6a5378808c0ead5a4b24319ce9;
wire [flogtanh_WDTH -1:0]        Ie67275a4b3fdc050f0f6e7ac7d1eebfc;
wire [flogtanh_WDTH -1:0]        I9ca81c841a75a9ac242835956509e0fe;
wire [flogtanh_WDTH -1:0]        I41f9acc96650353174155a5f378d5cc5;
wire [flogtanh_WDTH -1:0]        Id50f18f642f3b00ffa34986f78a0eae6;
wire [flogtanh_WDTH -1:0]        I0d73c905b2ed777acd71d560928dcf0b;
wire [flogtanh_WDTH -1:0]        I75838ca09e301b8e1301cbf603a1f8c2;
wire [flogtanh_WDTH -1:0]        I2b6b1c25caf8b00d19ccc98156a8ca2b;
wire [flogtanh_WDTH -1:0]        Id968b34075e351ab01d65abcb4ed8cca;
wire [flogtanh_WDTH -1:0]        I28ea2b207bcd3518a85ff150466a6a08;
wire [flogtanh_WDTH -1:0]        I84da4ce7441e132e775167c1cd81dbe5;
wire [flogtanh_WDTH -1:0]        I7d0a1c64b2e85e1bf0bf99423321466b;
wire [flogtanh_WDTH -1:0]        If19dc22d45cc4664c85a043ec4c00617;
wire [flogtanh_WDTH -1:0]        I3b9b9b41b54ff194314b572a15daf606;
wire [flogtanh_WDTH -1:0]        Ibf482db0f5058be72061267c42ebc292;
wire [flogtanh_WDTH -1:0]        Ic914f847e623d9c52e2d9ae5076c21c3;
wire [flogtanh_WDTH -1:0]        I6d2dbb953a58b91dafa7f0d34d41bdc3;
wire [flogtanh_WDTH -1:0]        I46fc20938dd554b23b5af5f7c3e39480;
wire [flogtanh_WDTH -1:0]        Ib393146d81d3cf031466543311cee2ad;
wire [flogtanh_WDTH -1:0]        I1fa8b37b4697ae60cf399285d9524b8d;
wire [flogtanh_WDTH -1:0]        I42564ec6a794ea803795f0b5b3523a93;
wire [flogtanh_WDTH -1:0]        I66c8261df769288836e188ecb32b6dc6;
wire [flogtanh_WDTH -1:0]        I4a0033a180d7edce81fcfef603532e28;
wire [flogtanh_WDTH -1:0]        I267714c8a5aa14bae9c74da272a60aa5;
wire [flogtanh_WDTH -1:0]        Ic7a21921e2716fba55aad2e351f4498a;
wire [flogtanh_WDTH -1:0]        I47a34c8d2174c12f96041e82ad835db2;
wire [flogtanh_WDTH -1:0]        I9a3f0b4867087790c78f674b719dbf7b;
wire [flogtanh_WDTH -1:0]        If99ca487495a015063fd8dc54ae596aa;
wire [flogtanh_WDTH -1:0]        I138f008a6206a1067bb0e22ce3d90990;
wire [flogtanh_WDTH -1:0]        I1043f1b92b49a8c304a23c0b5c615def;
wire [flogtanh_WDTH -1:0]        I48ad9b737892d7c49340ed679f46e034;
wire [flogtanh_WDTH -1:0]        Icafa102383ef33455236ba268b1b7460;
wire [flogtanh_WDTH -1:0]        I04a9c9765fd468a7e841577f09fc287b;
wire [flogtanh_WDTH -1:0]        I677fca8017154fed3e6cd54362e829db;
wire [flogtanh_WDTH -1:0]        I7b929c228c865112f00bc6b4dcc95b52;
wire [flogtanh_WDTH -1:0]        I826fe051a6b09d5cacf712431ce89b7c;
wire [flogtanh_WDTH -1:0]        I2b54a135e59945901e9c11580a29ee3d;
wire [flogtanh_WDTH -1:0]        I23f781ebfa449cec7975b94179d72259;
wire [flogtanh_WDTH -1:0]        I566221060f06e724676ec9bec861d7de;
wire [flogtanh_WDTH -1:0]        Ia383b5dc3b7ce1bc7987926535639668;
wire [flogtanh_WDTH -1:0]        Icd9a876a0feb16ea62bcad5be2004dac;
wire [flogtanh_WDTH -1:0]        I40ae857caffae41564c2ecb0c7e9777b;
wire [flogtanh_WDTH -1:0]        I8f8273c4cb2a9ace8a09847efd4bdec7;
wire [flogtanh_WDTH -1:0]        I569d56a2673a104f3050d851d767af8a;
wire [flogtanh_WDTH -1:0]        I96ef4b631a7f63e19f67f3920685f0e6;
wire [flogtanh_WDTH -1:0]        I2022005072d2979dae84b6e4491a3ce2;
wire [flogtanh_WDTH -1:0]        I9e2de71442b8f504358e582087a6d19f;
wire [flogtanh_WDTH -1:0]        I98524ad028e4d832ebbcd92956dac08c;
wire [flogtanh_WDTH -1:0]        I1fb13d7500f5ac3821c424bd3688cf4e;
wire [flogtanh_WDTH -1:0]        I4d24e2ba47093eee6669f537374ecce7;
wire [flogtanh_WDTH -1:0]        I2aabda12ff89e708d04b4399472b5203;
wire [flogtanh_WDTH -1:0]        I227232e7189020459c16b3413e881b80;
wire [flogtanh_WDTH -1:0]        I8c733a5d394e6b8d045eede5cc7451f6;
wire [flogtanh_WDTH -1:0]        If4359aebd4cc66c75cf2a44f681ccc72;
wire [flogtanh_WDTH -1:0]        I4f45dd50d2825ab338b8a2a8264096c0;
wire [flogtanh_WDTH -1:0]        I8d2e10b8c474f1a915825ec78072ad56;
wire [flogtanh_WDTH -1:0]        Ib45caf6b563d22144be3e9225a99a1cd;
wire [flogtanh_WDTH -1:0]        Ie5b3748f3c81d9eeec767d546b29cbd8;
wire [flogtanh_WDTH -1:0]        I9d6730140c690037b5ca58aa30103f5b;
wire [flogtanh_WDTH -1:0]        Ib764a6d1978dc61cb4499b15c45cb1b4;
wire [flogtanh_WDTH -1:0]        I9df5b63f66c162d517daa69f5d0e6095;
wire [flogtanh_WDTH -1:0]        I4fbe7db2d4288676183dc69ed56c9c68;
wire [flogtanh_WDTH -1:0]        I1b40adfd6fa6c943dfa8d230d9e65514;
wire [flogtanh_WDTH -1:0]        I99f0cc5986099cb57fbebf9e5e262c56;
wire [flogtanh_WDTH -1:0]        I0eb3df4d4094e09e6c4b3c788baed61f;
wire [flogtanh_WDTH -1:0]        I4f5bb7e206563a334d7e2dd100b37c35;
wire [flogtanh_WDTH -1:0]        Id6f7923a16cc5adc96a730083153ca6d;
wire [flogtanh_WDTH -1:0]        I59ecb14b5f34ebab3da4784709de66a4;
wire [flogtanh_WDTH -1:0]        Idf8ebc0d747ae143aa61866e33d458c0;
wire [flogtanh_WDTH -1:0]        I54f5a8caf0e1c2df9477b37157d94995;
wire [flogtanh_WDTH -1:0]        Id682e531735437bc24abbf3d3d51e18b;
wire [flogtanh_WDTH -1:0]        I77e1bed2da0ccf1475dcfe908d64f82c;
wire [flogtanh_WDTH -1:0]        I05ecce409cca00ea5b0df25de5a50cf2;
wire [flogtanh_WDTH -1:0]        I1a450ec193ccde2946f6ca20c0fa894c;
wire [flogtanh_WDTH -1:0]        I831d214dcb4f8d534b5ddaaeaeeb81ce;
wire [flogtanh_WDTH -1:0]        I01fbfc3b5c14733738f93a3487e54f35;
wire [flogtanh_WDTH -1:0]        Ia540866403683bc30504bace19bdda7b;
wire [flogtanh_WDTH -1:0]        Icff5d12020f78478c77210d9c692dfbe;
wire [flogtanh_WDTH -1:0]        I05fb1982415bd3fa78dd9a00af7a3d4a;
wire [flogtanh_WDTH -1:0]        I6eb28698ab4105a74c6510dbcfefbc3c;
wire [flogtanh_WDTH -1:0]        I977864efb0d94149cce7dc4d165f11de;
wire [flogtanh_WDTH -1:0]        I7cc0f835ad7a18683e1fdb5bcbfb7f2f;
wire [flogtanh_WDTH -1:0]        I9362b615a612599239e3b752a9334e8c;
wire [flogtanh_WDTH -1:0]        I9389a0dfe5a82a903c89e1a468f0ad57;
wire [flogtanh_WDTH -1:0]        I5d4fb4b5a5ad3dc48beebfa0e0cebbed;
wire [flogtanh_WDTH -1:0]        Idc4ce4afd846e212526d21a5e0cd1c14;
wire [flogtanh_WDTH -1:0]        Ifb9b29c43f435452cc761218c509f5df;
wire [flogtanh_WDTH -1:0]        I38a0ba1e69b467d4aed306e76ec3bfdb;
wire [flogtanh_WDTH -1:0]        If2143db72bf9a02b64eb45b3a4faa39d;
wire [flogtanh_WDTH -1:0]        I66279b0fa707a272f43ee929cb297945;
wire [flogtanh_WDTH -1:0]        Ice780b1695a8e80607a03dee3c426ffe;
wire [flogtanh_WDTH -1:0]        Ib091954846c14743e01fd4e7bafda1b5;
wire [flogtanh_WDTH -1:0]        I90b0296f5ef87dfaa6110fc2e9d6ed9d;
wire [flogtanh_WDTH -1:0]        I3b8663f2adecb8da2c84dbb37341e25f;
wire [flogtanh_WDTH -1:0]        Icd37da8ea84a606529e32b2db4eb7f5f;
wire [flogtanh_WDTH -1:0]        I19bc03089c6c288e1778bd1f197a3ce3;
wire [flogtanh_WDTH -1:0]        Ie626a24e3680f7d3995dd0c2ce60cbcc;
wire [flogtanh_WDTH -1:0]        I0988382a446b21da209d49d0d00bd6df;
wire [flogtanh_WDTH -1:0]        Iebee55168fb47664095b11c9f6641124;
wire [flogtanh_WDTH -1:0]        I19f5cb50b27b6c5e40012df9397aa288;
wire [flogtanh_WDTH -1:0]        Ic0954671eb1dc893c3932e456800fadf;
wire [flogtanh_WDTH -1:0]        I706ca74386e5778b30eca35432429bc3;
wire [flogtanh_WDTH -1:0]        Ia4131464996aabab8aae1db85f6a50e4;
wire [flogtanh_WDTH -1:0]        If6af0cc7a120b2897c3a69d54a554e86;
wire [flogtanh_WDTH -1:0]        I2de1ca2c390bdd3011fff4a359bb5332;
wire [flogtanh_WDTH -1:0]        I88ebe846173f486b07d2051a80bd055f;
wire [flogtanh_WDTH -1:0]        I6fb55222b69475b7168874423226ec9c;
wire [flogtanh_WDTH -1:0]        I2c577b130db6f4673704c858d454f3ea;
wire [flogtanh_WDTH -1:0]        I9b09b800a9dcd8ac36f25cb0324e748d;
wire [flogtanh_WDTH -1:0]        I383f23d4e769bbdc1c8acd9c660a0b3e;
wire [flogtanh_WDTH -1:0]        I74ac0327175f50f508a5013df298df02;
wire [flogtanh_WDTH -1:0]        Iea20a6ecf4bbf907d1a102bde797284f;
wire [flogtanh_WDTH -1:0]        Ica26f542586d50c56ce0f3c00f36b388;
wire [flogtanh_WDTH -1:0]        I77d655383c0c22b1af75d9308fab2e4f;
wire [flogtanh_WDTH -1:0]        I7c6862830daffc98cb2c1fc121d82c38;
wire [flogtanh_WDTH -1:0]        I4a4ebb2f3389d67c4b7671e12fc5cd92;
wire [flogtanh_WDTH -1:0]        Icf19dd665616a8c96146b3ab9f46c741;
wire [flogtanh_WDTH -1:0]        Ibc927d678e218397e23147b5c0654fd9;
wire [flogtanh_WDTH -1:0]        I97f2813ec39bbf1513faf66b3e38838a;
wire [flogtanh_WDTH -1:0]        Ib0358b6f47edcd54971935de215203f8;
wire [flogtanh_WDTH -1:0]        I716ee53e79883f69aa045380a357e913;
wire [flogtanh_WDTH -1:0]        Iaa6f2bbd8a343ebf878da57badb4572b;
wire [flogtanh_WDTH -1:0]        I25c324feaca84e80f58075597e8c448f;
wire [flogtanh_WDTH -1:0]        I823f1a0d2d757d5ca83dc7b5ca08e0f8;
wire [flogtanh_WDTH -1:0]        I7fc190647082a3d71614f46f670167bc;
wire [flogtanh_WDTH -1:0]        I1a650234a61a3ff90ea079e29d322069;
wire [flogtanh_WDTH -1:0]        Iebdf938a28594624f4d4a337356485cb;
wire [flogtanh_WDTH -1:0]        I70a7b1083c9593840759854430ee9d62;
wire [flogtanh_WDTH -1:0]        I3fd068d55154441ffd005999ea823fd0;
wire [flogtanh_WDTH -1:0]        I99aa55a3e285e62e9a8b50174e84b68c;
wire [flogtanh_WDTH -1:0]        Ic5ca74b66763c6e5591c7c2bfeeb0663;
wire [flogtanh_WDTH -1:0]        Ief099d2084b84e0e23599d98102a13b7;
wire [flogtanh_WDTH -1:0]        I5ab556386d2973354a5551ba9823e4ba;
wire [flogtanh_WDTH -1:0]        I84aa89bab681c2fc7a8c7c6b47200dec;
wire [flogtanh_WDTH -1:0]        I64f65df774d29696425ba460dda09b68;
wire [flogtanh_WDTH -1:0]        I101b9397639b59fd53a88d17425e0c96;
wire [flogtanh_WDTH -1:0]        I9e09c25be9f877c1e1aaf79bf12c7943;
wire [flogtanh_WDTH -1:0]        Ic302f050dba883d8f4bd20b1030ba14d;
wire [flogtanh_WDTH -1:0]        I42c1d469ff97913cbf15e3ebee6fdfa8;
wire [flogtanh_WDTH -1:0]        I848425f041888d7433b68900f259732a;
wire [flogtanh_WDTH -1:0]        If9f2a53dbf6e9b9a335a7657b7a2b468;
wire [flogtanh_WDTH -1:0]        I2b4671193178503f5329954e74a399b3;
wire [flogtanh_WDTH -1:0]        I495f8be463b15db906474c518e0741e2;
wire [flogtanh_WDTH -1:0]        I97b93c6d963d51a819b1dc9ab3bf28ea;
wire [flogtanh_WDTH -1:0]        I3e265a7dcf29687248b9275df49771fb;
wire [flogtanh_WDTH -1:0]        I2593b1b30f4c97845a1f77c3f558b263;
wire [flogtanh_WDTH -1:0]        Iffd94cf3a8a4681ff3327c90bf89bd8b;
wire [flogtanh_WDTH -1:0]        I3a4695c79b62f6baa47cdc939c4e2974;
wire [flogtanh_WDTH -1:0]        Iea71417e738c6ca54c50aa014cc38627;
wire [flogtanh_WDTH -1:0]        Ibc577b2948aec87c0696c860d7efa1d7;
wire [flogtanh_WDTH -1:0]        Ic8df04756f67e6dd29f3374c5f86d451;
wire [flogtanh_WDTH -1:0]        I08401e4e9a1766a0034f45933b5bb29a;
wire [flogtanh_WDTH -1:0]        I546122346a22ad64a6ab2b4978cde095;
wire [flogtanh_WDTH -1:0]        I5e5bb0de4fe6682a6beaa86f6cd1ca32;
wire [flogtanh_WDTH -1:0]        Icaae0fb0f460f68d690ab00697355a49;
wire [flogtanh_WDTH -1:0]        Ia487e80f0010e7cb34aa12471e62a62f;
wire [flogtanh_WDTH -1:0]        I42455e7e4d0c63f97702d204d18a446e;
wire [flogtanh_WDTH -1:0]        I3bee9305e2f4456aae800bbb174b7843;
wire [flogtanh_WDTH -1:0]        Iaec2f15665e83416bc140890f3cdde9a;
wire [flogtanh_WDTH -1:0]        I14f1aa0dbf6f1f0fbf6b5f996e229a04;
wire [flogtanh_WDTH -1:0]        I487391402b6aa27bf212724a37ea9c33;
wire [flogtanh_WDTH -1:0]        If87afc1cf342dca9986f798c38a69dab;
wire [flogtanh_WDTH -1:0]        Ia9f375709014a9d553d46cff2799b59f;
wire [flogtanh_WDTH -1:0]        Ibb1c020ea255a966e54c00fc7cc745b5;
wire [flogtanh_WDTH -1:0]        I34d428a56bd0142a9be9f627f1c3c87f;
wire [flogtanh_WDTH -1:0]        Icae8a2980dd7403caf72820ae508885b;
wire [flogtanh_WDTH -1:0]        I57db98eb439d59a895dabe029c6a3a8b;
wire [flogtanh_WDTH -1:0]        Ic8f858d7f7a16b771933741d31679dc1;
wire [flogtanh_WDTH -1:0]        I9937af6fcf9d834f308bc3683d524981;
wire [flogtanh_WDTH -1:0]        I9dcf19da38f352fe7fa27c22bff08c19;
wire [flogtanh_WDTH -1:0]        I463f4f370e1ecad71de44780eff10df4;
wire [flogtanh_WDTH -1:0]        I2bc787aa749db4a5f48bd917715a11d5;
wire [flogtanh_WDTH -1:0]        I53309409a6059c3bd39f037c23ec3458;
wire [flogtanh_WDTH -1:0]        I3d072e173fd12ac9d802a29a0ff4378c;
wire [flogtanh_WDTH -1:0]        I2603e0b8b93f6680e44c9c8883f6512c;
wire [flogtanh_WDTH -1:0]        I2115d62275a57ec7273e3631c0a32872;
wire [flogtanh_WDTH -1:0]        Iab354cc9ac1173335c0efeef694f3567;
wire [flogtanh_WDTH -1:0]        I91bc663fcd7f86a066b8b3f93b1dcfc2;
wire [flogtanh_WDTH -1:0]        I6c19936ca2edeb0e261e880a1055e964;
wire [flogtanh_WDTH -1:0]        I988c0d94f97329dd1cff7d913cb449e7;
wire [flogtanh_WDTH -1:0]        Ifebfa58419ecd22a334ed4b67f5c3581;
wire [flogtanh_WDTH -1:0]        If444a37a85774dcc2769ffd74b785e46;
wire [flogtanh_WDTH -1:0]        I71a28e8525f07dabeabe4b4f45f353d0;
wire [flogtanh_WDTH -1:0]        Idbb89639b8399b57b190efd898643328;
wire [flogtanh_WDTH -1:0]        I514830acdad20c4ff3d078477e939b4b;
wire [flogtanh_WDTH -1:0]        Ib1d70f302858eb7c78fb834071616a9b;
wire [flogtanh_WDTH -1:0]        I036342f6be0f2e2f1f4927099a5c4a78;
wire [flogtanh_WDTH -1:0]        I82bd4ea32da7ae3a0d5938fc8a1424c5;
wire [flogtanh_WDTH -1:0]        Iedb655aa25e5f0e35137ec6c3acdc527;
wire [flogtanh_WDTH -1:0]        I6964f2e681e9cdf63fbc0358cb6edcca;
wire [flogtanh_WDTH -1:0]        I0c59e8c82a31aacbf5977ff778a7ff49;
wire [flogtanh_WDTH -1:0]        I41aeb75239ce0d636288e8ceb0665b34;
wire [flogtanh_WDTH -1:0]        I1b6d20c64b9f23fb6c30f723546aa285;
wire [flogtanh_WDTH -1:0]        Ie0d3fd5e7c38c10fdcae3f1b217c28f4;
wire [flogtanh_WDTH -1:0]        I0d66aa55747362354aa81d96057bc4c2;
wire [flogtanh_WDTH -1:0]        Ia8b7d74eaf227e697c3eb58b31eb355f;
wire [flogtanh_WDTH -1:0]        I1ea33707e40a2e41513fdb3118371437;
wire [flogtanh_WDTH -1:0]        I79034cd4180d03348de2c101927048a7;
wire [flogtanh_WDTH -1:0]        I68c85727adecde0aa8aa66ed08c4b502;
wire [flogtanh_WDTH -1:0]        Id23895e0696cdd27e3087294fb52a65b;
wire [flogtanh_WDTH -1:0]        Iebd050e29044153d5881ef80b2db8c28;
wire [flogtanh_WDTH -1:0]        I43939a168f9f5e476262ace39c6ae483;
wire [flogtanh_WDTH -1:0]        I3c057d64cf4fca0238a874f0ced99c76;
wire [flogtanh_WDTH -1:0]        Ie5167faac3e6510d4b208a1bdc0cd44c;
wire [flogtanh_WDTH -1:0]        I066cd52173ec5dbce9a3f470d73325af;
wire [flogtanh_WDTH -1:0]        I1cad8b885a541dd049093ce60c3f8a06;
wire [flogtanh_WDTH -1:0]        Ic7ad59f6a232a997706d17b4098e0324;
wire [flogtanh_WDTH -1:0]        Icd2d69f12d4744ce7b09fce7f27ab830;
wire [flogtanh_WDTH -1:0]        Icf8cfc800f0a2aa5140a7f83f035b0cc;
wire [flogtanh_WDTH -1:0]        Ic9ee0243e36f66f462eb3d4ce93fdde9;
wire [flogtanh_WDTH -1:0]        I6bfbf7ff79ff0a6facc9ba5031239644;
wire [flogtanh_WDTH -1:0]        I5353c3239ddb4d7fa7094e413b5303b1;
wire [flogtanh_WDTH -1:0]        I78ade92efd265027807c861be44a10af;
wire [flogtanh_WDTH -1:0]        Idfca1b1d8041e5808799499e8c8dcf5e;
wire [flogtanh_WDTH -1:0]        I2bc5a10c587d89d10021aa5eaafb490a;
wire [flogtanh_WDTH -1:0]        I4710d61c763098027934286c6a9f3714;
wire [flogtanh_WDTH -1:0]        I30080cc6c03bbe933165d266558a822c;
wire [flogtanh_WDTH -1:0]        If6a04c29b7205c5db5f2ff3cf302c45f;
wire [flogtanh_WDTH -1:0]        I7e28234bdf66ab5489d36d15678db797;
wire [flogtanh_WDTH -1:0]        Ib5d9348a114627a8b1f56aca968d20b1;
wire [flogtanh_WDTH -1:0]        I74b3c9dd3a8168aacd4369b9ff68fdfd;
wire [flogtanh_WDTH -1:0]        I4e2b59a03731959106d469ffee7b7d33;
wire [flogtanh_WDTH -1:0]        Ia7046faae1ab05978e4b32bd44049fb9;
wire [flogtanh_WDTH -1:0]        Ic6d519691c7543b1bd0707a8c9899088;
wire [flogtanh_WDTH -1:0]        I0c5250aaca86185fed5978438c8861b6;
wire [flogtanh_WDTH -1:0]        Icc6bde490bd8df2ce5efe8cfb24cf5f5;
wire [flogtanh_WDTH -1:0]        Ic78949e07e643f571f23df7e8f15d9fb;
wire [flogtanh_WDTH -1:0]        I861bd8df5caf968dc6edd7a05d690033;
wire [flogtanh_WDTH -1:0]        Ifb8b3586a5b69b20cf03eabf51344ab6;
wire [flogtanh_WDTH -1:0]        I6f44882493f9eadbdbe1ac46a3d2a43b;
wire [flogtanh_WDTH -1:0]        I9ea09f27ce4484f2e7fc3a6b6d6ecb7c;
wire [flogtanh_WDTH -1:0]        I5a3ec39885fba8d015009d671a1cb544;
wire [flogtanh_WDTH -1:0]        If0b9225e759438be175c4128c78605ea;
wire [flogtanh_WDTH -1:0]        Ic4e6d76148a8170d1af0c95f370367a5;
wire [flogtanh_WDTH -1:0]        I33d941ad9d4858fcfb77f0f6cf99d2ec;
wire [flogtanh_WDTH -1:0]        I244bd772f9d750b4e1800e0b0ca67d63;
wire [flogtanh_WDTH -1:0]        Ia0868eee7e7e0640ce1a4d3ca9c001cb;
wire [flogtanh_WDTH -1:0]        I00c203d60e09f1cccdadb8ebff2de650;
wire [flogtanh_WDTH -1:0]        Icb3ab2c67a87b2ee158e0021b72fc186;
wire [flogtanh_WDTH -1:0]        I20c7780e77b49d31808e59cae58968a9;
wire [flogtanh_WDTH -1:0]        I5b64997d083769666741c794dd92fb7f;
wire [flogtanh_WDTH -1:0]        Ia332fad029505e5975156f8e13910358;
wire [flogtanh_WDTH -1:0]        I0a3323aac825506435068f6746aee974;
wire [flogtanh_WDTH -1:0]        I9cc95185621ad5718a905092c03315f8;
wire [flogtanh_WDTH -1:0]        Ibec442c099da091afcf75a7c970bf8ea;
wire [flogtanh_WDTH -1:0]        Iba2a341076f0506aeac3769e71b91f43;
wire [flogtanh_WDTH -1:0]        If3a79ede332c39a8d2a276de833242f6;
wire [flogtanh_WDTH -1:0]        Ic9e82f153d0e690d5ea47ee159523b72;
wire [flogtanh_WDTH -1:0]        I49ccb3e14fe61618806e791ecb4f4eae;
wire [flogtanh_WDTH -1:0]        Ia265b95249953a7867c611d475d01169;
wire [flogtanh_WDTH -1:0]        I461ebbf3a02ae63e2eb27531b1370f24;
wire [flogtanh_WDTH -1:0]        I5ef2899606d7f08aa6d0028f9f113e38;
wire [flogtanh_WDTH -1:0]        Ice66c108aa66981051df71e226cb0e4d;
wire [flogtanh_WDTH -1:0]        Idf3a6723fec1ef62c1e37a419590122c;
wire [flogtanh_WDTH -1:0]        I645ff0d8c0a87ba7f792fc83f342b958;
wire [flogtanh_WDTH -1:0]        I0bde2fc197586c74374ffb402956baf5;
wire [flogtanh_WDTH -1:0]        Ica94017f26e96fb22a47add326ee126e;
wire [flogtanh_WDTH -1:0]        I9182b3349816b6ddaffde1cbec78339e;
wire [flogtanh_WDTH -1:0]        Id32e7ad5b1aa825732d9b26d0fa02ca1;
wire [flogtanh_WDTH -1:0]        I5bf9702e2afd6c791b28c76c84aeb886;
wire [flogtanh_WDTH -1:0]        I51b5e641856239367cf43f9b5679b268;
wire [flogtanh_WDTH -1:0]        Ifbd7b868d9cb7e04bf2189922bcb9c92;
wire [flogtanh_WDTH -1:0]        I2d1a5645b126761fc7fb70d24e37189a;
wire [flogtanh_WDTH -1:0]        Ib78e7602e521bc064d5cd9efe10ec6b1;
wire [flogtanh_WDTH -1:0]        I49f5f87662fbb540d72c94bfd1acd060;
wire [flogtanh_WDTH -1:0]        I0497115b3dd67c6538039969368e03ae;
wire [flogtanh_WDTH -1:0]        I30253dc91301ca27b5732312c01145e0;
wire [flogtanh_WDTH -1:0]        Ieba8e28ee660b8e2d78909d61ced3233;
wire [flogtanh_WDTH -1:0]        I143f5e324716a94d24ada126886bf895;
wire [flogtanh_WDTH -1:0]        I12e6fe32f6159ce6bb8be6411af2b7bb;
wire [flogtanh_WDTH -1:0]        If64aa8c220b9ab6652e081da7e404e80;
wire [flogtanh_WDTH -1:0]        I03392e42f99b06cb65b38122c1e4dc81;
wire [flogtanh_WDTH -1:0]        I1092325b801600fa7ec85fa640167da9;
wire [flogtanh_WDTH -1:0]        I32270eb6cf0594020ee19abb2edfe93d;
wire [flogtanh_WDTH -1:0]        Ib028686da9c849e827cf249a744b7db3;
wire [flogtanh_WDTH -1:0]        Ib135d3d7d338f5ff3a1f504aec754bbd;
wire [flogtanh_WDTH -1:0]        I5f3ff7fa8686f7a380302d71b88cfb4b;
wire [flogtanh_WDTH -1:0]        Id9cbc2e4b0f437840f028c7273d49416;
wire [flogtanh_WDTH -1:0]        Ic01904f7c518990eff2dc1de127676c4;
wire [flogtanh_WDTH -1:0]        I98b5a84c247422b51abf63a705fbb5f7;
wire [flogtanh_WDTH -1:0]        I43f2ddd9780f86af489f8deae51168ec;
wire [flogtanh_WDTH -1:0]        I0ae39e89061b4f8c5c0e56eba2f48889;
wire [flogtanh_WDTH -1:0]        I0a013fff6c792363bd7feb03d9691db8;
wire [flogtanh_WDTH -1:0]        If612cf94a3cefcfb844d6e975ba4aada;
wire [flogtanh_WDTH -1:0]        I7cf8401bf6893eab0b9f33a0f91ddd05;
wire [flogtanh_WDTH -1:0]        I3dab04eb1045e1b3b6bb47e0f4c390ad;
wire [flogtanh_WDTH -1:0]        Ic7ccbeaf4ab94d0660eb7a0533723e24;
wire [flogtanh_WDTH -1:0]        I447db5cb14c9588418037bbb793a6274;
wire [flogtanh_WDTH -1:0]        I08043393cb7f2558c145a698ea6652c9;
wire [flogtanh_WDTH -1:0]        Ic1227b130f19411495bed64035ea317b;
wire [flogtanh_WDTH -1:0]        I84865c4f872c0845124b78fabf695c2c;
wire [flogtanh_WDTH -1:0]        I6861b48d33277dd057c6f09ba630d700;
wire [flogtanh_WDTH -1:0]        I57b9dd7a7deea6695dcd03439c9723cf;
wire [flogtanh_WDTH -1:0]        I022bebca44e2f0b8f9877dd0e709b29f;
wire [flogtanh_WDTH -1:0]        I1cd6b35bcdfd461db69a4c1bdb1d387f;
wire [flogtanh_WDTH -1:0]        I8e3d5a48955fe19e24975579d55f4e14;
wire [flogtanh_WDTH -1:0]        I40a1ecabded8add5bffe316f2d8beda9;
wire [flogtanh_WDTH -1:0]        I7ee915ffb1c7b8985788c5e6af532ce3;
wire [flogtanh_WDTH -1:0]        I7c52ae4af926267b5e27a530202fcce0;
wire [flogtanh_WDTH -1:0]        Ia897087d82c2deac4697755c31766241;
wire [flogtanh_WDTH -1:0]        I1a5c6c50817db8bde279d5f0b5095d76;
wire [flogtanh_WDTH -1:0]        I4c23326dc80b54231289f9f18c4db711;
wire [flogtanh_WDTH -1:0]        Idf0c1b85712fcbbbcc12915158ebff62;
wire [flogtanh_WDTH -1:0]        I8326b063a9b9688fb3014667c49ada1b;
wire [flogtanh_WDTH -1:0]        I6b32298e8c61e75d0a38bca3084c0528;
wire [flogtanh_WDTH -1:0]        Ic41133a438fcea4a1cad9f5e5ee05a03;
wire [flogtanh_WDTH -1:0]        I5b0d72cedc120406402076148e2d30b0;
wire [flogtanh_WDTH -1:0]        I1ac5e426032b874b250cb8adad5b345a;
wire [flogtanh_WDTH -1:0]        Iaf624549f73b0d13c1a73c850b99f810;
wire [flogtanh_WDTH -1:0]        If9aca7e28f987bf6c7f2fb9b6f11962f;
wire [flogtanh_WDTH -1:0]        Iaaf7efeae9f6dc9e8222dc2b10122000;
wire [flogtanh_WDTH -1:0]        Id98a58cd8017fd149ea4f5b295f7ec80;
wire [flogtanh_WDTH -1:0]        Iea1cd2321d2ac9b891b344e2ba2363d3;
wire [flogtanh_WDTH -1:0]        Ib9e45e75ce8cdd3b548eaf3e41a091ce;
wire [flogtanh_WDTH -1:0]        Ia544fa24b953fe91800978895e3e610e;
wire [flogtanh_WDTH -1:0]        I9fcedcbd532cefe1e66ec94b22457cf4;
wire [flogtanh_WDTH -1:0]        I7fa710c37f5f96c3cdc35612a702a71c;
wire [flogtanh_WDTH -1:0]        Ic627802cf228a709638c14adf83091f8;
wire [flogtanh_WDTH -1:0]        I98fd105696fca11c1075f9bd30013747;
wire [flogtanh_WDTH -1:0]        Ib6bd27a683e11d238fcb775bb44dd913;
wire [flogtanh_WDTH -1:0]        I61345963ceabdaa0f25f8a463fc9fe5d;
wire [flogtanh_WDTH -1:0]        I3affcbe66b25dc7f11f98b4e444937a2;
wire [flogtanh_WDTH -1:0]        I9e8375af6af10f4bac3e87e416d430ee;
wire [flogtanh_WDTH -1:0]        Ib537657951962c85ad92d43777458588;
wire [flogtanh_WDTH -1:0]        Ida1cd844022bbf1b8431225e66b2b78f;
wire [flogtanh_WDTH -1:0]        Id0af2b1d8b0aa3ba9764ea6a22fafc8c;
wire [flogtanh_WDTH -1:0]        I30e9ab592e97dbc5fb6ab58d2ffbf8d4;
wire [flogtanh_WDTH -1:0]        I3f934c17beeba9f2d2ca58b3677fe1f3;
wire [flogtanh_WDTH -1:0]        I2ec2a6de2be39b1bc259b0be72e35a0f;
wire [flogtanh_WDTH -1:0]        Ie3e094ae62dc2a694777f4792c78c886;
wire [flogtanh_WDTH -1:0]        Ic32e349efae2ca419e095ee5e15a501d;
wire [flogtanh_WDTH -1:0]        Idea1d2f5e910ebadc99d356dee8646bd;
wire [flogtanh_WDTH -1:0]        I1befb935ee9cb871c9a7476c1fc0da3f;
wire [flogtanh_WDTH -1:0]        I7cf160bea55d67417a4ee9ce9b252871;
wire [flogtanh_WDTH -1:0]        I01c57f697f2af7d2c6ae904319f10725;
wire [flogtanh_WDTH -1:0]        I196915263bfb62cc21659f81572438b4;
wire [flogtanh_WDTH -1:0]        Id580f8a2748efff9b6b747c497c16e9c;
wire [flogtanh_WDTH -1:0]        I548af5c4ccd2816978de565c0c02f176;
wire [flogtanh_WDTH -1:0]        I77b54488bd26318f14b4364035cd1836;
wire [flogtanh_WDTH -1:0]        Ifb7004286169cd9b229b083aea58a408;
wire [flogtanh_WDTH -1:0]        I786338397f55073dce91e1c8c5f8e298;
wire [flogtanh_WDTH -1:0]        Ib04408fcc6f4d26fcdb5599b03b1b534;
wire [flogtanh_WDTH -1:0]        I0e5931219d94c8e8e1f4af081404dcab;
wire [flogtanh_WDTH -1:0]        Ifda1a58a6f54318a30faa98dc1982e8e;
wire [flogtanh_WDTH -1:0]        I8d96b419b010f8076311420d7b9c8a18;
wire [flogtanh_WDTH -1:0]        I799ce64e6df49e2b62dc6beda4500146;
wire [flogtanh_WDTH -1:0]        Ife13f962c7a8df3845cde104a959f678;
wire [flogtanh_WDTH -1:0]        Ia592b65aa89be2fcd981cf144683a298;
wire [flogtanh_WDTH -1:0]        I7f701ff37ad3fc34d2f4efafe5ff5351;
wire [flogtanh_WDTH -1:0]        Ib52365bf14aedf524bb23a4a6fe10551;
wire [flogtanh_WDTH -1:0]        I43c815a8ce0b2df9744a525328969691;
wire [flogtanh_WDTH -1:0]        Ieba74e8bf3d692612c544af3ce6046fd;
wire [flogtanh_WDTH -1:0]        I6c4a1ded9bf39091cf302ebe0103e2f0;
wire [flogtanh_WDTH -1:0]        I6cc1587e659f3f97d636485b708b1eeb;
wire [flogtanh_WDTH -1:0]        Icd4ff8d14af2699db2b5168027894ebb;
wire [flogtanh_WDTH -1:0]        I84b09aba55d2335f19faa5762aeedb89;
wire [flogtanh_WDTH -1:0]        Ia79d52fe2130426c07890fcaa50137db;
wire [flogtanh_WDTH -1:0]        I3c4b9082ba72cade4d52924eff135135;
wire [flogtanh_WDTH -1:0]        I308aaa8ac500b5589aa4af533a9062bf;
wire [flogtanh_WDTH -1:0]        I65f6c14ae4e7139fd858d7637ec3fd46;
wire [flogtanh_WDTH -1:0]        Iac91f4037e542d9fda30fadafe7e79ac;
wire [flogtanh_WDTH -1:0]        I02425810db970e5ef0b791dc4be103a9;
wire [flogtanh_WDTH -1:0]        I8cd5970682bc84881489c12ff073212c;
wire [flogtanh_WDTH -1:0]        Id0bc7b00dec58136a8016979d8a9faad;
wire [flogtanh_WDTH -1:0]        I1ee27be7e1a38aff0039b21c45f406d1;
wire [flogtanh_WDTH -1:0]        I7c61892052c3c32343ed172d4ae354cc;
wire [flogtanh_WDTH -1:0]        Idf90f01353ad1057e11fd060442f4e53;
wire [flogtanh_WDTH -1:0]        I7cd312338aa5a86e1b05cc28ab7a2b23;
wire [flogtanh_WDTH -1:0]        Id45f4e0f142b6c3925f24a37dcf7c0ae;
wire [flogtanh_WDTH -1:0]        I88d4372b4f7bfddd2af726c2df391287;
wire [flogtanh_WDTH -1:0]        I52a9bcfbd2d3a763671f19cfeaf7bb8b;
wire [flogtanh_WDTH -1:0]        Ic8978ad86275ac6f4a0cf80ebefc5b27;
wire [flogtanh_WDTH -1:0]        Ia3cc6acf2cae41e560e09993007ffd2b;
wire [flogtanh_WDTH -1:0]        I99745124c45f37d3882064590394a0aa;
wire [flogtanh_WDTH -1:0]        Iba0d2f08788f2208a648ae7b5414195d;
wire [flogtanh_WDTH -1:0]        I33fe34f9be3c51b4b93f89c3f862e332;
wire [flogtanh_WDTH -1:0]        I9f7df6ad60284c812aeb522974578e0b;
wire [flogtanh_WDTH -1:0]        Iecda9a183e74f78b9fd5ce34e80d712e;
wire [flogtanh_WDTH -1:0]        Iab1fb7006598181bd8749ed90c519b13;
wire [flogtanh_WDTH -1:0]        I5293b996bbf152abf110df1205ad4856;
wire [flogtanh_WDTH -1:0]        Ieef3b299ec35075c71ef9fb10525bfc4;
wire [flogtanh_WDTH -1:0]        Ia99c08ee345bdc1489ce82a62481ef3b;
wire [flogtanh_WDTH -1:0]        I58a7c08adf48d0737c5803e2a818c045;
wire [flogtanh_WDTH -1:0]        Iaa314530e04145eb73672ebb150858af;
wire [flogtanh_WDTH -1:0]        I30a1c8fcd9a510a6ed559f07dd809b90;
wire [flogtanh_WDTH -1:0]        I05f7363bfcc34691280079e82f6f5449;
wire [flogtanh_WDTH -1:0]        Ic4f5e9d49419e1c57cfa387761ab643d;
wire [flogtanh_WDTH -1:0]        Ica5ce135e77ed1d7cbc8277344ffeaeb;
wire [flogtanh_WDTH -1:0]        Id3dd71ea0bf0f2996fbe42b8c3318762;
wire [flogtanh_WDTH -1:0]        Iac98c702c4d9d78460fc7c212bce7841;
wire [flogtanh_WDTH -1:0]        Ib834b91bf81067e8efa9d470023e8b9d;
wire [flogtanh_WDTH -1:0]        I1fe269380ba03e78a8e41c17aa4bd757;
wire [flogtanh_WDTH -1:0]        Ic6ead78ed741442f17a15a157cd6ef9c;
wire [flogtanh_WDTH -1:0]        Ib19549130ee3307413b69c50042f7302;
wire [flogtanh_WDTH -1:0]        I4e257dbd6f196a02dc0f5a2e5f6047d7;
wire [flogtanh_WDTH -1:0]        Iad6acaf97d307fdbe0f20bf010acb468;
wire [flogtanh_WDTH -1:0]        I3dbfbd34d1fdfd4f422d900154123b6b;
wire [flogtanh_WDTH -1:0]        I67c9882f9e19df5a7b9bd0d900bb2f75;
wire [flogtanh_WDTH -1:0]        I529b763dace1924613d184c6c70c2708;
wire [flogtanh_WDTH -1:0]        I3099768bc986a11350656e472fc21ac1;
wire [flogtanh_WDTH -1:0]        I7a600aeb6cf8c3311c10afa4d82767a1;
wire [flogtanh_WDTH -1:0]        Ifba5972f9d38199dbc675432a29934e4;
wire [flogtanh_WDTH -1:0]        I8c7aab31f8cb705ea13a41a5bd349303;
wire [flogtanh_WDTH -1:0]        I0934fb292b19451a050fb3374a7bd1a7;
wire [flogtanh_WDTH -1:0]        I171149dcaab2c0f0e2a10547ad95084d;
wire [flogtanh_WDTH -1:0]        I9a3d1741c77fb1bbc1a54383874de82a;
wire [flogtanh_WDTH -1:0]        I23b60ca4da2df0ec40c1df62d058deef;
wire [flogtanh_WDTH -1:0]        If89f2ce813bab91af88f73ddc570d5a1;
wire [flogtanh_WDTH -1:0]        I7978d2d800b4438d0644ae3df6bcac9c;
wire [flogtanh_WDTH -1:0]        Ibc0dfcffac26f4898d42808534f6588f;
wire [flogtanh_WDTH -1:0]        Ibc4eddc0f1768e9ec7e38e951a28ec42;
wire [flogtanh_WDTH -1:0]        I3a0a6f3d0141e8ad04d89c4bf306a96f;
wire [flogtanh_WDTH -1:0]        I1c97fd1d21a31af8b5498a79b1a3e7b6;
wire [flogtanh_WDTH -1:0]        I1c875571dd1be1bb28aa15554964b485;
wire [flogtanh_WDTH -1:0]        Ie4f063eeaf7ee3f033e2a01ffaca623e;
wire [flogtanh_WDTH -1:0]        Ide5d5fdcf86b369b015890030a222a0a;
wire [flogtanh_WDTH -1:0]        Ibb3d57d510cad00064a331f61f6400a2;
wire [flogtanh_WDTH -1:0]        I7cf6e8d40e7bd7685a7260638523690c;
wire [flogtanh_WDTH -1:0]        I9485ae915474a31562ce358666d66245;
wire [flogtanh_WDTH -1:0]        I52ccac771cc9a1c1797862bc781e1f58;
wire [flogtanh_WDTH -1:0]        Ia54b6f7044a831020e49f1bf48bc063a;
wire [flogtanh_WDTH -1:0]        I9db2090916f2535b14ed3292e78baa32;
wire [flogtanh_WDTH -1:0]        Ie71c7babb5d17378d40444b6bbd4e7a6;
wire [flogtanh_WDTH -1:0]        I5b77a8ce7f495ae61315d1590bfd71b8;
wire [flogtanh_WDTH -1:0]        Ia0977b79857bdbf058535c30e338c38a;
wire [flogtanh_WDTH -1:0]        I4e4bb795cf09757c8ad3933c9ce4686f;
wire [flogtanh_WDTH -1:0]        I600ea1371a2be66430ac9534583b512b;
wire [flogtanh_WDTH -1:0]        I78c29808e737dab48b5144b232dd02f6;
wire [flogtanh_WDTH -1:0]        Ife5b9afdbb30c122b84d5378f9cb366d;
wire [flogtanh_WDTH -1:0]        Ie2ae83a457d79fbddc640d49d626171c;
wire [flogtanh_WDTH -1:0]        I27556d599dd1a27ee8f49e819ccbf29a;
wire [flogtanh_WDTH -1:0]        I3711e49a4eec517e47897fb731d75958;
wire [flogtanh_WDTH -1:0]        Icce595233ce089eafcca3eae5e71e5f8;
wire [flogtanh_WDTH -1:0]        Ifda4e727eb6275266f583badb6d4a9ed;
wire [flogtanh_WDTH -1:0]        Icc3cadf40c09be1a8c2847caf0e3e63c;
wire [flogtanh_WDTH -1:0]        I2be66a82c7b58e3c14b5816522b46969;
wire [flogtanh_WDTH -1:0]        Ib43886d923b8c683004713ff25b2f90d;
wire [flogtanh_WDTH -1:0]        I826fe7ad9e67061800d5d6543d779864;
wire [flogtanh_WDTH -1:0]        I132d9671c582876568c0f7f5335f5227;
wire [flogtanh_WDTH -1:0]        Ic0c9069041758b53f56a46da81dd2d60;
wire [flogtanh_WDTH -1:0]        I0859c80b42a8c60dade8f05d58ee3701;
wire [flogtanh_WDTH -1:0]        I6f4c5a8de7690fec959861f43c134915;
wire [flogtanh_WDTH -1:0]        Ib3690ec149adde94343d3e617931a287;
wire [flogtanh_WDTH -1:0]        I14f1005a8c0fbdc5ca02c032b8891c2b;
wire [flogtanh_WDTH -1:0]        I41f2bf9ff00f983ad1298c8c83b041cb;
wire [flogtanh_WDTH -1:0]        Iacd30dfb96f6572ec56eff0a4094ec04;
wire [flogtanh_WDTH -1:0]        Ib5414585cd6976cfce42e42190cc08d7;
wire [flogtanh_WDTH -1:0]        I1c748b8fe4979331bc3fe5aff4b6f9f4;
wire [flogtanh_WDTH -1:0]        I1ca59325ff30db83df5bf0a2cd9706b6;
wire [flogtanh_WDTH -1:0]        I158c7973974f36c2793127964e50d1bd;
wire [flogtanh_WDTH -1:0]        Ie2f5b03f3b136e651b8aba92a30d298a;
wire [flogtanh_WDTH -1:0]        Id5ea6ba2402275cb925a1848b31ec2e1;
wire [flogtanh_WDTH -1:0]        I312ce79a8dd2ce3d37c930d42640509b;
wire [flogtanh_WDTH -1:0]        I3862f7017bc2bc69844b73f2a79f47f5;
wire [flogtanh_WDTH -1:0]        I467d5e2554ef25873e0b44e947ee0011;
wire [flogtanh_WDTH -1:0]        I4ed41fde5449b7112baf000a05484ac4;
wire [flogtanh_WDTH -1:0]        Ice73b514709469fd21cd254bf4ceadd9;
wire [flogtanh_WDTH -1:0]        I40c4db2872b602bf9d6a4fc4ba5ac34d;
wire [flogtanh_WDTH -1:0]        I45ba06a6d6f00c174b1439a6f226a085;
wire [flogtanh_WDTH -1:0]        Ibe5ab52bd0f220f7a6aac244c0e3867e;
wire [flogtanh_WDTH -1:0]        Ic8a272f82736fd599fb3250e970edf9b;
wire [flogtanh_WDTH -1:0]        I36668064f280c70f9143ee9f39973015;
wire [flogtanh_WDTH -1:0]        I5b9710b16effc8bf0695517c6e651836;
wire [flogtanh_WDTH -1:0]        Ief92462253c5a03a42d46ed7087caf9a;
wire [flogtanh_WDTH -1:0]        I038b42a83025f5eaebf45799d1ebe7b0;
wire [flogtanh_WDTH -1:0]        Idf196345491ff3290796ba7827d31c17;
wire [flogtanh_WDTH -1:0]        I73ddd7cf9272ceab5a663e2244e72d7e;
wire [flogtanh_WDTH -1:0]        I2230f0e48899877bc2bcb3538be81bfa;
wire [flogtanh_WDTH -1:0]        I16507fab8f9076bfeb419896fa7cdc1d;
wire [flogtanh_WDTH -1:0]        Ibc0ec83d6b8e6be89ddc88ef83f0b03d;
wire [flogtanh_WDTH -1:0]        I3dd1f28cf199299aba54e47a429c9b11;
wire [flogtanh_WDTH -1:0]        Ifc59c1b26ec09b3a7fe5a2b90511c93b;
wire [flogtanh_WDTH -1:0]        I49d9203dc6f8c17f17383e8f7e01f005;
wire [flogtanh_WDTH -1:0]        I9c6fc8e09cd63551f40accc98d784a44;
wire [flogtanh_WDTH -1:0]        Ibeec86c75d950ee00dd63a2930f08a24;
wire [flogtanh_WDTH -1:0]        I26692a6aab1d81d71219a436bee5e10b;
wire [flogtanh_WDTH -1:0]        I47b2438c3680b2d816168df37d7c491c;
wire [flogtanh_WDTH -1:0]        Ieb50592e17305d0f74cbf216be947862;
wire [flogtanh_WDTH -1:0]        I5983bf2c6c90b872ee6cf58b5e520311;
wire [flogtanh_WDTH -1:0]        I0071f023f1be4400541c13bc68278417;
wire [flogtanh_WDTH -1:0]        I6745cacecb7ee86cf3c7ad7eeee6048f;
wire [flogtanh_WDTH -1:0]        Ib2f1635b38ca6090e5ff633cbfa13273;
wire [flogtanh_WDTH -1:0]        Ib9672d20643d856ff31905ab14c0ac87;
wire [flogtanh_WDTH -1:0]        Id2c0bc90fd26e82fe91b5aef7bdd3a29;
wire [flogtanh_WDTH -1:0]        Ib9dfea1f34a120eda30d5bd919365a6a;
wire [flogtanh_WDTH -1:0]        If4a723ce836f5327b85e234ebd195bd9;
wire [flogtanh_WDTH -1:0]        Ia7bf82c9e5ca4467b5e50beeaeb975e9;
wire [flogtanh_WDTH -1:0]        If63dd5997e033817126a9ebaf38c1955;
wire [flogtanh_WDTH -1:0]        I327c9acb8934729b4ea5486787afa2e8;
wire [flogtanh_WDTH -1:0]        Ie2ee6baf8ec357f6131dff92fb480e42;
wire [flogtanh_WDTH -1:0]        Ieddef08050c38d07e5d38f5bb7b099c0;
wire [flogtanh_WDTH -1:0]        Ibff4d4fca3681fe10807414ed84e4157;
wire [flogtanh_WDTH -1:0]        I39f9e8430db114991bfb27cc46ef3e39;
wire [flogtanh_WDTH -1:0]        I4540d74c919f50e9b6e40ef6b8cfd279;
wire [flogtanh_WDTH -1:0]        I56aa548618a4a15e9a35e04f5eeb823f;
wire [flogtanh_WDTH -1:0]        I01637ffca829d72accbb5dcee48817ca;
wire [flogtanh_WDTH -1:0]        I1908897b529ca04df7e7da395be4a8ce;
wire [flogtanh_WDTH -1:0]        I7e8af960e934c7cc3cb163d6f8e7d597;
wire [flogtanh_WDTH -1:0]        Ib2bbd59cd6098608ed53ac556036534f;
wire [flogtanh_WDTH -1:0]        Ifd80d371c8851b9e16193a3e62ddf79a;
wire [flogtanh_WDTH -1:0]        If004552b2047ab1cf23bb50375460b01;
wire [flogtanh_WDTH -1:0]        I19d2c4bc969133fa59d22f7f2d8cfd4a;
wire [flogtanh_WDTH -1:0]        If97092e1e2147de199c94a23831cf6b9;
wire [flogtanh_WDTH -1:0]        I532326ad245909d441134296dae9a5d4;
wire [flogtanh_WDTH -1:0]        Ibf74a4dfaab7f7f538d2b5fac7394b63;
wire [flogtanh_WDTH -1:0]        I6ca7199e28b480ac5816bf5b4cfb1eef;
wire [flogtanh_WDTH -1:0]        I991a7a7d562eb0a8b4b8d8f008ef2225;
wire [flogtanh_WDTH -1:0]        I0d5b26d24fbce6b236120b5697d0db6b;
wire [flogtanh_WDTH -1:0]        I64c3d7be41abaa17d6992f9af8e72789;
wire [flogtanh_WDTH -1:0]        I618d329f2b0f18617d80aa350b79601c;
wire [flogtanh_WDTH -1:0]        Icb91e63ebabc7a75a54eb7c731df4fa0;
wire [flogtanh_WDTH -1:0]        I58e3a5e842e14d09de91959839798a67;
wire [flogtanh_WDTH -1:0]        I673d1d0d0daab99bd940c46cc14ef55a;
wire [flogtanh_WDTH -1:0]        Icdecd5095ef818a0915ff3fcb395db5b;
wire [flogtanh_WDTH -1:0]        I62cadbd70b07a6a7a2974c7c392696b3;
wire [flogtanh_WDTH -1:0]        I236f843994d3065b6ee70c41f390a3d0;
wire [flogtanh_WDTH -1:0]        Icd8257d7f53d93db989eb56eaeb7e593;
wire [flogtanh_WDTH -1:0]        I7a9001d6c1d1aa8af79d9b152e596b70;
wire [flogtanh_WDTH -1:0]        I05931ceae6eff26e5a66a44a54d628ae;
wire [flogtanh_WDTH -1:0]        I56a43a072d463792d9e676c4907b3e76;
wire [flogtanh_WDTH -1:0]        I306fec0aa68a0396053a6e0fa1cda38f;
wire [flogtanh_WDTH -1:0]        I336a86e85d3a8a42c4b6458ccb92ae05;
wire [flogtanh_WDTH -1:0]        Idee8c8144207d676d1f2f9064bbdff45;
wire [flogtanh_WDTH -1:0]        Id97f66b78f1e3b6bf0b962b85ca1cde7;
wire [flogtanh_WDTH -1:0]        I5855124d566af739caa6511f8598f2c5;
wire [flogtanh_WDTH -1:0]        I52c7f0a8f9b4533052b5acd1b5bd5e17;
wire [flogtanh_WDTH -1:0]        I50729db4a8e04f18979707df14cb2419;
wire [flogtanh_WDTH -1:0]        I3b1db672b1a94502b90451260062a274;
wire [flogtanh_WDTH -1:0]        Ia3cb3ea64576a3e7332e1fb55953aa3e;
wire [flogtanh_WDTH -1:0]        I1a83f91eb1262911ae8d99e305294bf8;
wire [flogtanh_WDTH -1:0]        I3cb1f233951d49f985b0deac6e052bfd;
wire [flogtanh_WDTH -1:0]        Id01bfbd86b6321a843e239ca97cec514;
wire [flogtanh_WDTH -1:0]        I7015def91103398e54f446ce3e43af01;
wire [flogtanh_WDTH -1:0]        I26b769b58e1c21b68dd95c9f38c0362b;
wire [flogtanh_WDTH -1:0]        I04874bd1bf257f205b5189c8c20e5a12;
wire [flogtanh_WDTH -1:0]        Ic86f9988281398adfe43152beb722c1b;
wire [flogtanh_WDTH -1:0]        I937e3a8ede2305ea7c1750283224a870;
wire [flogtanh_WDTH -1:0]        I9d8ac6c29c2f5df7c2d124dface59e35;
wire [flogtanh_WDTH -1:0]        Ia7206430a739a11af4d860096eedd6c3;
wire [flogtanh_WDTH -1:0]        I56b46c426895409b40c3be9b79365a8a;
wire [flogtanh_WDTH -1:0]        Ibf4c2c00f8e012e9498361bfd3c5b06e;
wire [flogtanh_WDTH -1:0]        Ic63de8464f79ae05f27f05c935dbf495;
wire [flogtanh_WDTH -1:0]        I899e5f03cd1d52d11f898959559aaeea;
wire [flogtanh_WDTH -1:0]        I4d21ee443e5921532d5bf1db7ef93f82;
wire [flogtanh_WDTH -1:0]        I59c80c7ec26f43308b1a646c47160568;
wire [flogtanh_WDTH -1:0]        Ieb5fa20abbdb29a7f75021b7afafea31;
wire [flogtanh_WDTH -1:0]        I8a954a331d36266465a0813d2e8b319b;
wire [flogtanh_WDTH -1:0]        I16a12326344aadf4226bd149424a53a8;
wire [flogtanh_WDTH -1:0]        Ib49e53ca8efd9564ee9572eb3089bb51;
wire [flogtanh_WDTH -1:0]        I07f36b533b48344c13dbb133739712f4;
wire [flogtanh_WDTH -1:0]        Icbde2c6230e9cc67ef12031e38bb344f;
wire [flogtanh_WDTH -1:0]        I7a0072bf1e5fb0c4de85c6e4447878a4;
wire [flogtanh_WDTH -1:0]        I2e22e867f6f84a7807b82f64a147022e;
wire [flogtanh_WDTH -1:0]        I320bafc5a1775d6933bcb9f2d2c84576;
wire [flogtanh_WDTH -1:0]        Id9704e1d8096cd28577c5c357d30b7a4;
wire [flogtanh_WDTH -1:0]        I5ec61756ff7237146f2d83f17eb5bb3a;
wire [flogtanh_WDTH -1:0]        I4b8554cab486a4fc1e14884a6495016e;
wire [flogtanh_WDTH -1:0]        I382008a17338641e68fa859ac2af1d20;
wire [flogtanh_WDTH -1:0]        Iaa235d085a5916a3b0814c3ed2a9026f;
wire [flogtanh_WDTH -1:0]        Ifd375ad8038ea2455c0e3b1463b83b7e;
wire [flogtanh_WDTH -1:0]        I5d86ce0b58c0b281d747116a9069ef33;
wire [flogtanh_WDTH -1:0]        I0b75763235278d8eca6ca72fc97fb83c;
wire [flogtanh_WDTH -1:0]        Id20394136fb036435bb4680aac64581f;
wire [flogtanh_WDTH -1:0]        I9bc4c3b77a9635bb77ad31527d961952;
wire [flogtanh_WDTH -1:0]        I8a16afac6e470ca69634d7fe9656387a;
wire [flogtanh_WDTH -1:0]        Ief93f4a7eaaa1f43ea1788dc4629c093;
wire [flogtanh_WDTH -1:0]        Ic4e7f690bc050f1d1f84eae7ca193e1c;
wire [flogtanh_WDTH -1:0]        I34b86fbc3949cb2083931ad8edd2444d;
wire [flogtanh_WDTH -1:0]        Ia60421aa427236540b4d0d08d52ff507;
wire [flogtanh_WDTH -1:0]        I560c163fb55aa4b56da25f96e9b8ef6c;
wire [flogtanh_WDTH -1:0]        Icace650ee3865bd7bbddd2d9435c5561;
wire [flogtanh_WDTH -1:0]        Ib3c46d34c5bc3d2651147b3e764d9786;
wire [flogtanh_WDTH -1:0]        I7d27d070b96b7810f667e1d1845342d3;
wire [flogtanh_WDTH -1:0]        Ie5e2ba4fe22870afc81d6cfc708570be;
wire [flogtanh_WDTH -1:0]        Ida7ec09c913caa0e78a2c4cbaae517c8;
wire [flogtanh_WDTH -1:0]        Ibf3bde181da4f960537516d6c0b2a72c;
wire [flogtanh_WDTH -1:0]        Ic5eba898858be1f768841ead792d6d86;
wire [flogtanh_WDTH -1:0]        Ia93f96aa0718f8755e9ebb8cc5d8f405;
wire [flogtanh_WDTH -1:0]        I72197797a307c611fa8952533e63d7bf;

reg                              I3c62d5bd891bd3750b7bd1d32612f589;
reg                              I699819696b0299ab80e7233d054ec590;
reg                              Iac11baea9832d6493626d2fe40fd385f;
reg                              I92354deea988f3beb25bfba90735c6ac;
reg                              I6d3acefe6d7dfb94a5d66dcaa1bbbb76;
reg                              Ibd047e2643dc68affb5b4f25b82ded31;
reg                              I65e382d77592c7d1af308d171b27ff3c;
reg                              I7d4dc5e91ba3d952184d90de12f67bd3;


reg  [fgallag_WDTH-1:0]         Ifeb14203f4daf31c7701a6a742be57cc;
wire [fgallag_WDTH-1:0]         Ic188ebb37ff178022c61400613f4f3dc;
wire [fgallag_WDTH-1:0]         I5a11c8e7d2b7d4c0253df9015b7f3ab5;
reg  [fgallag_WDTH-1:0]         Ib581c19864deecf01268595049268b19;
wire [fgallag_WDTH-1:0]         I3f80921fd94cff373648fa34fcadd4d2;
wire [fgallag_WDTH-1:0]         Ib0740d8c9ab158e682432a0e3ec89798;
reg  [fgallag_WDTH-1:0]         I661d84af541e30828bcbd962d72baba3;
wire [fgallag_WDTH-1:0]         I229f7430f590d86a323b48806beec48c;
wire [fgallag_WDTH-1:0]         Ibb6505392d5b3be76542bb0303d46876;
reg  [fgallag_WDTH-1:0]         I1c6928cccb4bf7ea7dfd74e425b9624d;
wire [fgallag_WDTH-1:0]         I26fa0a5f87600d9535e8f83fa1a11136;
wire [fgallag_WDTH-1:0]         If23edf1bc3801016b24252fbc3d33508;
reg  [fgallag_WDTH-1:0]         I6eabc5c074fb1e2183a5f1ecee87a518;
wire [fgallag_WDTH-1:0]         Id87360986474c9bfa5266a90b59a9a8b;
wire [fgallag_WDTH-1:0]         I47478ccbfc4c3b944d130a192fb4fb5a;
reg  [fgallag_WDTH-1:0]         I0107769bbd7c239685b4818731334437;
wire [fgallag_WDTH-1:0]         Id63daaeb52208682533b5f136480a29c;
wire [fgallag_WDTH-1:0]         I40b126fdab110e58eac80ea13bcc699d;
reg  [fgallag_WDTH-1:0]         If723180430080198d18a08d6775ab208;
wire [fgallag_WDTH-1:0]         I1e9d5c2338b6f89e43c30c0ad71f675c;
wire [fgallag_WDTH-1:0]         Ib12b389fb2603e428b72d1e712975e40;
reg  [fgallag_WDTH-1:0]         I44abc734d6acf92a8e8209186d7a1676;
wire [fgallag_WDTH-1:0]         I11cce7dd119eb0e3acafc12dbc6d3536;
wire [fgallag_WDTH-1:0]         I22b0cc5517631526be6455fc60dd5323;
reg  [fgallag_WDTH-1:0]         I72aa55988d58c664f3291b5786fc8ceb;
wire [fgallag_WDTH-1:0]         I934b111c08439d3797cb8928c7238f23;
wire [fgallag_WDTH-1:0]         Ib8aba28214fb9ee1693cafe9175831e1;
reg  [fgallag_WDTH-1:0]         Ie69528583db8155917ab3d32a446de04;
wire [fgallag_WDTH-1:0]         I508cb12fa71441b216fd7c1899d00e24;
wire [fgallag_WDTH-1:0]         Ia03282a7ed4a337981d4f5b01f564a1d;
reg  [fgallag_WDTH-1:0]         Ib22b47d95b72871e74069fe80a191680;
wire [fgallag_WDTH-1:0]         Ic69c6ea6b4f360efae87611c00b00fdb;
wire [fgallag_WDTH-1:0]         Icf75bf863d8867b0fe354017921aeae1;
reg  [fgallag_WDTH-1:0]         Id9451e945bd26b8dcb4cb83ab4ade73b;
wire [fgallag_WDTH-1:0]         Ifccbe59b7ebe3f692f5b7e7564ca50ba;
wire [fgallag_WDTH-1:0]         Ia65c174738acf41b82f75be972e9022e;
reg  [fgallag_WDTH-1:0]         Iba4627d3d3ef91f168068ed128c04113;
wire [fgallag_WDTH-1:0]         Ifd7275bc534fe9da81b12b25ed218e91;
wire [fgallag_WDTH-1:0]         I587a0e70cecf4d054cc0ab53150876e0;
reg  [fgallag_WDTH-1:0]         I39bef4d462b0a3f88ce1485a58d66da0;
wire [fgallag_WDTH-1:0]         I01a99ac2a3f919f4fc1680edb11c576b;
wire [fgallag_WDTH-1:0]         I7dc71f64f9b3940721569574db6e18d0;
reg  [fgallag_WDTH-1:0]         Ib95e457d5ae9fc89e197c249414abbcd;
wire [fgallag_WDTH-1:0]         I322b3879383d75c43c55535f01fdfdd6;
wire [fgallag_WDTH-1:0]         I935ba9f8f6e9c68f75a7cb576655cab5;
reg  [fgallag_WDTH-1:0]         I2be28be47a38e9ca9d3b9167327d3d59;
wire [fgallag_WDTH-1:0]         I1adc689464e0b81fa165eb17e71310fa;
wire [fgallag_WDTH-1:0]         Ibdc981a062c989ada978f733ddff0f71;
reg  [fgallag_WDTH-1:0]         I2ee6154b613d0d86c2354604e93a9a57;
wire [fgallag_WDTH-1:0]         I2bdc0908c3d365d25f8026263dc4a258;
wire [fgallag_WDTH-1:0]         Ibcbc5e2720516c24359870ac790373f4;
reg  [fgallag_WDTH-1:0]         Ia7479d4940b575cf918cb8421f041e44;
wire [fgallag_WDTH-1:0]         Icf6c6fcfa42c48f16a1b30cd325c139f;
wire [fgallag_WDTH-1:0]         I11fdefe51f8f028fba7698870d198df6;
reg  [fgallag_WDTH-1:0]         I3c5b1cddd608ad869e0182ad68bd0494;
wire [fgallag_WDTH-1:0]         Ife8337f33629521c096d4dcfde96e879;
wire [fgallag_WDTH-1:0]         I10f17104471f87c53a589926534fc9fe;
reg  [fgallag_WDTH-1:0]         Ic4425ae997c479e05e12347a803213dd;
wire [fgallag_WDTH-1:0]         I8afa93d48ae589bb90cc74897defe4de;
wire [fgallag_WDTH-1:0]         I8fdaa3f282af2d5f053d77216c659146;
reg  [fgallag_WDTH-1:0]         I3a0518d0d382758ae579acd7e6cd634a;
wire [fgallag_WDTH-1:0]         I56d0b4df55f7f4181a51f58187d399e4;
wire [fgallag_WDTH-1:0]         I167ee185ac7beee082544897898b27fa;
reg  [fgallag_WDTH-1:0]         Ifd28c1cd286b7a483891bdd094b70db1;
wire [fgallag_WDTH-1:0]         I8ae9260d2a5dd6c2ed4b6157946e38d4;
wire [fgallag_WDTH-1:0]         I5264a25f96edda24a763298d92cdf8c1;
reg  [fgallag_WDTH-1:0]         Iadf7734be049c645819d9d023b58c4dc;
wire [fgallag_WDTH-1:0]         Ie405c3459c9caf16c0a257a059a9fa96;
wire [fgallag_WDTH-1:0]         If7d5260450e23711760a6f9e5f7aa820;
reg  [fgallag_WDTH-1:0]         I5f23af0d0853ea6de084ccf77702b78d;
wire [fgallag_WDTH-1:0]         Ie76a46f18cbb52a93a4fad65462da3e8;
wire [fgallag_WDTH-1:0]         Id1265b30a8ed85169b1837aa1b656aa2;
reg  [fgallag_WDTH-1:0]         Ic5c99c42e9ebe5dded369ac78a1bedb5;
wire [fgallag_WDTH-1:0]         I0445dbe40692ef21353aacc7b4f7a4c9;
wire [fgallag_WDTH-1:0]         I84e6c5099aaef8094f4c2bbc82989c4c;
reg  [fgallag_WDTH-1:0]         I4f2498bec0e96802b82f0419d97c527f;
wire [fgallag_WDTH-1:0]         Ie3be0f770c8ddbdf301ae23881499e9d;
wire [fgallag_WDTH-1:0]         Ibf4bfa16424f7051e80b2947ff7f5533;
reg  [fgallag_WDTH-1:0]         Icaf86e0abee612aa972388c0b6f90763;
wire [fgallag_WDTH-1:0]         I3a4d175e3b015a17f7a49cc6bacbd12f;
wire [fgallag_WDTH-1:0]         I0e138642d8ed7e30cc254d4e259e3d51;
reg  [fgallag_WDTH-1:0]         I478c4f13c05651605a2045bb5fd6b60d;
wire [fgallag_WDTH-1:0]         Id85473220f4909f9182711939cf6a978;
wire [fgallag_WDTH-1:0]         If1c79ab7bbf50d343ba3f758a31d6786;
reg  [fgallag_WDTH-1:0]         Ide67911b52687d67ef0c25f2aadf14c5;
wire [fgallag_WDTH-1:0]         If77ecdb29d692c01752be0908c4f4392;
wire [fgallag_WDTH-1:0]         Ic2d209d919c7e43f467c3f2d093c9a8c;
reg  [fgallag_WDTH-1:0]         Ie9e7630af25f39a0e820181918edd029;
wire [fgallag_WDTH-1:0]         Ia188482ea4a2696f188f637912aa6f3b;
wire [fgallag_WDTH-1:0]         I6c59651ae65c67edfa963ce797b98234;
reg  [fgallag_WDTH-1:0]         I0e1f07f30cfe36f189e9dcb4e713b5c8;
wire [fgallag_WDTH-1:0]         Ibd0c9231ee029200ca39013c839bc4ae;
wire [fgallag_WDTH-1:0]         If4b95101c6d8670411a018ed1ae697d3;
reg  [fgallag_WDTH-1:0]         I31cee5e2a93635987776b0ea477e6211;
wire [fgallag_WDTH-1:0]         I0fed2eb07a75f701ff7b7ca9dbcddb81;
wire [fgallag_WDTH-1:0]         Ib1e406a5bb0569ac2c25e7021ec58edb;
reg  [fgallag_WDTH-1:0]         I84721f2bc5ae10db78d2e7e07cc28d94;
wire [fgallag_WDTH-1:0]         I96140f2ad00cb9a1249b5135ea251bc8;
wire [fgallag_WDTH-1:0]         I8198f75286b8c817d3b69cf7537b1c38;
reg  [fgallag_WDTH-1:0]         I6c6d057e910da53aa47441566f95153e;
wire [fgallag_WDTH-1:0]         I34fecbd6c558b25e7f8d08fb10b224f4;
wire [fgallag_WDTH-1:0]         I9431b10311eda8240d91bed96a969523;
reg  [fgallag_WDTH-1:0]         Iecbf70768fbaaab8da98eaa9a2b956ee;
wire [fgallag_WDTH-1:0]         I8df49bd85a846a4c4c32af63798f3e0e;
wire [fgallag_WDTH-1:0]         Ib623d99c3d272f39c518b6a41dd03e8d;
reg  [fgallag_WDTH-1:0]         I71b8492d70b423e95938995c07395def;
wire [fgallag_WDTH-1:0]         I05be7b5c657867c4331ed3df72a1aec5;
wire [fgallag_WDTH-1:0]         I388b66a7b7e9225f7aef4699521e9250;
reg  [fgallag_WDTH-1:0]         Iae469bcbba9598bb46aa7ccf9fa06a37;
wire [fgallag_WDTH-1:0]         Id47eecb4e17f799da48d80451cb47b5d;
wire [fgallag_WDTH-1:0]         I532db075ab1b0a5a37a2085ecd0611c3;
reg  [fgallag_WDTH-1:0]         Ie2e854376f4b6509ec41507401173269;
wire [fgallag_WDTH-1:0]         Iedabb8b1ffd46b983fd74b9f6010dcca;
wire [fgallag_WDTH-1:0]         I357c21c29061134ed6e5c872836f4759;
reg  [fgallag_WDTH-1:0]         I7b1401c3c2c389d9bf05658c88ff6b40;
wire [fgallag_WDTH-1:0]         Ib032a08190a75ceb242a9dc8272b4a02;
wire [fgallag_WDTH-1:0]         I5a1d671b8b8877192d2c129be7f149c0;
reg  [fgallag_WDTH-1:0]         I88ee95aeb6c744eca0e127e8497b5dc9;
wire [fgallag_WDTH-1:0]         Ia870db84a0411e463b6e15f502323810;
wire [fgallag_WDTH-1:0]         I4d1c830053fedd74930d9992732e9542;
reg  [fgallag_WDTH-1:0]         I5573e18ade3430ef3eff5e6d960e44eb;
wire [fgallag_WDTH-1:0]         I8105600a0847cabdb96310074840bdb7;
wire [fgallag_WDTH-1:0]         Ie53c31ded4a5c8977f956e968dd5a9a7;
reg  [fgallag_WDTH-1:0]         Id6260fa8a9be077673e82344c736b1c4;
wire [fgallag_WDTH-1:0]         I7d6591184fd95d3f288f481734e85c02;
wire [fgallag_WDTH-1:0]         Id5355c3ed75d1aed52250f6f0d00b1a0;
reg  [fgallag_WDTH-1:0]         Ic052eadb342350c52d89e73d5fea80bb;
wire [fgallag_WDTH-1:0]         I69c3d2866b040d67900eeb991b7c2981;
wire [fgallag_WDTH-1:0]         Ib43ca9d864e41a89bec5344ece17fd10;
reg  [fgallag_WDTH-1:0]         I98b8d024432fc54ebf2f15d99968f2e0;
wire [fgallag_WDTH-1:0]         Ice61d34abe5e2a9593bfb911da54e959;
wire [fgallag_WDTH-1:0]         I6c7b0be00e8302794aa3a79fb2acf100;
reg  [fgallag_WDTH-1:0]         I98f54ab8454940141a484332f2a05369;
wire [fgallag_WDTH-1:0]         I7dfe4eb1588a68b8a35dec39978d06eb;
wire [fgallag_WDTH-1:0]         I144843095a5e8952e26bb5c9943f0cad;
reg  [fgallag_WDTH-1:0]         I9d94ad2da06ac1fef4da7dcc56abffca;
wire [fgallag_WDTH-1:0]         Ica59cc444ecf8f8700bf1ce16a254b89;
wire [fgallag_WDTH-1:0]         I0b6cd5372e2cc6a72c1c8f984279cb69;
reg  [fgallag_WDTH-1:0]         I51262e3abe460148e3c2d2b74989c2b8;
wire [fgallag_WDTH-1:0]         I0d69f1eb92a8b30d86ffbe0c153197f2;
wire [fgallag_WDTH-1:0]         Icd143823913eb777c0cba42d8a5802e9;
reg  [fgallag_WDTH-1:0]         I560583680bb2f5a0b5ede42ceaafcf8b;
wire [fgallag_WDTH-1:0]         I5a48ea253b357c8e6441be01918bc57c;
wire [fgallag_WDTH-1:0]         I02a575305a6112f734bc3ebf6b883b90;
reg  [fgallag_WDTH-1:0]         I389f83346ffaffe8186fb0074d71f43c;
wire [fgallag_WDTH-1:0]         Ic3c81f609bf98f2ded891b55bacbd453;
wire [fgallag_WDTH-1:0]         I20f0ea42718bdd84caf3da4a1b32c5a1;
reg  [fgallag_WDTH-1:0]         Ie89c2a1b3943d12197bb972bd12595b0;
wire [fgallag_WDTH-1:0]         Ie38b3f5ad91f2c983d519c9b1200559c;
wire [fgallag_WDTH-1:0]         I11489ad40e6ff10933319784981fe59f;
reg  [fgallag_WDTH-1:0]         Ic7be56919976a2d1088114c21c3c1ffb;
wire [fgallag_WDTH-1:0]         I1e5e2679a0e75104cc0be107ecadd01c;
wire [fgallag_WDTH-1:0]         I10fe1f517735fad803f3d5d75fa3d406;
reg  [fgallag_WDTH-1:0]         Icb5dab0df062ab46bd3d1a73e85ef4c2;
wire [fgallag_WDTH-1:0]         I903e174feff2be7109cdb19fa15a63ec;
wire [fgallag_WDTH-1:0]         Ifed41503f4acb3625530d3c74b5ccb52;
reg  [fgallag_WDTH-1:0]         I27a568cfc2df13cf689d366a25e5d05f;
wire [fgallag_WDTH-1:0]         I6893d09bc4fca46b4ad33c42d1950790;
wire [fgallag_WDTH-1:0]         Ic9550361e9ae769b5095df4857041e60;
reg  [fgallag_WDTH-1:0]         Ia6688964078f1ea87b742352877aac45;
wire [fgallag_WDTH-1:0]         I4ec84e063fb84d278ae90b84751b1bcc;
wire [fgallag_WDTH-1:0]         I29cedb22eb565264529effcf107e167f;
reg  [fgallag_WDTH-1:0]         I180deab4fe0d03104cf2ee035f6a9b8c;
wire [fgallag_WDTH-1:0]         I33998829023b087dbfa2e568d77291b3;
wire [fgallag_WDTH-1:0]         I229b8819c94a612ca986936c96ffa9a9;
reg  [fgallag_WDTH-1:0]         Iff6cd034bb64d13c21910c11bd92266e;
wire [fgallag_WDTH-1:0]         I5bc68432bc0a9ea8cd024d7fc3d3fdc8;
wire [fgallag_WDTH-1:0]         I62c0db0621c1a71960770d14c332dc0d;
reg  [fgallag_WDTH-1:0]         I7c34057a77f2bdda93c422506959818d;
wire [fgallag_WDTH-1:0]         Ib84e5271ffa3584148ce87dcf2a4f2a2;
wire [fgallag_WDTH-1:0]         Id94e17f3fb5b4fe7a5fbe8e25d02ec27;
reg  [fgallag_WDTH-1:0]         I7ff7d3fd63fa67cd72d1591c1a373180;
wire [fgallag_WDTH-1:0]         Ib633998a5fd0df508b47ba9c2f7c390a;
wire [fgallag_WDTH-1:0]         I10cb83fe0a939bf2784eb93ca1d7b3c5;
reg  [fgallag_WDTH-1:0]         If910e75bf10cf02a5b414cbb4fad1304;
wire [fgallag_WDTH-1:0]         Ie36cfd3519810d325d5cdc5150380fe0;
wire [fgallag_WDTH-1:0]         I8f8b2e93ca65e789d13d66ecea733894;
reg  [fgallag_WDTH-1:0]         I266697a6eca2b73a76fd375a0ad72a05;
wire [fgallag_WDTH-1:0]         I6ac3755ff9de4d43d0493891b2a5758d;
wire [fgallag_WDTH-1:0]         I2527b288272a0ee2127436252a47a6aa;
reg  [fgallag_WDTH-1:0]         Iba188abd7715fcbdad3b1f3d985c6fc3;
wire [fgallag_WDTH-1:0]         I5f0212d2ffe8f85614891882390bbc25;
wire [fgallag_WDTH-1:0]         I743dd733d1c20868da7a802ea99b23bb;
reg  [fgallag_WDTH-1:0]         Ic60c640562e3e45c89a1de78af509b6a;
wire [fgallag_WDTH-1:0]         I1e009fcbec9031954637f055cb9cfe01;
wire [fgallag_WDTH-1:0]         I5dacf7fba8d457b393930fcc76135b39;
reg  [fgallag_WDTH-1:0]         I0456494b33e4ec852c123cb3003b9886;
wire [fgallag_WDTH-1:0]         Ia6caeb0fcc8e7486e4d55b72a0d499a5;
wire [fgallag_WDTH-1:0]         Ic50ab0fdec011923b02c0c0d717befa5;
reg  [fgallag_WDTH-1:0]         I2ed7c217fe3e21fcb27e04f68b95dd6b;
wire [fgallag_WDTH-1:0]         I631e31da7dccd5b9311a4fa73e6a0227;
wire [fgallag_WDTH-1:0]         I3afc7e76861fb1fa36291ac8d5508483;
reg  [fgallag_WDTH-1:0]         Ifda5780b42bf451a7ce834f17b3fdd20;
wire [fgallag_WDTH-1:0]         Ib152eea9af905931ab45c4f9d89fa50b;
wire [fgallag_WDTH-1:0]         I7c06d7efe631bc01f98ca137df06876e;
reg  [fgallag_WDTH-1:0]         Iadca92fd39d1fd6032feb8415ca5246f;
wire [fgallag_WDTH-1:0]         I94118c50e80e5fed4294d16358d41579;
wire [fgallag_WDTH-1:0]         Ifd5f5f8f7ac4238cdb3a5fb2e86eecad;
reg  [fgallag_WDTH-1:0]         I613453382f19dd7eb9bdf51e945a33b0;
wire [fgallag_WDTH-1:0]         I1269d97f8ab4f5dddc002acf38b4a189;
wire [fgallag_WDTH-1:0]         I17e9d58c80d0da6e6093836deecfa743;
reg  [fgallag_WDTH-1:0]         Ideafa683e6a3a38848fb8bee22eba11b;
wire [fgallag_WDTH-1:0]         I89a793ddaf4887ddb8dbaaba13225d08;
wire [fgallag_WDTH-1:0]         Icd18edbcc227111c037023bf2b57ee5a;
reg  [fgallag_WDTH-1:0]         Ie4226e7e17c7971f07aaf0cfaeae495a;
wire [fgallag_WDTH-1:0]         I2b4fe952791866aecbbbcf01257d527b;
wire [fgallag_WDTH-1:0]         Id22f8eb74ec1e8499e150278e438359d;
reg  [fgallag_WDTH-1:0]         Ifbbfa268bd4c31c7eed45cd43fe6a405;
wire [fgallag_WDTH-1:0]         I797321bb9e3c2d7d3727af9a4cf5418b;
wire [fgallag_WDTH-1:0]         Id10ed140128d500e98d984a15b479fb4;
reg  [fgallag_WDTH-1:0]         Ib2d99d95f7a31e4745211c5ff96f851c;
wire [fgallag_WDTH-1:0]         I5eeb78b1511aa7b76765d82328323a4c;
wire [fgallag_WDTH-1:0]         If89f8e436166d9beeca9937c45b2c7d5;
reg  [fgallag_WDTH-1:0]         I692c0a91b415b400a3640e2d9a40edad;
wire [fgallag_WDTH-1:0]         I55f8232fcfcb929a35717f724f44eb4c;
wire [fgallag_WDTH-1:0]         Idfd24573e271b5cdd6f051496cb6ba8f;
reg  [fgallag_WDTH-1:0]         If8c4dc70212e8873167e1cad8e8e5692;
wire [fgallag_WDTH-1:0]         I7a7705607e93fca1cf1e7b1c92c4e3cc;
wire [fgallag_WDTH-1:0]         I145c31d89636b936f18a19bf50966bbe;
reg  [fgallag_WDTH-1:0]         Ib2f75e91bf9e1d32a3f170fc85244139;
wire [fgallag_WDTH-1:0]         I7e2e0ffb2b5622ba6e03a47755a9a1dc;
wire [fgallag_WDTH-1:0]         I15cae93770d041e2ef681a81e8256059;
reg  [fgallag_WDTH-1:0]         I3606dc61f24567cb1ace443cea62a43b;
wire [fgallag_WDTH-1:0]         I5f50e835526833015a2087dbdb77686e;
wire [fgallag_WDTH-1:0]         I6a86457e1b16bfc515084fe599281818;
reg  [fgallag_WDTH-1:0]         Ie402c9f793b7306323efb8fe23533250;
wire [fgallag_WDTH-1:0]         I98f32439ec64d796ebb157815b259aa2;
wire [fgallag_WDTH-1:0]         I2453c39e5805313c3a8fd0d074058916;
reg  [fgallag_WDTH-1:0]         I54652565023310e2eccfc4cb87c56b43;
wire [fgallag_WDTH-1:0]         Id59ca1b1cff93a8544c54c6d4ee22b2f;
wire [fgallag_WDTH-1:0]         I34636cc42b16776295078bd349a76ac6;
reg  [fgallag_WDTH-1:0]         I616b7a5987edbc001e0ae1b638f25a39;
wire [fgallag_WDTH-1:0]         I726538434626c5202d53d29faedddd56;
wire [fgallag_WDTH-1:0]         I48f8d5589f772fbb4b3923fbd213e7f7;
reg  [fgallag_WDTH-1:0]         I06604bac478ee906b3fe8ff307cdf046;
wire [fgallag_WDTH-1:0]         I8ea236c734f7b96620a37750134d3872;
wire [fgallag_WDTH-1:0]         I83e4b71b0a0a3a82fc0a9fb56f803fa9;
reg  [fgallag_WDTH-1:0]         I135dd8a85aca863db660f2ad4f80ca2e;
wire [fgallag_WDTH-1:0]         I259d7244226dbcbd1d02df5ca164afdc;
wire [fgallag_WDTH-1:0]         I2abd0942d4d5e3aff2d24db9656c025f;
reg  [fgallag_WDTH-1:0]         I8715d73b58270dfa33b903e9cfb50be8;
wire [fgallag_WDTH-1:0]         I086375f289b769938edfc8b9b5146714;
wire [fgallag_WDTH-1:0]         I0fa19f52fef5a583890e3096eb23f1db;
reg  [fgallag_WDTH-1:0]         I7f60cb59895af6d314f5d0f401c80350;
wire [fgallag_WDTH-1:0]         Icb82f8092f14511d62f7cbe821af9faf;
wire [fgallag_WDTH-1:0]         I0e4a9bf26a9df3551a69edced6128e30;
reg  [fgallag_WDTH-1:0]         I3e25e6e9de5ee9242a472ce957056762;
wire [fgallag_WDTH-1:0]         I7e8df00362c29bd3924ecbe3dd1db23c;
wire [fgallag_WDTH-1:0]         Icd359ef9d3a983f4258cc4441110cc97;
reg  [fgallag_WDTH-1:0]         I4c5f36517aaf872e7f05de2f7f76a6ce;
wire [fgallag_WDTH-1:0]         If1014cbbd6e267aaacbcf3c8ba33a98b;
wire [fgallag_WDTH-1:0]         I31d6000373f248b1dde9fc0108bfd280;
reg  [fgallag_WDTH-1:0]         I0e993e6f98616632f17835a2994f45e3;
wire [fgallag_WDTH-1:0]         Iae4dfe3ede67923e8b740dd575b216b6;
wire [fgallag_WDTH-1:0]         I445cd3125f69b7e29d582a4803709c8f;
reg  [fgallag_WDTH-1:0]         I281f996740b16568b9d29ca41a3fa50d;
wire [fgallag_WDTH-1:0]         Iccfddf46ea48242ca751b5d53f98d270;
wire [fgallag_WDTH-1:0]         I2a8dcc8d3db0d8b5bb54bc7fae5e6ca7;
reg  [fgallag_WDTH-1:0]         I55bbb73d68871d9dbce4d590c029aeab;
wire [fgallag_WDTH-1:0]         I804705ac9a613b4107c8ceaac4127386;
wire [fgallag_WDTH-1:0]         Ibbf4549a33d4916489e7e325a811add1;
reg  [fgallag_WDTH-1:0]         Ida491561008f4984480d1b0f09d2fa77;
wire [fgallag_WDTH-1:0]         I8f40972503fbfdab92676a32f351dfe6;
wire [fgallag_WDTH-1:0]         I9a2d80bf2bbc2101c8e426cfc1c8277b;
reg  [fgallag_WDTH-1:0]         I624e237f248d292c0417ff85056857b0;
wire [fgallag_WDTH-1:0]         I8fc9ec077c7c6ce5e2660a4530a234ae;
wire [fgallag_WDTH-1:0]         I71c9904d29e88f0a5e6d7f8ec88de592;
reg  [fgallag_WDTH-1:0]         Ic7c1fd79ba76dbb254c6183017f40b3e;
wire [fgallag_WDTH-1:0]         I3e3bf3c2155f584784863ae41cb73c7d;
wire [fgallag_WDTH-1:0]         Ic6c8869890916818213809df90b52856;
reg  [fgallag_WDTH-1:0]         I546d683af76dc209a5205c6274abe908;
wire [fgallag_WDTH-1:0]         I9cc24d95a0ddbe4145d144003778eebc;
wire [fgallag_WDTH-1:0]         I3c61b092287e1f2c446aa7346b3dfcfb;
reg  [fgallag_WDTH-1:0]         I7b4bb785489c5bb22c84d9778192fe44;
wire [fgallag_WDTH-1:0]         Ib9b96de1e217660c2ac9f7815249c6a2;
wire [fgallag_WDTH-1:0]         I8f94e1fe9df14c5dd75421cdfe8b1efe;
reg  [fgallag_WDTH-1:0]         Ifc6af7d7aeb7162d554b8604a44f3361;
wire [fgallag_WDTH-1:0]         I2cc498e11d3d487d1e8319df8521ff6d;
wire [fgallag_WDTH-1:0]         Ie2a432bd8429925297936c8aebf7282f;
reg  [fgallag_WDTH-1:0]         I5b650c4c3291670b480a7f1095093dfb;
wire [fgallag_WDTH-1:0]         Iae3d8158d13c8179719cbe12fdd7f9ab;
wire [fgallag_WDTH-1:0]         I309c99cc023e0c7804b2574821d63f10;
reg  [fgallag_WDTH-1:0]         I2f5f88cb5e5e4723bd8a83c5fa80cc4c;
wire [fgallag_WDTH-1:0]         Ieadf1b0e427ecddd261297ae4054a0bd;
wire [fgallag_WDTH-1:0]         I5806c65240e9ce9f9d0804d063c2674e;
reg  [fgallag_WDTH-1:0]         Ic174b361182c98486e65b7f87b073274;
wire [fgallag_WDTH-1:0]         I8dbe4e03db655e1f691254835fb58798;
wire [fgallag_WDTH-1:0]         Ib73d05919f3373f122b121be5a038f4b;
reg  [fgallag_WDTH-1:0]         I7ba2f7201745258dbf224de087a25233;
wire [fgallag_WDTH-1:0]         I14b22818be28bc385f91920399012555;
wire [fgallag_WDTH-1:0]         I84136dfec9c8ab98228801deffbe8c19;
reg  [fgallag_WDTH-1:0]         I131a4bd335fc23ee10f7ccb1881ab9cd;
wire [fgallag_WDTH-1:0]         Id2878a17128a23eee2272c7e39743bd3;
wire [fgallag_WDTH-1:0]         I09e9850f90a7f073169e66c9e2339f51;
reg  [fgallag_WDTH-1:0]         I90cb3e06b42f25956b788a792eef371f;
wire [fgallag_WDTH-1:0]         I3701d2d2e74c43b3ae347902c0efff20;
wire [fgallag_WDTH-1:0]         I1260922a3e6cd464e43f215299d70ef1;
reg  [fgallag_WDTH-1:0]         I56302770a8d56932e7bb5dcff56c71e2;
wire [fgallag_WDTH-1:0]         Id6487b559b7ebad725aa43382f09bab3;
wire [fgallag_WDTH-1:0]         I97cf4612b19722d7f5f4cf9a867a9b22;
reg  [fgallag_WDTH-1:0]         Id3b8c058b3838c388eb5ddcb31dfc799;
wire [fgallag_WDTH-1:0]         Ib6ea830665d44628aef5041b2fa46328;
wire [fgallag_WDTH-1:0]         I4856ddf90e056e12eb6ec14d66f776b3;
reg  [fgallag_WDTH-1:0]         I7ca8ce63dfb821d10304958bada71737;
wire [fgallag_WDTH-1:0]         Ia6181e1acc2ea46a85626a22983e2662;
wire [fgallag_WDTH-1:0]         I370986beb4c411ce7154bb1c7045c5d8;
reg  [fgallag_WDTH-1:0]         I06ad44414b45d262f9542015d2dead8d;
wire [fgallag_WDTH-1:0]         I8b38fb1f95f036393933d07e0a60b875;
wire [fgallag_WDTH-1:0]         I0b22c5487df5e2b47d2ac3e16ca195b9;
reg  [fgallag_WDTH-1:0]         I833ef4acfed17e4699d65cbaa3e7dbd5;
wire [fgallag_WDTH-1:0]         I33d76ad1185bbf80de5e8ff0ad52b15f;
wire [fgallag_WDTH-1:0]         Ic7437fa32ca344b6eaa895d35d335e57;
reg  [fgallag_WDTH-1:0]         Ia77e3db939408af719e0a8555dcb68ed;
wire [fgallag_WDTH-1:0]         If2c522a90684b77b18f0058d1d2b14d8;
wire [fgallag_WDTH-1:0]         I1dcfffaaabc223ae08cd9d08d6e968d2;
reg  [fgallag_WDTH-1:0]         I57ab4999187992eda55a82bf0f09b31f;
wire [fgallag_WDTH-1:0]         I869e040de179572cdfd9373a4de8b31c;
wire [fgallag_WDTH-1:0]         I16bb10e8ddda86c2c8a1df7b0ec4c133;
reg  [fgallag_WDTH-1:0]         I21f7b5402ae8e8954d99931bd5108250;
wire [fgallag_WDTH-1:0]         I3fb8890ee1f1cb30ecdf50d69e4ac0fa;
wire [fgallag_WDTH-1:0]         I50ab3193dde101b550b508744be5a775;
reg  [fgallag_WDTH-1:0]         I3627708869b47d460182bc5040092f9a;
wire [fgallag_WDTH-1:0]         I6b60e2478c009889776de20209929ee0;
wire [fgallag_WDTH-1:0]         I022ed4e5e55e9c3cd418bca5475beb82;
reg  [fgallag_WDTH-1:0]         Ifd88f0f0abd1c037434dc16e34550d2a;
wire [fgallag_WDTH-1:0]         Ie6b559c2f0bd388d072b660341eebe31;
wire [fgallag_WDTH-1:0]         Ie44afe129f71022f34e9f9cb5ac4eb3d;
reg  [fgallag_WDTH-1:0]         I27eec53da48406e7e1202345a0810e08;
wire [fgallag_WDTH-1:0]         Ia46aa3a3e6a01d4690dfe0e7f1eab548;
wire [fgallag_WDTH-1:0]         I38c8f2c90a4d997e5597b462e7e8c613;
reg  [fgallag_WDTH-1:0]         I682d42afaaf103550ce4fbdba6192c88;
wire [fgallag_WDTH-1:0]         Idb7244908662bcd97fe8fe0db4b1abdc;
wire [fgallag_WDTH-1:0]         Ib38a5e546fdc5837a97c4ff3a627777d;
reg  [fgallag_WDTH-1:0]         If225534847db8723768941c3819ed7c0;
wire [fgallag_WDTH-1:0]         If570b3495ea5b3f250cf4873f5dd0bb9;
wire [fgallag_WDTH-1:0]         Iaebf3465f121a3c054c87227d7e9e167;
reg  [fgallag_WDTH-1:0]         I43a91b2232a47d1f6731bafc15ced5db;
wire [fgallag_WDTH-1:0]         I50bbcccc40af5e9700b97e682953c8c9;
wire [fgallag_WDTH-1:0]         I6fd1108c6ac90f5c69db5aca76055a32;
reg  [fgallag_WDTH-1:0]         Ic54026604afd19b0c7c71ea1ac0f1c4e;
wire [fgallag_WDTH-1:0]         I5422f11a7e0b646dd4fa254602f91b34;
wire [fgallag_WDTH-1:0]         If6f92d3b43974c88963a188a26bc3009;
reg  [fgallag_WDTH-1:0]         I218bd69f079aa21f0dda241ae6e387ad;
wire [fgallag_WDTH-1:0]         Ic5c34f86b03fffdcf723ff4116822e3f;
wire [fgallag_WDTH-1:0]         I19fb6cacc6841dec5653ef273676f18f;
reg  [fgallag_WDTH-1:0]         Iaaacca4d06ad0f202d839fd7674f1829;
wire [fgallag_WDTH-1:0]         I2ebd72fb063702a7c36b4b546f4b94b8;
wire [fgallag_WDTH-1:0]         Ia0abbf270f98b4bf4f29b56611db23b6;
reg  [fgallag_WDTH-1:0]         Iecddac410bb2121da0df2d73c2d23cb8;
wire [fgallag_WDTH-1:0]         I6328eca7325eea20ccf30adf8b928edb;
wire [fgallag_WDTH-1:0]         I38ad3c494c777f3985d61eef7cab8fb6;
reg  [fgallag_WDTH-1:0]         I1aabc0c0b7b602297ad592ae48b23452;
wire [fgallag_WDTH-1:0]         Ica13fd6daec896ddb0fa6be797edf6bb;
wire [fgallag_WDTH-1:0]         Ieb8d87fc8ecfad97cb9840b3739d6ea4;
reg  [fgallag_WDTH-1:0]         Ida3aaf7237b1383cfe95eeccf3971a8e;
wire [fgallag_WDTH-1:0]         I970c832cf68b5178f3d8111c9fed3b5a;
wire [fgallag_WDTH-1:0]         Ic1087bae156ef4dd5fe218537432b0ed;
reg  [fgallag_WDTH-1:0]         Idd2a8ed39edf6697b0988ee4eb4f2d95;
wire [fgallag_WDTH-1:0]         I65f78ccc122f96f97fee54955d370288;
wire [fgallag_WDTH-1:0]         I6655118cfe24b706e6557438ffa1711a;
reg  [fgallag_WDTH-1:0]         I735c660d5232e03dd8fb129e2ca4b445;
wire [fgallag_WDTH-1:0]         I5f77d7804a3e4adb641908be74f3ea19;
wire [fgallag_WDTH-1:0]         Ia12b8e62d6e1d52861589818deb6a851;
reg  [fgallag_WDTH-1:0]         Ia04d6065987df3f007658614406cbc28;
wire [fgallag_WDTH-1:0]         I9263e4ab78ca05f93ff921c4fd9ff787;
wire [fgallag_WDTH-1:0]         I59260857d96064096680b8361521b588;
reg  [fgallag_WDTH-1:0]         I7aeddde5b60828ac7f8b6c2addaf220b;
wire [fgallag_WDTH-1:0]         I6f8f253cfb1fe1c2254e557f732a9b22;
wire [fgallag_WDTH-1:0]         Iee39a5d6276b276729abd14472262ed1;
reg  [fgallag_WDTH-1:0]         I150c28296847348d69cce123f20656c3;
wire [fgallag_WDTH-1:0]         I3f247e74edd47e346d3bbb5dc3408844;
wire [fgallag_WDTH-1:0]         I20aa2879f47abd3c368f7494d944222d;
reg  [fgallag_WDTH-1:0]         Ib94d38d19b3791fa2d1b42fdfde8435e;
wire [fgallag_WDTH-1:0]         Ie0b33e2c1def11ccdaaae4ed2b042df6;
wire [fgallag_WDTH-1:0]         If0192b9580e5fdb8d71b422ccb28666f;
reg  [fgallag_WDTH-1:0]         I94865622898b2e481e86a244f7aa2759;
wire [fgallag_WDTH-1:0]         I39448514454c92ce93c3b0bc1d0e5d50;
wire [fgallag_WDTH-1:0]         I5095a3f4dd1c3bca218d17f5c609b667;
reg  [fgallag_WDTH-1:0]         I1a4a432e735367f515ca747cef7d7d04;
wire [fgallag_WDTH-1:0]         I677e9047c3ede581db9512b4fe072ea9;
wire [fgallag_WDTH-1:0]         Iea2a2368935757fe57b3d283fdccdb3e;
reg  [fgallag_WDTH-1:0]         Ib3a2b744d8f38671a63da6f8f8f1a6a1;
wire [fgallag_WDTH-1:0]         Ief6fbe6927f26b7a037f8e0bcb7751d8;
wire [fgallag_WDTH-1:0]         I36cd8882960099f242551ff3cbf8e4bd;
reg  [fgallag_WDTH-1:0]         I87716ad5a64592abb812ffe041ccc163;
wire [fgallag_WDTH-1:0]         Ie1e5c12afad8f2d8c2abef26473b7d9c;
wire [fgallag_WDTH-1:0]         I3ac47b1ac8e31b0082c7acfab65e222c;
reg  [fgallag_WDTH-1:0]         I71b259faefbea7ce8f47e0ffb556a0be;
wire [fgallag_WDTH-1:0]         Ic8f2ae80147ee27c548de195dfefa382;
wire [fgallag_WDTH-1:0]         I2a4914c71690073767e6f5fe13f26178;
reg  [fgallag_WDTH-1:0]         I2161b2ff3514dbdbb79d25da87eeec2b;
wire [fgallag_WDTH-1:0]         I533eb0729cc85339e2fcd1847930adc9;
wire [fgallag_WDTH-1:0]         I99903b3dad6af712c1148c2f43194da0;
reg  [fgallag_WDTH-1:0]         I860a3c9fca8d240c68ce3825192353b0;
wire [fgallag_WDTH-1:0]         Ic68fd0a9ea4b641913aadb7fe011d8ab;
wire [fgallag_WDTH-1:0]         Icccc370bf2f48ce93f479d13fa7075e9;
reg  [fgallag_WDTH-1:0]         Ie4eb18c7e906c9a25c12e9980a9f61cb;
wire [fgallag_WDTH-1:0]         Ica1f13759a67176573842e56bcdf09bd;
wire [fgallag_WDTH-1:0]         I5b5a0ccc2f5f9a7554d6d55b0dc61d76;
reg  [fgallag_WDTH-1:0]         I20a24846a74af76fa4470d6350546a9a;
wire [fgallag_WDTH-1:0]         Ifed30886099cbeb5da64d1d0696bb5de;
wire [fgallag_WDTH-1:0]         I0cd3d6b7cb85a87bfbebc1982c5fddf7;
reg  [fgallag_WDTH-1:0]         I90d40f6e9721a7d075512b8b81907453;
wire [fgallag_WDTH-1:0]         I317b34a0f6e16550b4a3e887cdd0c250;
wire [fgallag_WDTH-1:0]         I38a9b558c3289d954fe0de802b473be4;
reg  [fgallag_WDTH-1:0]         Ifc4525a25f38affb399004b057d1318c;
wire [fgallag_WDTH-1:0]         I39fa2bacef89a2f523f91b1e7f3cbe90;
wire [fgallag_WDTH-1:0]         Iacadd2fc2b7446edd7c45341a0670cb7;
reg  [fgallag_WDTH-1:0]         Icc93649a2050b9ded1e625be936b411f;
wire [fgallag_WDTH-1:0]         Id01272140c18ae29a8c75e493cf01268;
wire [fgallag_WDTH-1:0]         I316810ae743e5626556ad8f3176849bc;
reg  [fgallag_WDTH-1:0]         Ibcc30c960ae0f29c4efb1266c9e490ac;
wire [fgallag_WDTH-1:0]         I4d981fbbadbaa97ef98429ac12ca6710;
wire [fgallag_WDTH-1:0]         Ib9d5224a4d0b87aeb65cd6cf030ee52e;
reg  [fgallag_WDTH-1:0]         I3b2ffa79fd2227a24c6468a89f2bd989;
wire [fgallag_WDTH-1:0]         I2a1672224d3a3c513f2f04bb4dc123e0;
wire [fgallag_WDTH-1:0]         I92246b941db36e725ce7cbb1c9b4a0b5;
reg  [fgallag_WDTH-1:0]         Ib489a11dfdd8a2b3ad561c965b3d7d2a;
wire [fgallag_WDTH-1:0]         I364afb3546858e133a2bb541798e7886;
wire [fgallag_WDTH-1:0]         I62b8229b8e21a4bfd043c23450ff50e5;
reg  [fgallag_WDTH-1:0]         Ifa51cf9f9d3d1b91c72387f5daf05c79;
wire [fgallag_WDTH-1:0]         I9908671d65856b8714d43d83f0811a17;
wire [fgallag_WDTH-1:0]         I49266ae645036370bba4d99a1a85bc6f;
reg  [fgallag_WDTH-1:0]         Ifda20d77c574c8f13816620c56fff950;
wire [fgallag_WDTH-1:0]         I3e3f06cade9b6c8ea10e45996449e405;
wire [fgallag_WDTH-1:0]         I242c35248366a124753da854841595a7;
reg  [fgallag_WDTH-1:0]         I03ce0915d3a170429959221b6c8cd16c;
wire [fgallag_WDTH-1:0]         I9525b42d4dc80c42608cfa0ea10b8b2d;
wire [fgallag_WDTH-1:0]         I347dd57356eb6e025dada067d0f661b9;
reg  [fgallag_WDTH-1:0]         I9c2da511df8277b7e61cf8611d04dd32;
wire [fgallag_WDTH-1:0]         I94361c7eb9f16c4b20dfcdb7b8ad8cf3;
wire [fgallag_WDTH-1:0]         I6bb3031e93da171fac995de3e23c8b71;
reg  [fgallag_WDTH-1:0]         Ib8c628f3d97ffdf8a8b5db0fe90bbfa8;
wire [fgallag_WDTH-1:0]         Idc043493a919ec50417594df96f4d669;
wire [fgallag_WDTH-1:0]         I88cede4b89eb0f3917530d0ce2468c3a;
reg  [fgallag_WDTH-1:0]         I42e0e42ae26723497a1da5e86e855499;
wire [fgallag_WDTH-1:0]         I9e051ecfe79c36a913b15a0c7fe27f4d;
wire [fgallag_WDTH-1:0]         I3a590077bea5f1023ac006b321083554;
reg  [fgallag_WDTH-1:0]         Id7e44a94fcaa2ca22ac9eb6756ecb830;
wire [fgallag_WDTH-1:0]         I5479857f4f724aaea25ba124c9edb232;
wire [fgallag_WDTH-1:0]         I2bac571cd0d32e8a1bd527245a76f11b;
reg  [fgallag_WDTH-1:0]         Ie91db5e628b828dfaa8c1bd7d614d986;
wire [fgallag_WDTH-1:0]         Id2ed64cae3cb1e0ada8e3fb4ebb2dc78;
wire [fgallag_WDTH-1:0]         Ic1c911bc20d03275c7d20ab993e9a54d;
reg  [fgallag_WDTH-1:0]         I683ebfd7677d9e175d7a86479a5b42c6;
wire [fgallag_WDTH-1:0]         I16b9849d3f2edd7f9ed7accb138d2c02;
wire [fgallag_WDTH-1:0]         Iff207077a60c0196ac33f68e37d7d824;
reg  [fgallag_WDTH-1:0]         I11090ba16ce17a70438618b474837c33;
wire [fgallag_WDTH-1:0]         Ibcfe38455aa7aa33ae950172fb915dc5;
wire [fgallag_WDTH-1:0]         I0980811a7928bd72e415daf24b41137f;
reg  [fgallag_WDTH-1:0]         I845dd61995152e9d39cea7f0370b5a4d;
wire [fgallag_WDTH-1:0]         Ic9d9832294a3707b4041b2c4d8f92615;
wire [fgallag_WDTH-1:0]         Ie5a8e0e3d35d27fbb680552444f2ae65;
reg  [fgallag_WDTH-1:0]         Ia3e4dff8c98b38b6aebec9094ed26421;
wire [fgallag_WDTH-1:0]         I3ef9641c53e7aa6a588481b57b865aa3;
wire [fgallag_WDTH-1:0]         I91e4dd08f282857ab4c275bb1441c9d7;
reg  [fgallag_WDTH-1:0]         Id69a54dc4854348a482f052c64a736ca;
wire [fgallag_WDTH-1:0]         Ie838f76c6fc041e4fa66441094ae477c;
wire [fgallag_WDTH-1:0]         Iea26a1265fd6c48c038993b2038d2747;
reg  [fgallag_WDTH-1:0]         I0f56c52253603ac01a22f3b942429262;
wire [fgallag_WDTH-1:0]         Ice9f8149ed08f537da5e146b417085e0;
wire [fgallag_WDTH-1:0]         I7920256f397f35450287256339769d4b;
reg  [fgallag_WDTH-1:0]         I718f82404f82fe0e822ee20d33ad20a2;
wire [fgallag_WDTH-1:0]         I71f6bd2fe34731aab306cfb89a3335ca;
wire [fgallag_WDTH-1:0]         Ibad06757b56b14755f0e50620a53dc6c;
reg  [fgallag_WDTH-1:0]         I6c86073aaa32b64a43d06eb1a2d9fba8;
wire [fgallag_WDTH-1:0]         I5dd57cfd0d7ce83fcbdb3f560ac713fb;
wire [fgallag_WDTH-1:0]         Id76592cbf9ad537e9cab20469c5e5861;
reg  [fgallag_WDTH-1:0]         Ie0c8e27167e6ba97a83dd238086f45e6;
wire [fgallag_WDTH-1:0]         I239498228bdcb1c2a8b2cbef48e850a6;
wire [fgallag_WDTH-1:0]         Ibc80d98586cca13a6849ae053b68e5fb;
reg  [fgallag_WDTH-1:0]         I6bb5e8ee16a2bc0c3b77c882cfb659e7;
wire [fgallag_WDTH-1:0]         I82fc4233a3d2840670eb9b9adf6c9215;
wire [fgallag_WDTH-1:0]         I257237e7bef8b0e4cb27bc9a3a93aba6;
reg  [fgallag_WDTH-1:0]         Ieef625ad664ddadc849be46d1c083748;
wire [fgallag_WDTH-1:0]         Ieb08f6a94aa827632606608d014e26d3;
wire [fgallag_WDTH-1:0]         I1980cdd5ecb000134e55f507f369af66;
reg  [fgallag_WDTH-1:0]         Ice91b069200a91b2ad48fbf87bb2e766;
wire [fgallag_WDTH-1:0]         Ifdbb9947713ac574738236fcb5c6ae07;
wire [fgallag_WDTH-1:0]         Id0efde1d7f80f8848613c26fa4637c37;
reg  [fgallag_WDTH-1:0]         I9d4c7c85b4da5f7003ff05ed3a240a2e;
wire [fgallag_WDTH-1:0]         Ia737ee8f2c01feba1db87fe3e1a2388c;
wire [fgallag_WDTH-1:0]         I76952d4ed281844c1c1795290b1ddc05;
reg  [fgallag_WDTH-1:0]         Ia8f1616f8a65025446a5ab4cc1624f9b;
wire [fgallag_WDTH-1:0]         I5d8e065dba640832d9d8db3e4338fbb5;
wire [fgallag_WDTH-1:0]         I7fa89ba905b099ebafe001878c4f0bed;
reg  [fgallag_WDTH-1:0]         I29848deb21ad480cdf155d849dc7bd48;
wire [fgallag_WDTH-1:0]         I3b3e36ffb1cff2c07bc9a61afdde10c1;
wire [fgallag_WDTH-1:0]         Icd841b02588f755a3133b72f8c625897;
reg  [fgallag_WDTH-1:0]         I1ae69988f89b200bd0e48f640211321c;
wire [fgallag_WDTH-1:0]         I2c8137e5ee04a1067858d7bb8d09d65b;
wire [fgallag_WDTH-1:0]         I52945b9d986280c3dab4248e69247005;
reg  [fgallag_WDTH-1:0]         I7ddcc3c9f4d21aacc07d8eb285dee83e;
wire [fgallag_WDTH-1:0]         I38eb22d29ad9f4192499980fc17898b4;
wire [fgallag_WDTH-1:0]         Ia0319e76fc112b3457f20662a7a51603;
reg  [fgallag_WDTH-1:0]         I28f7cf50ea7ac81667ff1353e0e121bd;
wire [fgallag_WDTH-1:0]         Ib714941df0aaca40e7573e030d97b3f1;
wire [fgallag_WDTH-1:0]         I7a82bbf1146a3c68f01abf488a2e3c8f;
reg  [fgallag_WDTH-1:0]         I09b7dd699ae0c4d34a7d1588efc90452;
wire [fgallag_WDTH-1:0]         I47bcab5b082a8ce6312244224c162d39;
wire [fgallag_WDTH-1:0]         I05b26dca2316a9d527da24deb63c4756;
reg  [fgallag_WDTH-1:0]         Ic937101cc53e67403e56ac85011aa9ba;
wire [fgallag_WDTH-1:0]         I68ded74f52dbd02ceb1da62a79d619d2;
wire [fgallag_WDTH-1:0]         I256d84c23de18bd9a03cb41c0e3e4b8e;
reg  [fgallag_WDTH-1:0]         Ib42b03d2f76b8939ff3183008b17a969;
wire [fgallag_WDTH-1:0]         Iaa113fd5f1e0c51d9f47240fe81b5604;
wire [fgallag_WDTH-1:0]         I619aafd5767c45229765838152161b71;
reg  [fgallag_WDTH-1:0]         I4b99f00b1c2cdcee6bf4f1d2e8199ee4;
wire [fgallag_WDTH-1:0]         I907bf413f65fad54303751c054687b29;
wire [fgallag_WDTH-1:0]         I4bbb9f6eb1d79d41c7b5d61df854bd16;
reg  [fgallag_WDTH-1:0]         I01e153b020e1349eb66b47de581408df;
wire [fgallag_WDTH-1:0]         I7b727f2e9454f90d4fa4ef2cf69ddf23;
wire [fgallag_WDTH-1:0]         I997c88ff27fe957ec35a2b7146dd56f0;
reg  [fgallag_WDTH-1:0]         I8ca1a48206ed8f1dc7ca57d77d0331a2;
wire [fgallag_WDTH-1:0]         I6fc1f37134064dd7514b46ce7d27ceaa;
wire [fgallag_WDTH-1:0]         Ide7fdb7a17f3d99a7840a648e0873bec;
reg  [fgallag_WDTH-1:0]         I40e8430f50206db37e500c22f461b0c7;
wire [fgallag_WDTH-1:0]         I7856585e0374651fc5f9921f69706a0b;
wire [fgallag_WDTH-1:0]         I93dc025ca2d2cc3002c62c5d2e13d45b;
reg  [fgallag_WDTH-1:0]         I521128b7d945e025ded04037494c850a;
wire [fgallag_WDTH-1:0]         I79b1967c2128c611ee4fe0d14bced1f4;
wire [fgallag_WDTH-1:0]         I9c656300bb176deba4be8400371f0ef2;
reg  [fgallag_WDTH-1:0]         Ic24dbb1a30bb9a32c1992afcba90d4fb;
wire [fgallag_WDTH-1:0]         Ib8aeaf62789d1d7a5a23d7492ff551b2;
wire [fgallag_WDTH-1:0]         I141a53fdaada1994dc38d694fd03b5e3;
reg  [fgallag_WDTH-1:0]         I06cc903106b42e397fa7c4bc6c5edea4;
wire [fgallag_WDTH-1:0]         I9a8e8c3ce2c6323acee0877d445a2268;
wire [fgallag_WDTH-1:0]         I1d81174ecfb84b8c906126d13900178e;
reg  [fgallag_WDTH-1:0]         I765dff22de01d419a6626919d23850f2;
wire [fgallag_WDTH-1:0]         I701a3c05ad8e6ac5cea30b78707e77d1;
wire [fgallag_WDTH-1:0]         I92ab5c30a7bfae4e698a74d2e48cde1a;
reg  [fgallag_WDTH-1:0]         Ie9538b63a057a50371de2d17898d3ad7;
wire [fgallag_WDTH-1:0]         I75fefd09122859510021931c16051262;
wire [fgallag_WDTH-1:0]         Ifd41e7ed8ef5fa870c1abf043b5d5f2d;
reg  [fgallag_WDTH-1:0]         If93a5596528db9017b8783fa0cf1dbc2;
wire [fgallag_WDTH-1:0]         I2779af0ff280ea511af850df795d1fb6;
wire [fgallag_WDTH-1:0]         I983825ee77db3cbd86c937e5fe4707fd;
reg  [fgallag_WDTH-1:0]         I68016caaf170fbe2734c5b6aaf089894;
wire [fgallag_WDTH-1:0]         I2eb84b0b6b12b9269bb791ae03e5094d;
wire [fgallag_WDTH-1:0]         I715efc0ca41f678f8c582aaa3f255767;
reg  [fgallag_WDTH-1:0]         I169b0fac6d01a713986b636bf8dfc3fb;
wire [fgallag_WDTH-1:0]         Ie42cb87efb2b87d88eed6139132bb23e;
wire [fgallag_WDTH-1:0]         I764815deb8bceeb1b9929de2dfd46235;
reg  [fgallag_WDTH-1:0]         Iddb14d68b464d04fe9e0b4e62789601a;
wire [fgallag_WDTH-1:0]         Id2e2722999e300df1bc7ea89dbf5689d;
wire [fgallag_WDTH-1:0]         I1b869d6b94307bc9bea28db11161e61e;
reg  [fgallag_WDTH-1:0]         Ie5b71f77beb734a6ab7f7be6c6f9c252;
wire [fgallag_WDTH-1:0]         I2b7e1a65c52821f3f7e194a443b0117d;
wire [fgallag_WDTH-1:0]         Idf695c6735d8d8aafa37ad4cbd5a5872;
reg  [fgallag_WDTH-1:0]         I59f9fa0b81ca88915c338ece1d1e08d5;
wire [fgallag_WDTH-1:0]         I8b31aa4edbc800c99628c5851cad8770;
wire [fgallag_WDTH-1:0]         Ib9114ddde15c1908595081b52ba00c48;
reg  [fgallag_WDTH-1:0]         I4f27922ccb21b65dcfe2dc0fcc97cdf3;
wire [fgallag_WDTH-1:0]         Id40d461c28ecc2017d9b7d2eadf5ea44;
wire [fgallag_WDTH-1:0]         I3d52a609547a0ac3cd6d0481f09d00f2;
reg  [fgallag_WDTH-1:0]         Idd7ae55ba748fb36e49684037212936d;
wire [fgallag_WDTH-1:0]         I4b8f58440e6848610f2e7e06efbc64fe;
wire [fgallag_WDTH-1:0]         I45abcbcdc3951ebaef039e6cb2562d4d;
reg  [fgallag_WDTH-1:0]         Ib8da505d1572487e814e7b0682e6dfa9;
wire [fgallag_WDTH-1:0]         Ica1d5cc8dc277e91787ec1bf0f2ed65c;
wire [fgallag_WDTH-1:0]         I5bed8ad020614972a82bf3ad66300f12;
reg  [fgallag_WDTH-1:0]         Idedb59a6fa2f6ad049f81ac652c645d8;
wire [fgallag_WDTH-1:0]         Ie5d481ac7a371e1fd3c48c5cf9649a67;
wire [fgallag_WDTH-1:0]         Ic7ec84d03001998a8504a79afb1f0d5c;
reg  [fgallag_WDTH-1:0]         I7d50b49718ab2007accda67ac77a65d0;
wire [fgallag_WDTH-1:0]         I9786bf468ba8540d7e75d762fc832709;
wire [fgallag_WDTH-1:0]         I43cfed51e8dec917304dff4f44a984c6;
reg  [fgallag_WDTH-1:0]         I27e0600689451a7475a36143f0eb1079;
wire [fgallag_WDTH-1:0]         Ib093fabefab0a1b46d2199c1c948abc8;
wire [fgallag_WDTH-1:0]         If34baa3a92291d91308582e9c268ccaf;
reg  [fgallag_WDTH-1:0]         Iba6724b61ecb74552b9bb3cab96480c6;
wire [fgallag_WDTH-1:0]         I9b53bbb22003297175c6c4655ef83c93;
wire [fgallag_WDTH-1:0]         I8c00e1f1c7faa04600505a6f30e32ccc;
reg  [fgallag_WDTH-1:0]         I0abb44bd896fbc695e880fee67fb0c42;
wire [fgallag_WDTH-1:0]         I9df2a441fadba7dc49effc5eecf4b0e8;
wire [fgallag_WDTH-1:0]         I225a03b34b73fee071973985a66f9213;
reg  [fgallag_WDTH-1:0]         Ifd714548110aa979e735cc6e13d3ef57;
wire [fgallag_WDTH-1:0]         I102372ac8a06119e5d827d83f172bbd2;
wire [fgallag_WDTH-1:0]         I4b819b7da7ced2a32e77b3b26682168f;
reg  [fgallag_WDTH-1:0]         Ieeb6c7cdf1379ee3d2933d81bc812dbc;
wire [fgallag_WDTH-1:0]         I5cad4cd564b0956b08f22cd42d594b01;
wire [fgallag_WDTH-1:0]         I3d1050efa384172a3af1fa5f259a3877;
reg  [fgallag_WDTH-1:0]         Id682af5250edce8e3811d418ecf2dd10;
wire [fgallag_WDTH-1:0]         Id685ced1c37d97c75b49b2f790dbabad;
wire [fgallag_WDTH-1:0]         I66de52bc354a661ccda6f4d6d744bfdf;
reg  [fgallag_WDTH-1:0]         I1d02127e28fb2e9aaf352815627960e7;
wire [fgallag_WDTH-1:0]         I219e400c87948e7b2bf715745a4b152c;
wire [fgallag_WDTH-1:0]         Ib9a88f5ea722553569167ca7b186fd50;
reg  [fgallag_WDTH-1:0]         Ibee34260749dc92b8523e83cd64d6a40;
wire [fgallag_WDTH-1:0]         I3372567dacc350adf991928753209605;
wire [fgallag_WDTH-1:0]         I68904155ce7e8d722b67725f81af7f06;
reg  [fgallag_WDTH-1:0]         Ie9a2a59c7b3571194198dca0c679c5f6;
wire [fgallag_WDTH-1:0]         Ibf50476ac553bceaedcb121b28093394;
wire [fgallag_WDTH-1:0]         I7bc807d9f1b67d68e11c8a064b218963;
reg  [fgallag_WDTH-1:0]         Ie4b5a941feb385e88498a98e5f8ddc01;
wire [fgallag_WDTH-1:0]         I5d20fcccde5844e36b83d7fd7034c413;
wire [fgallag_WDTH-1:0]         Id1b5740fd8ce883d3cf724bd7410f27e;
reg  [fgallag_WDTH-1:0]         I30b2b34a0cecfdbdeecba5f286befccd;
wire [fgallag_WDTH-1:0]         I47e720341773b3a11f4c71b4e9644525;
wire [fgallag_WDTH-1:0]         I12c6efa1dbc88f222ebcb8866946eea1;
reg  [fgallag_WDTH-1:0]         I8ce739ddc344cacb2de7f2c88a882170;
wire [fgallag_WDTH-1:0]         I0251d8ecec82a24878ce494f0b417ce3;
wire [fgallag_WDTH-1:0]         I9c9d28abad8610fa2cecb74d18a1c9e3;
reg  [fgallag_WDTH-1:0]         I8b00260bb93e928e66e9d4aaeb0d9b55;
wire [fgallag_WDTH-1:0]         Ibeef795b2235c98439628da8d7c094e0;
wire [fgallag_WDTH-1:0]         I21af49923adfeca8b24188a7bba54b1d;
reg  [fgallag_WDTH-1:0]         I9c1ca916654bad308af37d040b486cf8;
wire [fgallag_WDTH-1:0]         I61769f7c08a0b9cf78068455410b6bb2;
wire [fgallag_WDTH-1:0]         I46c921b6dbb398813ad0d6c06e2eb33a;
reg  [fgallag_WDTH-1:0]         I05749703a8a131453c563ed2264680a7;
wire [fgallag_WDTH-1:0]         I77fe52c685b1075c294ac3c0a5b0d63a;
wire [fgallag_WDTH-1:0]         Ifa087dd71378f388142d351fa18806b5;
reg  [fgallag_WDTH-1:0]         I4b76fe5f9863a41733b76decf9867d16;
wire [fgallag_WDTH-1:0]         Ia688029a35b4a62417906c9aa1cd7719;
wire [fgallag_WDTH-1:0]         I3f3c345d02438bc96a1f7b162315ea43;
reg  [fgallag_WDTH-1:0]         I2805bb16fd574a64de548b39a532cd8a;
wire [fgallag_WDTH-1:0]         Ifaaab2c6f368b133936a7295eeb9b45d;
wire [fgallag_WDTH-1:0]         I7577c4409a32ebf50e5a187f71c84b1e;
reg  [fgallag_WDTH-1:0]         Ide6a696c06f17f455d56bb28cad98bd0;
wire [fgallag_WDTH-1:0]         Ifbe064ac0a5f4bbf6caae486064a983d;
wire [fgallag_WDTH-1:0]         Iec97b82162ff77d0b123feeb5b5904e6;
reg  [fgallag_WDTH-1:0]         I39bce1f71ede4663c187ddfd6501eda1;
wire [fgallag_WDTH-1:0]         I439ac39c831e0ca87a40f49e439ce24f;
wire [fgallag_WDTH-1:0]         I2206f864d477e44a18769ea9cc01d8ee;
reg  [fgallag_WDTH-1:0]         Id0e769bee61ae0a90c167fab061f5965;
wire [fgallag_WDTH-1:0]         I5c616021ebd98fc8e0fcf5b19732175c;
wire [fgallag_WDTH-1:0]         I9b67c7138cc6e8c9ef36b5cb28932c9e;
reg  [fgallag_WDTH-1:0]         I83e03af8657a4a237641a9da7922e502;
wire [fgallag_WDTH-1:0]         Id3a6c8114a92efaf5f6c280f897bef71;
wire [fgallag_WDTH-1:0]         Ic295c2717dcc256113776b8d39368802;
reg  [fgallag_WDTH-1:0]         I7565e071282ca6e77bb469afc522f1a2;
wire [fgallag_WDTH-1:0]         I854d4e2867b459da2e2fc06c438e6077;
wire [fgallag_WDTH-1:0]         I4875abaa409c919efee2cde0c90e1e7d;
reg  [fgallag_WDTH-1:0]         I5d0dc5d40385ab67bc7f540f212b6a97;
wire [fgallag_WDTH-1:0]         I3b334e8064cbfe97e70a0f4055496f04;
wire [fgallag_WDTH-1:0]         I0bcc0953acf369ba9571d11e68511af4;
reg  [fgallag_WDTH-1:0]         I548cac395730b8386670cc4c7a64319a;
wire [fgallag_WDTH-1:0]         Iff92d12470884efa033800c88e1983e3;
wire [fgallag_WDTH-1:0]         I4d92612c245b6ebb246d2f41b3dd4107;
reg  [fgallag_WDTH-1:0]         Ic6d9bbbfb7890540edd10aa5758b0c4b;
wire [fgallag_WDTH-1:0]         I3d167f5af41902dc0a6477d55cf0abfd;
wire [fgallag_WDTH-1:0]         I53a8be01a8f8067f67e0498c48cfa2a8;
reg  [fgallag_WDTH-1:0]         I7beb1f915a881a302f93c869d81417d1;
wire [fgallag_WDTH-1:0]         Iaa7edba3767735cad1ec76479b5548b0;
wire [fgallag_WDTH-1:0]         I036d8ab76c1f8c3b52ddcad50c6c8a6c;
reg  [fgallag_WDTH-1:0]         I5fc389bbc1ce31f7b326da719dc576d4;
wire [fgallag_WDTH-1:0]         Ifaa7aff0fb2af9d3e04b2641b13cf884;
wire [fgallag_WDTH-1:0]         Idaffa51af26a79990b50e9422da6074c;
reg  [fgallag_WDTH-1:0]         I922e6f05f7c6e0f6f0b1a5c9548df238;
wire [fgallag_WDTH-1:0]         Ia78b9e9a1faddb38b4a1472f5eea3939;
wire [fgallag_WDTH-1:0]         Ia17748dd92434f8658e49a3f7ed682e8;
reg  [fgallag_WDTH-1:0]         I8c6bb234a1ca3deba637adf746672194;
wire [fgallag_WDTH-1:0]         I367d25430d8ec417123931f9534f3eba;
wire [fgallag_WDTH-1:0]         I1ecdfded32659bd57c752928f0cc12eb;
reg  [fgallag_WDTH-1:0]         Ide24ebd7423d4c4f43577b019f2e30e4;
wire [fgallag_WDTH-1:0]         I38a19bd51c6ee4fcb38493d869b7808a;
wire [fgallag_WDTH-1:0]         If7bcd20651da485996362af6b633fec3;
reg  [fgallag_WDTH-1:0]         Ifc412122eab7560c9021a17d7f8700c4;
wire [fgallag_WDTH-1:0]         I0fe662c7d5cce9cf3cac56b6125852ff;
wire [fgallag_WDTH-1:0]         I7a04a2c4768a6703cb98c2adfd53088f;
reg  [fgallag_WDTH-1:0]         Ia5a56ed2c6b98e72002c6c5f946e7264;
wire [fgallag_WDTH-1:0]         I6867bb41ee0a7f4c6ae0071e7975526d;
wire [fgallag_WDTH-1:0]         Iebc9456956b29940df3df4dddae0619f;
reg  [fgallag_WDTH-1:0]         Ia888ed8885f66084b777f66e25cef1e7;
wire [fgallag_WDTH-1:0]         I74d3dc7b6116f47b27dbfd112d7afd5d;
wire [fgallag_WDTH-1:0]         Iefb9092502c1c93656c9050bf74e6849;
reg  [fgallag_WDTH-1:0]         I248229aecef00b87a70ce88920e407f5;
wire [fgallag_WDTH-1:0]         I13440021cb8441969d3242de4fc6a0b5;
wire [fgallag_WDTH-1:0]         I42edf14a24cb1e19924e0f5531f97ed9;
reg  [fgallag_WDTH-1:0]         I3d162a0ec918f220a7d5f4efdf89cb58;
wire [fgallag_WDTH-1:0]         Id3c71879c307df1390bbc60c55a5f249;
wire [fgallag_WDTH-1:0]         Ia332b7b61c57cee58ef4a1733da2afc6;
reg  [fgallag_WDTH-1:0]         I1ca0372f60e48f2f803778c9017023c0;
wire [fgallag_WDTH-1:0]         I2e1fa8e49bf48184e6a669d18f5c8ced;
wire [fgallag_WDTH-1:0]         Ib4450f5e900229ff87baede34be883b4;
reg  [fgallag_WDTH-1:0]         Ieb9693d54f0808b0ba463fd3c316a80e;
wire [fgallag_WDTH-1:0]         Ibc9c9339a0bcbc6addcce833051a8cd0;
wire [fgallag_WDTH-1:0]         Ie7d8f527db720e17a73a57400a5360a5;
reg  [fgallag_WDTH-1:0]         I63da03315d7e51fcacb0bc0298e506ed;
wire [fgallag_WDTH-1:0]         I2c0a2ad9eef6e84c60d1a6503aa836db;
wire [fgallag_WDTH-1:0]         I7c420e9724fd4bc31071a57ac1ba5293;
reg  [fgallag_WDTH-1:0]         I918f5a12e96bb96941f019940f27a5be;
wire [fgallag_WDTH-1:0]         I3b06c3a23b2068e8f45870524c4af870;
wire [fgallag_WDTH-1:0]         I5a38174a83eaebe2678ca70fe5915c02;
reg  [fgallag_WDTH-1:0]         Ib4fb115f442ff544fa3d21b4e9d3f075;
wire [fgallag_WDTH-1:0]         I87d44c01b261e9c13add415e6b3cc5ba;
wire [fgallag_WDTH-1:0]         Ib3639c700fe97648415fd4dfc8a6466b;
reg  [fgallag_WDTH-1:0]         I387403482432a3196109484d1120d584;
wire [fgallag_WDTH-1:0]         Ifc15e0dd91741676f23cc20fc542ec14;
wire [fgallag_WDTH-1:0]         I5228b59565a0ae5f56237e5332ddefa1;
reg  [fgallag_WDTH-1:0]         I619af17eaa4a56726d6ab322a74dd0a4;
wire [fgallag_WDTH-1:0]         I50fdfffb4e2dbcf33282b3653f595ad0;
wire [fgallag_WDTH-1:0]         I87188c070d52012c107a5b37e718a5d4;
reg  [fgallag_WDTH-1:0]         I7a67ed3bb370520d0d25ce407ab8cd8b;
wire [fgallag_WDTH-1:0]         I4e9786ec39d388cdce110c86bb436ae3;
wire [fgallag_WDTH-1:0]         I7d0ebb3f7a7e77362b41f9ec9b98c9af;
reg  [fgallag_WDTH-1:0]         I7629b35ca548190a81021a2c13d8919b;
wire [fgallag_WDTH-1:0]         I47cb30eb341ae7ce99042a16cd109f26;
wire [fgallag_WDTH-1:0]         I1c2e01ba53fb12e4c3e44e4a9ef97888;
reg  [fgallag_WDTH-1:0]         I004851d3828f135ebe4d2e6ab83936bf;
wire [fgallag_WDTH-1:0]         If004fa1c4e6bbe1f458c2d2a4f1f6e03;
wire [fgallag_WDTH-1:0]         Icf7e609c4a537e6f2a7b86b7035717d3;
reg  [fgallag_WDTH-1:0]         I0e2c382b2e62ed43b76697230e34b719;
wire [fgallag_WDTH-1:0]         I7c9910ade59c54e170c4f10822b5aff4;
wire [fgallag_WDTH-1:0]         I39d74e21fb67539c0d310571b99a3e22;
reg  [fgallag_WDTH-1:0]         I36dac27d10701db70fb2b5996a3f038f;
wire [fgallag_WDTH-1:0]         I98939499dd98e583a4788cacc66c7fc4;
wire [fgallag_WDTH-1:0]         I395b85e88acd203dd93e519710aea79b;
reg  [fgallag_WDTH-1:0]         I51d62ebd160eb0d073a7efb64d20079a;
wire [fgallag_WDTH-1:0]         Ic530781e13180026815873e12550e405;
wire [fgallag_WDTH-1:0]         I850e5fd50416aaad26283152c4a49ddc;
reg  [fgallag_WDTH-1:0]         Ib3545a88d68631af1c94ca2cb1f379af;
wire [fgallag_WDTH-1:0]         Iba43927cdbcb6a80953fced163686073;
wire [fgallag_WDTH-1:0]         Ide38f5cac19b1bc82b26bfa12e5f9d8c;
reg  [fgallag_WDTH-1:0]         I81ad7b044118734f4dc32a1a4e8eba31;
wire [fgallag_WDTH-1:0]         I29aefee3f95a7d2838ec5068515f69b0;
wire [fgallag_WDTH-1:0]         Ib2d8874232a27b78a8c664e0fa2af512;
reg  [fgallag_WDTH-1:0]         I5ad8c235d46349b6d310d0f175f84288;
wire [fgallag_WDTH-1:0]         Ib964c4dd0a0ce2553766251b73018699;
wire [fgallag_WDTH-1:0]         Id002a482b2a09d2d17b9fa903882e8e0;
reg  [fgallag_WDTH-1:0]         Ibc00920378e2427df2a63a47dc3eaded;
wire [fgallag_WDTH-1:0]         Ifd870cf74e7e3e5b348ad55af7242c27;
wire [fgallag_WDTH-1:0]         I359451948e89283ee89d89cebf689445;
reg  [fgallag_WDTH-1:0]         Ic5195bbaa69d95059cca6e152dc9f705;
wire [fgallag_WDTH-1:0]         Ic4ba744721cdd747affca302b2b926d4;
wire [fgallag_WDTH-1:0]         Ifffc8f779e22eedf06f7d1c24da411cb;
reg  [fgallag_WDTH-1:0]         Ia01f20e0bcf35c2ee4963e9c392c1004;
wire [fgallag_WDTH-1:0]         Id381e35622a3ac2c549a8c9b702ec020;
wire [fgallag_WDTH-1:0]         I3ccf7fbf7a13aef5daa7905b485d6e3a;
reg  [fgallag_WDTH-1:0]         I9f6f48fea88d1cd73ef2b24c7e819964;
wire [fgallag_WDTH-1:0]         If49e3943165e2782c928a7da86847145;
wire [fgallag_WDTH-1:0]         I9deead4d27ef61f468a1bac90adfa27e;
reg  [fgallag_WDTH-1:0]         I847feea780cc8a06caea2d2ea79ad281;
wire [fgallag_WDTH-1:0]         Ie4d85aa4951d1a918d698c9e411b1ab2;
wire [fgallag_WDTH-1:0]         I6c050a19b5031493dcc7163509b00012;
reg  [fgallag_WDTH-1:0]         I7ef6f4aeda7fd6775839c068c681f9bc;
wire [fgallag_WDTH-1:0]         Iff6a8d4bc8f5f37d0ccc2d41f469ca86;
wire [fgallag_WDTH-1:0]         If74b57fb1d88f063bfef26ae6b74ff2d;
reg  [fgallag_WDTH-1:0]         I0645e741da20a4957747188273a655b1;
wire [fgallag_WDTH-1:0]         I6bed9b6e8b499c11d719f869467d2322;
wire [fgallag_WDTH-1:0]         I9fc7952b3920da1adf39777e9a1cd13f;
reg  [fgallag_WDTH-1:0]         I71125dffdd2d37e44dbb46143c1e8d9a;
wire [fgallag_WDTH-1:0]         Id1db54a136ab42fe675fa77b2b7fd2de;
wire [fgallag_WDTH-1:0]         Ic013de8383ced83cb6cb368e54cd0f43;
reg  [fgallag_WDTH-1:0]         I50c166f958b22ce866cd40334918274c;
wire [fgallag_WDTH-1:0]         Ia6ed9442d22d3228ce14749ffdacfab2;
wire [fgallag_WDTH-1:0]         If71eac564bbca0cf2967a8803a24f586;
reg  [fgallag_WDTH-1:0]         Icd225144fd331b870847044b4d02bed0;
wire [fgallag_WDTH-1:0]         I32e0c22a86e88cadc6a956c213ff992c;
wire [fgallag_WDTH-1:0]         Ib19bf2920a5486af62d38fa181293a47;
reg  [fgallag_WDTH-1:0]         I5e876482090ce6007c2a2f2101c24654;
wire [fgallag_WDTH-1:0]         I1b0dcddcb3e0a398857f038d3a52e719;
wire [fgallag_WDTH-1:0]         I92a94b468b025e5c1d103b2f8c92709e;
reg  [fgallag_WDTH-1:0]         I026ded06f56d9ca93f47fd85aec4f7ad;
wire [fgallag_WDTH-1:0]         I8c6bcabb8814607901102aca5f820293;
wire [fgallag_WDTH-1:0]         I76fe38786c53eb9f57d6512adb920d5b;
reg  [fgallag_WDTH-1:0]         Iec596e94ec168a564bccbbaa7df833c9;
wire [fgallag_WDTH-1:0]         I731089de22b5becf3621097ed7a81b7e;
wire [fgallag_WDTH-1:0]         I7878eb8ad885ea4193b8534015a445bb;
reg  [fgallag_WDTH-1:0]         Ib514e01c261e43a725582a10596eed32;
wire [fgallag_WDTH-1:0]         Ifb3674681315fa8cf6739996b823a7aa;
wire [fgallag_WDTH-1:0]         I5b26270d07cd79afa7019dac72898e3c;
reg  [fgallag_WDTH-1:0]         Ic19a62cdecb2329370f7e11c48d3738d;
wire [fgallag_WDTH-1:0]         I2d5ef5bf9c28065a2a4ab718fbc8ba3e;
wire [fgallag_WDTH-1:0]         I167dccb5e632afc0686602b35f9dea42;
reg  [fgallag_WDTH-1:0]         Ib2f5691baa59adfbaad62f6ffc71fb05;
wire [fgallag_WDTH-1:0]         I7c5f9c301a0bdbf642f7b3f33e9bfc66;
wire [fgallag_WDTH-1:0]         I3cb81e29fa5d50fadebe311acca6d090;
reg  [fgallag_WDTH-1:0]         I9bdfaca6112385deb86e24ad7e45bbaa;
wire [fgallag_WDTH-1:0]         I7bde3bcef8556c1b1e4c7d2192196e00;
wire [fgallag_WDTH-1:0]         Ia25c11794a51c0937e0600032133a6dd;
reg  [fgallag_WDTH-1:0]         I0e647bb8351cfe7828423e7099525585;
wire [fgallag_WDTH-1:0]         Id13f3a39b334d8a80b7c8286b09bd1e1;
wire [fgallag_WDTH-1:0]         I95b38f00928726b7b701405baf74f66a;
reg  [fgallag_WDTH-1:0]         I185b758fb3e50bcfb1464fe2ab593cfe;
wire [fgallag_WDTH-1:0]         Ie6443f42260e0a2983927d0940c82a06;
wire [fgallag_WDTH-1:0]         I32c90cfef12eece5e90200ef79c7231f;
reg  [fgallag_WDTH-1:0]         Ie25e944f9e3100c39b69bb38dffca177;
wire [fgallag_WDTH-1:0]         I43003b2ef41b34363169f004a6668a59;
wire [fgallag_WDTH-1:0]         I0b27fcbbc4514fa212fe3d023bdb526c;
reg  [fgallag_WDTH-1:0]         I8e77032a54376578b3d16799e30c97f7;
wire [fgallag_WDTH-1:0]         Ic385923d90d69cd387eb9fb5f62fd9ba;
wire [fgallag_WDTH-1:0]         Ic420c6e4d3748dafd05197706f316f62;
reg  [fgallag_WDTH-1:0]         I4cd2a7f8f8ec378200b00d03e447ac92;
wire [fgallag_WDTH-1:0]         I2f642acd0cb0bd30177bc0d65751ed99;
wire [fgallag_WDTH-1:0]         Ifd760e2ecefe198d6f583146e8cbe9fc;
reg  [fgallag_WDTH-1:0]         I1b3c55aca0da232cf3f81d6d0914729f;
wire [fgallag_WDTH-1:0]         If1064670adff5b00cbf7809e2621cfd5;
wire [fgallag_WDTH-1:0]         I8078293bd2540592bffc91383fa5ad38;
reg  [fgallag_WDTH-1:0]         I34c76f1a126120c4474e750e9b51e034;
wire [fgallag_WDTH-1:0]         I72311a2c7557be2b6cb95b3bc6f511a5;
wire [fgallag_WDTH-1:0]         I1c0777b46bd3a7e2126f614d55703204;
reg  [fgallag_WDTH-1:0]         I0edb624c344787066a2267757052196b;
wire [fgallag_WDTH-1:0]         I79ee4c7277f713aa710ae8cf7c470aa1;
wire [fgallag_WDTH-1:0]         I2a719cff60bf0985e451a32aa71c82fe;
reg  [fgallag_WDTH-1:0]         Ia8443f199838742595ac114f35c00143;
wire [fgallag_WDTH-1:0]         I32bfef7a7ecaa533e3bf92fb560e657b;
wire [fgallag_WDTH-1:0]         Ia1af17b99a087b22fecb7ff79a370363;
reg  [fgallag_WDTH-1:0]         Ib25b8a538c9d64880e114bf4a80ca42e;
wire [fgallag_WDTH-1:0]         If4a6b6a8b44d2c55c93b111d20525ec6;
wire [fgallag_WDTH-1:0]         Id75247b073a7993bff1992cfe1874ff6;
reg  [fgallag_WDTH-1:0]         I25f6a3d7bb869082e4dbbd0ee8574c95;
wire [fgallag_WDTH-1:0]         I7d41f27ff64d549b7e5df6b172969d8a;
wire [fgallag_WDTH-1:0]         I63a6ad22f067ea29cf79e51ebc011f8d;
reg  [fgallag_WDTH-1:0]         If96057023747a1538d9f06966af48bc2;
wire [fgallag_WDTH-1:0]         Ie3a2d4d85d4e4ac011887cbd329bd9b7;
wire [fgallag_WDTH-1:0]         Ic3b5918c230369180edc94c5b01046e7;
reg  [fgallag_WDTH-1:0]         I199e995390462e06853b1f5cdbd46e0a;
wire [fgallag_WDTH-1:0]         I3bc9fcec69ab6a1efb2d86e03804415c;
wire [fgallag_WDTH-1:0]         Ifdf2c8ac7eb668b49ed3cf950d08c179;
reg  [fgallag_WDTH-1:0]         Iec6325d585ddd0a9f86bb5cd0229960d;
wire [fgallag_WDTH-1:0]         I9ee16e46a399d1445fcdf251757a5e43;
wire [fgallag_WDTH-1:0]         I644ff86dfecc5a20a1431f9cc67ee6f9;
reg  [fgallag_WDTH-1:0]         I4be1ccfec148a522fbf5b8375245cbb3;
wire [fgallag_WDTH-1:0]         I45cf986a60a429a68051f76beb8188fb;
wire [fgallag_WDTH-1:0]         I56a7bd438035251cd67dfb97b3a345d7;
reg  [fgallag_WDTH-1:0]         I074386ff6a3d8d644f4b2501c69f26c7;
wire [fgallag_WDTH-1:0]         I4e48461fcd58a133a09d856852887a4f;
wire [fgallag_WDTH-1:0]         I00c294596fc87af7f1b8377260232832;
reg  [fgallag_WDTH-1:0]         I83b378e5534c553b57beb22c5178a3ce;
wire [fgallag_WDTH-1:0]         I901714025da5b89ee929ea2859f3e6c7;
wire [fgallag_WDTH-1:0]         I7af09468b60d8e594a1aa85ad74911d5;
reg  [fgallag_WDTH-1:0]         I14f79d67f75af6a495d6eb2986210cda;
wire [fgallag_WDTH-1:0]         I976786b0539b07b056dad0f050eeb53f;
wire [fgallag_WDTH-1:0]         Ic0ed40d42c2af78809ecb381660ef229;
reg  [fgallag_WDTH-1:0]         Iacd805413ec1eb001b3083554f187554;
wire [fgallag_WDTH-1:0]         I8e1ad4f44dcac3e770dd862413b25a4e;
wire [fgallag_WDTH-1:0]         Ie03547bf9963c8a716e20e4aaef52dc7;
reg  [fgallag_WDTH-1:0]         I3e61e09fcc81a0011a79f5c5ce77bc46;
wire [fgallag_WDTH-1:0]         Iaf5caa6558f0a98b91fb72db734bbec4;
wire [fgallag_WDTH-1:0]         I26e996666f3436cfa998f34c3a05f7db;
reg  [fgallag_WDTH-1:0]         I6e6cbb7dba8eb3c02b5b4e4469e23cea;
wire [fgallag_WDTH-1:0]         I7b37d3b1b23f09c6ac46a94cf2c4ead7;
wire [fgallag_WDTH-1:0]         Idfc51f66e038c5ae625e98b615a7beaf;
reg  [fgallag_WDTH-1:0]         I8b25822c33f7d506ef69216af3fdab44;
wire [fgallag_WDTH-1:0]         Ief8b577d924f257ae5e1dd47009b0db2;
wire [fgallag_WDTH-1:0]         Idedf5a83a99278f57c6c9294b66b69eb;
reg  [fgallag_WDTH-1:0]         I06fd642cbc8aa2f65197801d7459cfa2;
wire [fgallag_WDTH-1:0]         Ie59366fcd6132a48f3e9be1bb5b600c6;
wire [fgallag_WDTH-1:0]         Idf55d61336e413c5aa3226b3b44f27b1;
reg  [fgallag_WDTH-1:0]         I22202e6c3de9b06c04ce9514af28933e;
wire [fgallag_WDTH-1:0]         I273c1e28c3ed897b7d0f6b36a3a8def9;
wire [fgallag_WDTH-1:0]         I05ce5256e568621df7129058c50e9fa6;
reg  [fgallag_WDTH-1:0]         Ib991cdbb91133cb82e154c575e00a174;
wire [fgallag_WDTH-1:0]         I64b507fe58b933919d0766631985a74e;
wire [fgallag_WDTH-1:0]         Ib8af108fab1636823714995f78c9d575;
reg  [fgallag_WDTH-1:0]         I5590364df6874420e169aa444ab520b9;
wire [fgallag_WDTH-1:0]         I7c0376cbc3660f3d82a5da22806ef5e3;
wire [fgallag_WDTH-1:0]         I166d54ee9aa9002c59a0aca2834632f5;
reg  [fgallag_WDTH-1:0]         I43a9e393037fb4aa84741dca22648459;
wire [fgallag_WDTH-1:0]         I3884d561185660e7e0f461b3487fdfd4;
wire [fgallag_WDTH-1:0]         Ib5f971498046dd212d853ff440c553cc;
reg  [fgallag_WDTH-1:0]         Ibb4d8301d90c66fdfac92b3fbc53c019;
wire [fgallag_WDTH-1:0]         I4b991f90354e3f74d105a64929a97d6f;
wire [fgallag_WDTH-1:0]         I325d401c6a1f445dcb7a83d90d2da75e;
reg  [fgallag_WDTH-1:0]         Ibae217fa4b808e4accbeb8f4a9a976ab;
wire [fgallag_WDTH-1:0]         I9534939768f7d2532ca4e6757dfafb72;
wire [fgallag_WDTH-1:0]         I91eeb6252974a1f69908b7e7114b95f5;
reg  [fgallag_WDTH-1:0]         Ia8bd7a3594f7084a57e64da023bf784c;
wire [fgallag_WDTH-1:0]         I090228a60e5919fa88d842b1638ee296;
wire [fgallag_WDTH-1:0]         I898cf70b6c6b57d256490f44d257fd84;
reg  [fgallag_WDTH-1:0]         I3ce4b9d41f5472bf60ed2802a2ab10eb;
wire [fgallag_WDTH-1:0]         I8994d511d611a3c1b7a8122cd3d2825e;
wire [fgallag_WDTH-1:0]         I256f73600515ae5c410454c425b66696;
reg  [fgallag_WDTH-1:0]         I93ec9bc6fbd056e7e52496546493e727;
wire [fgallag_WDTH-1:0]         I43d14ec8853bfd211aa6b887c7ebdd5a;
wire [fgallag_WDTH-1:0]         I362d1818937fd8d777531b85e86b4145;
reg  [fgallag_WDTH-1:0]         I2374b90dde1cf481baa40af31e1a43e3;
wire [fgallag_WDTH-1:0]         Icd810cceba64ffbb087600155338911c;
wire [fgallag_WDTH-1:0]         I21dda2280e7aa79b6abd7820829583e1;
reg  [fgallag_WDTH-1:0]         I0cee595f488a909ade8a3b4c90dbb0c7;
wire [fgallag_WDTH-1:0]         I33ddd4cdef0a0704f204f4fdb14fd859;
wire [fgallag_WDTH-1:0]         I94a6499c7bd1d40e4f363a58db1aa114;
reg  [fgallag_WDTH-1:0]         Iba4c3d91d492b000ab1de7add9f171a9;
wire [fgallag_WDTH-1:0]         I0c87f78f08ac77246d7b3b8604dfd700;
wire [fgallag_WDTH-1:0]         Ifb6f3d60109d87ffd54e72b3958c7e80;
reg  [fgallag_WDTH-1:0]         I2b4152aa4c51cc1c1ffabac78cea267c;
wire [fgallag_WDTH-1:0]         I54745c58c61eba829e4717cd842d519d;
wire [fgallag_WDTH-1:0]         Ia3fca25225f6cd049ec92b44cdb57049;
reg  [fgallag_WDTH-1:0]         Ie4c3dd5c191aff00a6d62006223c2b76;
wire [fgallag_WDTH-1:0]         I9e278d7b6cccaa39163d0867427709ed;
wire [fgallag_WDTH-1:0]         Iefa9788b8791b23ea0ca3d756d7e4019;
reg  [fgallag_WDTH-1:0]         Ie4c0ba9510f9b924999bb5f432137271;
wire [fgallag_WDTH-1:0]         I3e5d8af6fed6b47aebf2eef7010afa8b;
wire [fgallag_WDTH-1:0]         I2b790f210029547ce774150b5390eb12;
reg  [fgallag_WDTH-1:0]         I5bad544a17b384973d5672acbe0ac0d5;
wire [fgallag_WDTH-1:0]         Ie96538fd32c8f8d7a3144012d10b29a5;
wire [fgallag_WDTH-1:0]         I5c474a60ee2779b8f1477d07f4ca88d1;
reg  [fgallag_WDTH-1:0]         I231bfb8e19e1d9c4bbd29a0bd75c1ed3;
wire [fgallag_WDTH-1:0]         I050a226112c903de442358e2d5be8274;
wire [fgallag_WDTH-1:0]         Ie542464c6c79a43b078a8314c4def3b6;
reg  [fgallag_WDTH-1:0]         I1ecf87e33de04d02db9e64590bcaffde;
wire [fgallag_WDTH-1:0]         I4df410c6a7eea67fd73cc33c791e7aa0;
wire [fgallag_WDTH-1:0]         I0ae4560405030e9485f14f6eca025625;
reg  [fgallag_WDTH-1:0]         I60c97bf58193f004e3fcfdbd6a03ce6e;
wire [fgallag_WDTH-1:0]         Id7e318f124e0534c8e0538f99616ed01;
wire [fgallag_WDTH-1:0]         Ic14dfb6df2b9a62e5c9471684c0cb07f;
reg  [fgallag_WDTH-1:0]         Ib71065a3fe70d3ab5f05b0c393278631;
wire [fgallag_WDTH-1:0]         I66ba7e48a07f5fdfe16d23b0dc243514;
wire [fgallag_WDTH-1:0]         Ia744719b1036a2236173a80ce326bb7d;
reg  [fgallag_WDTH-1:0]         I984074a5c77445ad266463e20d77899e;
wire [fgallag_WDTH-1:0]         I62e6e8be411f12cd5c4d63f1825521f3;
wire [fgallag_WDTH-1:0]         Ic3f0e0640b27dd1a3bd39f6b9507c7fe;
reg  [fgallag_WDTH-1:0]         I50bb40691aa09c42e0b64a076b50a971;
wire [fgallag_WDTH-1:0]         I2f94d5aad80c081124e3efa3804af183;
wire [fgallag_WDTH-1:0]         I82fa0db281b140ed781dcf5c53625117;
reg  [fgallag_WDTH-1:0]         I753bff437b6c563f5fddf19685405504;
wire [fgallag_WDTH-1:0]         I7a91b23716bf81bea4956eafb467c96a;
wire [fgallag_WDTH-1:0]         I5dfa454e544e731a6254e73c97d79e06;
reg  [fgallag_WDTH-1:0]         I21f2ec69bcc507756e2a5f85d3ead3e8;
wire [fgallag_WDTH-1:0]         I17572136bb435e84505c016523a6ec88;
wire [fgallag_WDTH-1:0]         I3a57ff68cdc9b93c07bc79f8cea77473;
reg  [fgallag_WDTH-1:0]         Iddec4486996054e475499d370016a685;
wire [fgallag_WDTH-1:0]         I9b0ac56afa21022e8bc69f5d20d17b66;
wire [fgallag_WDTH-1:0]         I2f363d2944c634905ef5ec14c9cedf52;
reg  [fgallag_WDTH-1:0]         I3d3edd06f8907f4369b825062348da87;
wire [fgallag_WDTH-1:0]         Id9468cba18d4c67a84cb2b16d2cf495e;
wire [fgallag_WDTH-1:0]         Id15ed601c43171647305818c6f30ace5;
reg  [fgallag_WDTH-1:0]         I72467ef10ecced8395a6870a39525787;
wire [fgallag_WDTH-1:0]         I2bda0265c40a5cedc359dee75fb15b4c;
wire [fgallag_WDTH-1:0]         I75bed085cf80c0672fb41df1d6fc4545;
reg  [fgallag_WDTH-1:0]         I9b74b672f55e7bf7560ba4dd2d0c79fd;
wire [fgallag_WDTH-1:0]         I318ebdf91ab8e83b80a880395879fc77;
wire [fgallag_WDTH-1:0]         Ib7f95eeae4f4565133ae98a0538e56c3;
reg  [fgallag_WDTH-1:0]         I285b012d2fb5e2279a79cf8edca24ac8;
wire [fgallag_WDTH-1:0]         I8ac8dbc25a20c0c27e09240a5cd1bfd2;
wire [fgallag_WDTH-1:0]         I5a7c45c0b4ce4206080f2b50cb0a169f;
reg  [fgallag_WDTH-1:0]         I8faf911a7d1ea8b0abe54f6688068ca0;
wire [fgallag_WDTH-1:0]         Id8c4e5d6318622bd8ec2974684f542b6;
wire [fgallag_WDTH-1:0]         I27cba499cffd339eddcdb4e2c846ee69;
reg  [fgallag_WDTH-1:0]         I3dca974bf2d5631a47ebf8b945efab20;
wire [fgallag_WDTH-1:0]         I8df19e0871c18890419c593410596b59;
wire [fgallag_WDTH-1:0]         Ifafce4fed1394ac5fa8849145960f2b5;
reg  [fgallag_WDTH-1:0]         I12141c45d147b058a9e392f3b7d7d06e;
wire [fgallag_WDTH-1:0]         Ifb977d4c5bac50b9d7f2f814a500f0f2;
wire [fgallag_WDTH-1:0]         I1d6de59e71e329f79055285b3a50c2b4;
reg  [fgallag_WDTH-1:0]         Ia527c96e30b782f837bc6206961400e4;
wire [fgallag_WDTH-1:0]         Id9a1f5bd846dc7d093ed9392722317be;
wire [fgallag_WDTH-1:0]         I9265fbbb34a66f13193ea1220ecb0589;
reg  [fgallag_WDTH-1:0]         I6adbdb64422a08be9bf9e538db97463b;
wire [fgallag_WDTH-1:0]         Ic886ecf946cd5c297012444cb34980ab;
wire [fgallag_WDTH-1:0]         Ifcc01d5d37df8c68972086c44575e8d6;
reg  [fgallag_WDTH-1:0]         I958cdf5367c7b0bd58b70b763d3af8aa;
wire [fgallag_WDTH-1:0]         I37085a233f195dce1a76d05b0157fcac;
wire [fgallag_WDTH-1:0]         I57c25f5b2fecd18092653842e49e8d11;
reg  [fgallag_WDTH-1:0]         I91b7b8e8887b5dd9853297463c55b78d;
wire [fgallag_WDTH-1:0]         Ia2812d1ba8ca6831a2f059eb23384b38;
wire [fgallag_WDTH-1:0]         I4b70004412f2ef37ac00fc19592b1f30;
reg  [fgallag_WDTH-1:0]         I6162978f0c57958ad0403246fb0530dd;
wire [fgallag_WDTH-1:0]         Id176f2681568337762559e78cde29ba6;
wire [fgallag_WDTH-1:0]         Ib952f8ef85514b1832324867adc72ce0;
reg  [fgallag_WDTH-1:0]         I508142e70fd04513977130556aa574ef;
wire [fgallag_WDTH-1:0]         Ia0c4e9942a4b08f69c2a027a712c9e39;
wire [fgallag_WDTH-1:0]         I08494381ebeda641f05b917fa31910a8;
reg  [fgallag_WDTH-1:0]         I2afab673e4b803ffd888f187de47fa49;
wire [fgallag_WDTH-1:0]         I2da299005fed6f2b710e25acd48ebe91;
wire [fgallag_WDTH-1:0]         I3f0568074c465ac281150bb70bbd76ec;
reg  [fgallag_WDTH-1:0]         I7a56f81596920126a9ea2c9fb3a19285;
wire [fgallag_WDTH-1:0]         Ia1038e3b807e16a30f6f4564509ddd30;
wire [fgallag_WDTH-1:0]         Ib6b79505990d6499127f78e3186cc2a8;
reg  [fgallag_WDTH-1:0]         Ic6252de2c819f2243476ddf82e22d137;
wire [fgallag_WDTH-1:0]         I25d94516522c19c0e53b5f52f4480216;
wire [fgallag_WDTH-1:0]         I5404c19d5b4c44dddcca70138fbe79de;
reg  [fgallag_WDTH-1:0]         Ieea8672b2f23711c6ba893de5c5d8bc2;
wire [fgallag_WDTH-1:0]         I4b96be53e3d059113bb74b27ffe30179;
wire [fgallag_WDTH-1:0]         I7265ecc942bf501ad034704f517d4e8d;
reg  [fgallag_WDTH-1:0]         I3a4dbdf517b8f9c93b567f91870e6160;
wire [fgallag_WDTH-1:0]         Ic091d8daff9f609c53cb191ed6b6ddeb;
wire [fgallag_WDTH-1:0]         I1c114e8dfd37b1d182028679b3974a1b;
reg  [fgallag_WDTH-1:0]         I4731ee7a0e08c69e2bd2a8bcea0838c2;
wire [fgallag_WDTH-1:0]         I2468caeaf9733c8bc6a485542b6b263f;
wire [fgallag_WDTH-1:0]         I9fa799fd606c85184ce84138a90f03e1;
reg  [fgallag_WDTH-1:0]         I1b6cbbcf01a65cd1c2f1e241f849c904;
wire [fgallag_WDTH-1:0]         I6611d1fa58dd253fe6344a41584d7e22;
wire [fgallag_WDTH-1:0]         Id8b3ba6e7ffd04674b2ae10b928f26f0;
reg  [fgallag_WDTH-1:0]         I663aee79f824c854f57c19e87207529b;
wire [fgallag_WDTH-1:0]         I8afb33eced17e8675a8e2bd90d16030b;
wire [fgallag_WDTH-1:0]         Id4cc4e9883ae7b27bed350ba292d9349;
reg  [fgallag_WDTH-1:0]         I34ff7299c9d83affa4512b7da302c199;
wire [fgallag_WDTH-1:0]         Idac55755226133905d3250273b1eccb8;
wire [fgallag_WDTH-1:0]         I5c3099cb6fc046e62863a69945ae3e04;
reg  [fgallag_WDTH-1:0]         I70ca6c9d0a5c99e0036479f7b5dd760a;
wire [fgallag_WDTH-1:0]         I4cd564459b8d65976195b2994e7d44f2;
wire [fgallag_WDTH-1:0]         If48b274e1e1809931eb2be69a565a443;
reg  [fgallag_WDTH-1:0]         I835bb7345787eaadc41816858e0a71a1;
wire [fgallag_WDTH-1:0]         I2280162ee1c08ccc9f0c17d1ca0e3628;
wire [fgallag_WDTH-1:0]         I1667cbf3caf9a10527531b6aa69df847;
reg  [fgallag_WDTH-1:0]         I3c7f6fdd0e9cc7426df76027912d1ccb;
wire [fgallag_WDTH-1:0]         I28b3ba64175358f277427fd790a9228b;
wire [fgallag_WDTH-1:0]         I80ddcee29ed7af07148977eddab4bccd;
reg  [fgallag_WDTH-1:0]         I9ff512085174a7720705d0fb37c4ec34;
wire [fgallag_WDTH-1:0]         I6c03138440f9bd0cb2cfe12abf619c10;
wire [fgallag_WDTH-1:0]         I32ab257af6a54e78706c6d83b579bcd6;
reg  [fgallag_WDTH-1:0]         I6a69cdf2bae1ea68c9be56dcc4e76a59;
wire [fgallag_WDTH-1:0]         Ib3709eb9dfc3a594d38ea5a0ef0cd444;
wire [fgallag_WDTH-1:0]         I907f4db1352049380285f358cac2b439;
reg  [fgallag_WDTH-1:0]         I855ddead34ac131137ba644afbfea2b7;
wire [fgallag_WDTH-1:0]         I44cf5ba18d7d029df13f446f09191b2c;
wire [fgallag_WDTH-1:0]         I22cd5fb22f122d99e37e6c1ca2666301;
reg  [fgallag_WDTH-1:0]         Ib1a463388daf270eb0ce698d7b5ded4b;
wire [fgallag_WDTH-1:0]         I6aa1e5acf0c2b01c94438bd1cff484c6;
wire [fgallag_WDTH-1:0]         I892abe227878c5232de3ccd90e8c13e5;
reg  [fgallag_WDTH-1:0]         I74e4bb7530c02073f9b15a6389659d4b;
wire [fgallag_WDTH-1:0]         Ia23629f3881e4119c36576f7da58ceaa;
wire [fgallag_WDTH-1:0]         If5086f7447696a697be414fe50ad91fd;
reg  [fgallag_WDTH-1:0]         I6721b13abeddc76139bdc7380434cc2a;
wire [fgallag_WDTH-1:0]         I2f12d1fa0b815564cefafc28ceb3de82;
wire [fgallag_WDTH-1:0]         I9dc20c15b19d9351497997c81511c744;
reg  [fgallag_WDTH-1:0]         I84fba239c5705bcd92096e204cc9438c;
wire [fgallag_WDTH-1:0]         Ib09ac099bcf61b09922b353403b29987;
wire [fgallag_WDTH-1:0]         I254c64de80d2a159aa0b3f3170042079;
reg  [fgallag_WDTH-1:0]         I4d46e4d50176768fda897949545e2125;
wire [fgallag_WDTH-1:0]         I3c2b6da8e286d0a7b628ba1071f29424;
wire [fgallag_WDTH-1:0]         I4dae38e87f09d78c748974da00f274f8;
reg  [fgallag_WDTH-1:0]         I57086cfab3b163c3911c3cf7bfb3141a;
wire [fgallag_WDTH-1:0]         I550630b507ceec38b960ab2a86a57f1a;
wire [fgallag_WDTH-1:0]         Ic8edf24599f1eee2af3576dfb2a6829a;
reg  [fgallag_WDTH-1:0]         Ice174debd5dc911fdf5d5756cff8d731;
wire [fgallag_WDTH-1:0]         I795c1c91cb6b7870b7efb07d67085be1;
wire [fgallag_WDTH-1:0]         I144ca4c629cc3134a991414038cfc9cf;
reg  [fgallag_WDTH-1:0]         Ie369670edc5b602d305904f3a4a4381f;
wire [fgallag_WDTH-1:0]         I531b70d12349f3bc67e6a3ec53368d97;
wire [fgallag_WDTH-1:0]         I379ed527c944420bb59be58b85ab4704;
reg  [fgallag_WDTH-1:0]         I41f66f79339962ef42fab3b88e571170;
wire [fgallag_WDTH-1:0]         Id8a109043bc922b718c203bd5d60a999;
wire [fgallag_WDTH-1:0]         Id37ddd7be0621f84793d1600ce915236;
reg  [fgallag_WDTH-1:0]         I5cbd2fad4d90bd77ba3d2448a37ac60f;
wire [fgallag_WDTH-1:0]         Ic126109499ee1dc2787ab05b404e7ae2;
wire [fgallag_WDTH-1:0]         I20bbdbbee46a2be5c6caa56786345e8b;
reg  [fgallag_WDTH-1:0]         Id86a2869148e2885633d9e277f7041c3;
wire [fgallag_WDTH-1:0]         I1cd8ba53b876e2436901749e355f354b;
wire [fgallag_WDTH-1:0]         I02199c9dc39a2c8be49a1c96aa89de15;
reg  [fgallag_WDTH-1:0]         Ifb7b585189db23efabfb522c9b45bede;
wire [fgallag_WDTH-1:0]         I4e8ff51a6f70f8ca6a17a1dea8caf0a9;
wire [fgallag_WDTH-1:0]         I17b1742efeadf5df716128d6603ebe99;
reg  [fgallag_WDTH-1:0]         I7763f0d28d8065d8c94ef8df96b2ab06;
wire [fgallag_WDTH-1:0]         Ic1a27480c9acc1684f3fed116d74cb5f;
wire [fgallag_WDTH-1:0]         I68da2c2a43373cf8145e6f7072bb5ca9;
reg  [fgallag_WDTH-1:0]         I115ba88588187c7115977e95bd26ee5a;
wire [fgallag_WDTH-1:0]         I0df7a888610865486aa1aaa2703dd041;
wire [fgallag_WDTH-1:0]         I27f3ef61a2ffbd4154a7b683aacd4844;
reg  [fgallag_WDTH-1:0]         I6e7f2bdd0c8231a3689893ef4877fdba;
wire [fgallag_WDTH-1:0]         If6448c72403a3d0bd904beac87f8aa96;
wire [fgallag_WDTH-1:0]         I0726f4d2f2b1d495b1b439f998193435;
reg  [fgallag_WDTH-1:0]         I546c513d5357ac1a6fe669888dfaf717;
wire [fgallag_WDTH-1:0]         Iecf45496b391208d62e88544b5d2ca49;
wire [fgallag_WDTH-1:0]         I05e3c3e8567ed11012cf9f9d7ecb629a;
reg  [fgallag_WDTH-1:0]         Ib3e12c614471912d0b276cb9f0382b1b;
wire [fgallag_WDTH-1:0]         Ib0fd0a839c85f3da5ae7b221f6e623d6;
wire [fgallag_WDTH-1:0]         I210ade98fc479cdb069e2b028f1920d4;
reg  [fgallag_WDTH-1:0]         I7187a2499e3319da90b6d6fc64411b46;
wire [fgallag_WDTH-1:0]         Ie045750c9289c899860823f90a306f3c;
wire [fgallag_WDTH-1:0]         Ic89a704c9de69cff5b09d1b3bb220fe8;
reg  [fgallag_WDTH-1:0]         I9b46582473bb4dd5541a35ac708486f4;
wire [fgallag_WDTH-1:0]         I1627b19e0ca42f9c264b626809fb37b7;
wire [fgallag_WDTH-1:0]         Ic8ba8abf8a87610d08fb5a8174639f99;
reg  [fgallag_WDTH-1:0]         I929796fe327ee9c8a05e6bb683ae5d7c;
wire [fgallag_WDTH-1:0]         Ic9593f3fe23f258c2ab4ddcadaa8ca4c;
wire [fgallag_WDTH-1:0]         I9c0a1bb49be6604f75611b92d937c124;
reg  [fgallag_WDTH-1:0]         Ib6638da8b69373c2026d3f5305825cde;
wire [fgallag_WDTH-1:0]         Idc0085a6595a7de7e2bc87c789b7d935;
wire [fgallag_WDTH-1:0]         Iff70fe838ee16e8e35b1034135555acc;
reg  [fgallag_WDTH-1:0]         I28c26bf4cf9693d1807818b2ca7883ac;
wire [fgallag_WDTH-1:0]         Id029b4c310acea870263d3715689e729;
wire [fgallag_WDTH-1:0]         Ibb4daaccffcf82b4cb4c431923c71f3f;
reg  [fgallag_WDTH-1:0]         I291fc4eef4b80d1020c96488b869727e;
wire [fgallag_WDTH-1:0]         Iec123ddb8d1e623d03d85a667c97ef31;
wire [fgallag_WDTH-1:0]         I9c1fd2b57c1756bf67bc8cf5ed4a1912;
reg  [fgallag_WDTH-1:0]         I53006ed50f6211439681aa7659647e35;
wire [fgallag_WDTH-1:0]         I89f0b0713e165a454e187fa51e89c642;
wire [fgallag_WDTH-1:0]         I71d437815bcfb755e16fc442431b6f68;
reg  [fgallag_WDTH-1:0]         I47fe32973727237ae0cd4c306c7efbfb;
wire [fgallag_WDTH-1:0]         Id812cf3919ed50a5e3897d129eeb4b8d;
wire [fgallag_WDTH-1:0]         I4e3e1eb8ea6dfb08ea2634a9bab8319b;
reg  [fgallag_WDTH-1:0]         Ic3e0c7d71f13a56a9a63e158c7f2cfa8;
wire [fgallag_WDTH-1:0]         I2d65b5115be2a22ed1e29426be3f0d15;
wire [fgallag_WDTH-1:0]         I1fa2749e15c3bd7253a023eb01140cc7;
reg  [fgallag_WDTH-1:0]         If383f241447cbea4e18f4f79fcdbf144;
wire [fgallag_WDTH-1:0]         I47c8671569e2c5c2a21f27aff2d1f4b8;
wire [fgallag_WDTH-1:0]         Ie19e8502010d0c178f9f2da8df3fa63d;
reg  [fgallag_WDTH-1:0]         Ia05354d3b4f61299d5897832639df2c2;
wire [fgallag_WDTH-1:0]         Iaf2144dab2167cd2629067e40bea3053;
wire [fgallag_WDTH-1:0]         Ia512ada6f00f86ff495ae12ead6607d3;
reg  [fgallag_WDTH-1:0]         I9faec40665477e8b3237773d606af2f0;
wire [fgallag_WDTH-1:0]         I4c2b80e4bbbd4c5e8d0da28c5d0f681e;
wire [fgallag_WDTH-1:0]         If7b2398d3426250d73917539ff743c8a;
reg  [fgallag_WDTH-1:0]         Id231ab3133d4bed02aad7e5f560ee5f0;
wire [fgallag_WDTH-1:0]         I6300fbbd385ad9280c751076bc68d70c;
wire [fgallag_WDTH-1:0]         I6446a839157f78880fc3fc7d8c378c78;
reg  [fgallag_WDTH-1:0]         I13616c8c7be221cf4d2c13ae87c38bed;
wire [fgallag_WDTH-1:0]         Iea078843b3c5139a395997c54462850a;
wire [fgallag_WDTH-1:0]         I53504e8899a821cebe69ed590a3fd7fc;
reg  [fgallag_WDTH-1:0]         I8793bc728a4d423fb96a88c83bb9746f;
wire [fgallag_WDTH-1:0]         I654debf65019f2748e631a051f3b17ca;
wire [fgallag_WDTH-1:0]         If7d5fe39b147f24303884de3a30d669d;
reg  [fgallag_WDTH-1:0]         I2fb6af0f152232550a3cadd55656df20;
wire [fgallag_WDTH-1:0]         I1e88b57c19a1ddfc1c1f0e168b60f814;
wire [fgallag_WDTH-1:0]         I24c005d076b3c887d45d1285a4fe1bc5;
reg  [fgallag_WDTH-1:0]         I5144918fcd4ce1a061644240730fc52a;
wire [fgallag_WDTH-1:0]         Ibaf7ab7333434b0d7e76e436ee40a406;
wire [fgallag_WDTH-1:0]         I18e00688f19c522b305d223ead684fb7;
reg  [fgallag_WDTH-1:0]         I1821eb21cdf8208ff6c2f28d963f7bd6;
wire [fgallag_WDTH-1:0]         I1af14572832bd6d6b5890b8340b79ec7;
wire [fgallag_WDTH-1:0]         I0258ec63762460afb41bcd6e8869ec69;
reg  [fgallag_WDTH-1:0]         I80471575b1d4b69ef073056f798394ea;
wire [fgallag_WDTH-1:0]         I652d3ed935b39f8fda8d84296456d633;
wire [fgallag_WDTH-1:0]         Id1280129b20bd6389618695aec9efeed;
reg  [fgallag_WDTH-1:0]         I890bf9b72cc3c71351547178d72796e5;
wire [fgallag_WDTH-1:0]         I5e33cad360aae934f418852541f5f2bd;
wire [fgallag_WDTH-1:0]         I907fd3abdcadda1cd7149c7cf01e5751;
reg  [fgallag_WDTH-1:0]         Icc9d28b84fa91028ae96cc9b8bae7555;
wire [fgallag_WDTH-1:0]         If950e448e3cba7cc9aa7aff7718775f7;
wire [fgallag_WDTH-1:0]         I73f044469c4dbcd5a98c0f83d6d043c4;
reg  [fgallag_WDTH-1:0]         I0b0d167c415f8c14594bd61907d46d80;
wire [fgallag_WDTH-1:0]         I9adf8836419a1c85b146e5e36de68af5;
wire [fgallag_WDTH-1:0]         I2934a8783b90254606bcd933c629577f;
reg  [fgallag_WDTH-1:0]         I9577d49a74520355e53a1818f479db0e;
wire [fgallag_WDTH-1:0]         I0f2bcdf124dff4219fd1a35ed1db7937;
wire [fgallag_WDTH-1:0]         Id26b2a9c13424769e1627b1549159a7e;
reg  [fgallag_WDTH-1:0]         Ie6e888d582ba9e600e91b119e2804642;
wire [fgallag_WDTH-1:0]         Iae82e5de28b12f962bd7c5e221317ac2;
wire [fgallag_WDTH-1:0]         I2115e45deea528402794afadd17d9fe7;
reg  [fgallag_WDTH-1:0]         Iccfac3d489b4b110d6b6e005a5ba45d8;
wire [fgallag_WDTH-1:0]         Ia7b3cb9de8e18f41561c2a46dda8696a;
wire [fgallag_WDTH-1:0]         I978020f8aaeb98cc1cea9360ec06da22;
reg  [fgallag_WDTH-1:0]         I69a67481ca8fd01dc5400dbe887b4f83;
wire [fgallag_WDTH-1:0]         Id0119672c8b017bce6fdba53d4dccf8b;
wire [fgallag_WDTH-1:0]         Icded30641e4770e30ee34bbf8d2a5721;
reg  [fgallag_WDTH-1:0]         I1f36f045becec7f0528f4a935d3da2ff;
wire [fgallag_WDTH-1:0]         I4aaef2f654ba03b1dc05719c81d5da69;
wire [fgallag_WDTH-1:0]         I02e3cbacce4e97e3088360f0acccee44;
reg  [fgallag_WDTH-1:0]         I530fe7720e3bcda35e940aa4973a7da4;
wire [fgallag_WDTH-1:0]         Ia6355e548635a4107a11c7952aa8b3d9;
wire [fgallag_WDTH-1:0]         Icbdf81888af42710561aec48ce84e3cb;
reg  [fgallag_WDTH-1:0]         I03069dda9fa863172d8747408800eeba;
wire [fgallag_WDTH-1:0]         I0bd950eee6abde9d1eaaabbe902fff5d;
wire [fgallag_WDTH-1:0]         Iea3ce04a4b8cc466e892aab886e63744;
reg  [fgallag_WDTH-1:0]         Ie7f36ee89f2b092555fbf8031d2347d9;
wire [fgallag_WDTH-1:0]         I93caf487f67a2adce04a7b2cd7fff358;
wire [fgallag_WDTH-1:0]         I3ca9464d884ccc7e2f396a74baea5bb9;
reg  [fgallag_WDTH-1:0]         I18af7980562b28c537be3bea8dc5252b;
wire [fgallag_WDTH-1:0]         If68a9cc5609ea7d87062bad2ebddb1a8;
wire [fgallag_WDTH-1:0]         I7b8d02aa08cde64a409f3766f940233c;
reg  [fgallag_WDTH-1:0]         I22ec20f9396d28ed39c5fc4bf060c44a;
wire [fgallag_WDTH-1:0]         If201a7afedfd1c329b55048e6bbad629;
wire [fgallag_WDTH-1:0]         I86ad427fe92cd4346b32ecf3c99c93c7;
reg  [fgallag_WDTH-1:0]         I105eac4e38f4661c7c7ca32161e42baa;
wire [fgallag_WDTH-1:0]         I1f8936599ead5ce1cd85132e382533f1;
wire [fgallag_WDTH-1:0]         I6667614b2fe12d6f63ac7737bf069b42;
reg  [fgallag_WDTH-1:0]         I5030734bfa54065cbef20c1350cd647d;
wire [fgallag_WDTH-1:0]         I37eb148270af62adba8341c83411f9f2;
wire [fgallag_WDTH-1:0]         I909cbd582f015b4eabefd660b2039ccc;
reg  [fgallag_WDTH-1:0]         Ieccf25e3abd6bae7dcf08baf815f3439;
wire [fgallag_WDTH-1:0]         Ie4729048b95fede1806dbd006de01338;
wire [fgallag_WDTH-1:0]         Ie3433004b0ea3bba81f0b7502c69c821;
reg  [fgallag_WDTH-1:0]         I600c21fca7901299f8e95e8fa0ea0eb0;
wire [fgallag_WDTH-1:0]         I02330d212434a6e8c303db2c3d36a3e5;
wire [fgallag_WDTH-1:0]         If548fc27869a7e48fedc89bd5c8037f0;
reg  [fgallag_WDTH-1:0]         Ic4363dfd133124dd45ec2211499d0788;
wire [fgallag_WDTH-1:0]         Id89498cf205e0cdef4886afd878c48f6;
wire [fgallag_WDTH-1:0]         I7cc21b5c21f6bc0603c3d57c86feeb00;
reg  [fgallag_WDTH-1:0]         I7c0bc779c09847e3beb0a139e8826511;
wire [fgallag_WDTH-1:0]         I547ae5055196f12eeeb36d69c325b84d;
wire [fgallag_WDTH-1:0]         I9ce2b40cd4433999690bb6e5c368e9b8;
reg  [fgallag_WDTH-1:0]         If64db4386bf8f7d07292f14e3b313520;
wire [fgallag_WDTH-1:0]         I4871ccbe2f182791243b7bdcc9b8e286;
wire [fgallag_WDTH-1:0]         Ie102c1592ae8606ab75b1f7101b44918;
reg  [fgallag_WDTH-1:0]         Ibf51e537b992c4b4c0539dda9948f45c;
wire [fgallag_WDTH-1:0]         I12fd829f22ba908180290432320a3660;
wire [fgallag_WDTH-1:0]         I23ef94c5c29e674714d4ea1ad2d3f0e8;
reg  [fgallag_WDTH-1:0]         I9f83063bdc3c352024f702cb9dc71ce8;
wire [fgallag_WDTH-1:0]         I8f967710d03870e026564db0df46d146;
wire [fgallag_WDTH-1:0]         I990c1f1dbce95ae4dfc62588c9cc9e1f;
reg  [fgallag_WDTH-1:0]         I72127f6d422ec68dcd47126b87b3d3b1;
wire [fgallag_WDTH-1:0]         Ia347d80a70a49605c51d19bc2e696aef;
wire [fgallag_WDTH-1:0]         I9d2e71f9a6d7eb4221978fef3c10d678;
reg  [fgallag_WDTH-1:0]         I0b4a1b48d110b820d8d87f6e94d32988;
wire [fgallag_WDTH-1:0]         I730db85d3d11d8327c6d48b8b87a00a4;
wire [fgallag_WDTH-1:0]         I34754a80000aa92f8a7e4997b91f6d07;
reg  [fgallag_WDTH-1:0]         I2e3aeede695007fabe0d6247a93ed403;
wire [fgallag_WDTH-1:0]         I5c6a3ec08cb17d6646bb3e63411a9698;
wire [fgallag_WDTH-1:0]         I055273589d8d967bd5e255808051a101;
reg  [fgallag_WDTH-1:0]         I8c5ea3dc59fdcdea1c5f503dde1e815f;
wire [fgallag_WDTH-1:0]         I7b5baeec7b11eca457dcd9d2b2b64ac5;
wire [fgallag_WDTH-1:0]         I5142a2511a55a7ad420618d874b0dddd;
reg  [fgallag_WDTH-1:0]         I873c4dbe95220e40d7388870520261bd;
wire [fgallag_WDTH-1:0]         Ic4c7a9d491c560d7b6c410d8216f59bf;
wire [fgallag_WDTH-1:0]         I5e008272bf3a470d74ca6b5cf39bf28f;
reg  [fgallag_WDTH-1:0]         I561fa67a9bfbedffcb04e7a4d6b76a64;
wire [fgallag_WDTH-1:0]         I2151735079b41a7f8cbfe2b93f1b7470;
wire [fgallag_WDTH-1:0]         I5c31bbaf08a6e8971f585cdae36384f5;
reg  [fgallag_WDTH-1:0]         Ia55752d6c4f20378ff570a661ab31d9a;
wire [fgallag_WDTH-1:0]         Ia69e34af60619fa04e8478e2d04768bb;
wire [fgallag_WDTH-1:0]         I509af9c5f9d6bf3be233847dbd05e3fa;
reg  [fgallag_WDTH-1:0]         Ia13307be43e9155ed0333df62ccc8bf2;
wire [fgallag_WDTH-1:0]         I7f9984597d0e7bcda92f13fbb8805687;
wire [fgallag_WDTH-1:0]         I3182472e08e707cbc36d60ba54613129;
reg  [fgallag_WDTH-1:0]         I07b3d1451487a55fbbedda48b0cb6c73;
wire [fgallag_WDTH-1:0]         I342ef25fefdb6a326dac80d76052bbd9;
wire [fgallag_WDTH-1:0]         If2455c2d04521a8d8c59965759eb328b;
reg  [fgallag_WDTH-1:0]         I9f8cf1a6cd0182fba35a49bd232f062a;
wire [fgallag_WDTH-1:0]         Id1414254ab35ee805c4010432eb24243;
wire [fgallag_WDTH-1:0]         Ib759c72355cd6e146edb26ad106a0418;
reg  [fgallag_WDTH-1:0]         Ie2e488a8589559deeec8598cf6726f1f;
wire [fgallag_WDTH-1:0]         I8db7cc6cb4bf55131bee6b00e76baf46;
wire [fgallag_WDTH-1:0]         I6826c8a05953c4df79e31a19adfa2693;
reg  [fgallag_WDTH-1:0]         I9118ee5ff8c9ba9b125e5baa07bf52e0;
wire [fgallag_WDTH-1:0]         I355aec2468fa96e2f32c8c324c48c5f5;
wire [fgallag_WDTH-1:0]         I56122ba51d99f9ca67828649860d409e;
reg  [fgallag_WDTH-1:0]         I13b894057e2deae2c00787385de252a8;
wire [fgallag_WDTH-1:0]         Ic45ea6e09fd20a2285b7e6e2507910f4;
wire [fgallag_WDTH-1:0]         I1bcda37ae1a26452a3443142fbee54f9;
reg  [fgallag_WDTH-1:0]         I7797a3ea5b97b514a797243cf9fe890a;
wire [fgallag_WDTH-1:0]         I288b192ad6d04370df8084511c7f44ce;
wire [fgallag_WDTH-1:0]         I3f7dda67dc14fdf45bfb9c4e01dd7f38;
reg  [fgallag_WDTH-1:0]         I3af78697aacc410108d0be7fd13c686b;
wire [fgallag_WDTH-1:0]         I4d589e9479ee494636d90a910e530863;
wire [fgallag_WDTH-1:0]         I6fd4da8e1e3cb360964d6e425d174465;
reg  [fgallag_WDTH-1:0]         I871cb63247618a543b444aa3f888fffe;
wire [fgallag_WDTH-1:0]         Ib8fcb6e6569d34c67145861431ad5334;
wire [fgallag_WDTH-1:0]         I5f7baab0fcf12df1e886e17375732c04;
reg  [fgallag_WDTH-1:0]         I124404013f8fc6b302661900b9ad8ed8;
wire [fgallag_WDTH-1:0]         I5405b3c646988338f12191bb8cb02205;
wire [fgallag_WDTH-1:0]         I87303a5c7e205b0b1b196ae97a0c994f;
reg  [fgallag_WDTH-1:0]         I8e413271c9d13748a1aa2d1a018ff28f;
wire [fgallag_WDTH-1:0]         I371946ff4a809b62ceed2334a9656787;
wire [fgallag_WDTH-1:0]         I5ebd9eab33e2e8cd6b2f7c1f3bd2e39f;
reg  [fgallag_WDTH-1:0]         I4d799e93b4dfcabd69977ddb25634a69;
wire [fgallag_WDTH-1:0]         I6d5be8ddd471c1ddf781949169bd9807;
wire [fgallag_WDTH-1:0]         I7f4bd63152869ed52c49aa41eea5ea1e;
reg  [fgallag_WDTH-1:0]         I1487f0027b7d16f4bc85bb00e537cbaf;
wire [fgallag_WDTH-1:0]         I499f6bbf3456d23378ff02b6f65a5ae4;
wire [fgallag_WDTH-1:0]         Id243e47daf8a5e75fe52a828af95b5aa;
reg  [fgallag_WDTH-1:0]         I1a5cdaa10022adf0ffbbc0f58b3e690a;
wire [fgallag_WDTH-1:0]         I0c81821914371a777679053e2aa5a55e;
wire [fgallag_WDTH-1:0]         I62bd2c30206c591bcb87f31543bda72e;
reg  [fgallag_WDTH-1:0]         I98246759d003e9bc6676ceb2d093a06b;
wire [fgallag_WDTH-1:0]         Ief591e9d4759a4b1059574bb624e4ce6;
wire [fgallag_WDTH-1:0]         Ic1238f5f1f2011fa1869cdb2f50e6a30;
reg  [fgallag_WDTH-1:0]         Ia3c2dfb3c4a45091be7cfecfad11f3ec;
wire [fgallag_WDTH-1:0]         Ie40648c85ed87c979a54dfc1f85d1cc8;
wire [fgallag_WDTH-1:0]         I7f2885836616ac775eb9406e8f5d5214;
reg  [fgallag_WDTH-1:0]         I74cda651bcb24472a7697ba017f831a4;
wire [fgallag_WDTH-1:0]         I36956634f94d6053aa455b29bc0b7a0f;
wire [fgallag_WDTH-1:0]         If1608747d211db3fdf51ecf7464c494c;
reg  [fgallag_WDTH-1:0]         Id7ba55b14ac0f471142011dc2d57cc4b;
wire [fgallag_WDTH-1:0]         I05a652e83a9b8c2c38de64de6a70f8bc;
wire [fgallag_WDTH-1:0]         Iccd84e19d39b19bec98dad532ea5b3ce;
reg  [fgallag_WDTH-1:0]         I5890643c88c4255a0e5efd45f8af3ee2;
wire [fgallag_WDTH-1:0]         Iaefa87388884b85eed690e9917bc9d5b;
wire [fgallag_WDTH-1:0]         Idf7e508a586310bf4ca23c84f8240691;
reg  [fgallag_WDTH-1:0]         I4f53e4955e9e506a7169ae810da5dde6;
wire [fgallag_WDTH-1:0]         I98836c38732b8da439946aa5fcbbd963;
wire [fgallag_WDTH-1:0]         Ic8ef3162d3d0c57faf5dd1bddef1622a;
reg  [fgallag_WDTH-1:0]         Ifc7c1ea337b122fb720767f1890f1a6a;
wire [fgallag_WDTH-1:0]         I8ff116e234a1007cc47989f3fdcf88d6;
wire [fgallag_WDTH-1:0]         I68115420b3b9b8ca8ca584c260e924ec;
reg  [fgallag_WDTH-1:0]         Id40d6f3a8dd09678b25b3e579dd5fb68;
wire [fgallag_WDTH-1:0]         I53dfee31709f8eca30897d6bf1618418;
wire [fgallag_WDTH-1:0]         I5bac906cb51bae905ea33717fe015201;
reg  [fgallag_WDTH-1:0]         I7002830b0a5f40ba2a2fe7a00c7b6d58;
wire [fgallag_WDTH-1:0]         I3ac389b6b81baf93095cc3e9e9c3d8ef;
wire [fgallag_WDTH-1:0]         I9f261cb4883275f5f9187a1a6e8fee08;
reg  [fgallag_WDTH-1:0]         I3f377e8994959ef8182a08538e393d9a;
wire [fgallag_WDTH-1:0]         Ief52e91e9170809b980aa881bf76957a;
wire [fgallag_WDTH-1:0]         Iecfe32305d22e6d91c3f7d4af2ad9d2f;
reg  [fgallag_WDTH-1:0]         I71bf29f3519e3238cec112ef97ce0579;
wire [fgallag_WDTH-1:0]         Iebf813928bcad8ee3b6911057c59752b;
wire [fgallag_WDTH-1:0]         Ib30aa869fd577fb3315608a85947dc7d;
reg  [fgallag_WDTH-1:0]         Iaa4bc2f51984f383479b597e6cd4c873;
wire [fgallag_WDTH-1:0]         I57ae0d331753595cd56d45a28cd5c790;
wire [fgallag_WDTH-1:0]         I82209dd60aeaffa4b05b38230c27147b;
reg  [fgallag_WDTH-1:0]         I9066a5cf776f80ebf89bdac1f2edb4ac;
wire [fgallag_WDTH-1:0]         Ibd173152b9400b4c8011451d68b07e4c;
wire [fgallag_WDTH-1:0]         Ifa110a9cdb359c2b0567d25d4dba725a;
reg  [fgallag_WDTH-1:0]         I7319203d7231bebb6d6e52422cce5ed2;
wire [fgallag_WDTH-1:0]         Idc21b018b7b6f2e0bc627e8968e06eda;
wire [fgallag_WDTH-1:0]         I1451eec261d2367ec6e7b2d50a20679a;
reg  [fgallag_WDTH-1:0]         I4e8309976fd6011d78728cef935dc3c1;
wire [fgallag_WDTH-1:0]         I783423950d0e0229826b2249f5cfdf5c;
wire [fgallag_WDTH-1:0]         Id8f178b6565e3a57c5370aaad14f0639;
reg  [fgallag_WDTH-1:0]         I5ed502118c175d5bdb4607973554a3a3;
wire [fgallag_WDTH-1:0]         I6b8fc6d29fb4549e3f191f913bccff9e;
wire [fgallag_WDTH-1:0]         I67fb672706bbd331c27ab1eb386c24b5;
reg  [fgallag_WDTH-1:0]         If457f80b3d29b60b840f886fa928297c;
wire [fgallag_WDTH-1:0]         Idc98380b110c22495027a7cdb6f2029d;
wire [fgallag_WDTH-1:0]         I112661c3273bde5c91b800dd8ddb08a9;
reg  [fgallag_WDTH-1:0]         I7e0f785ec7554540c9a4a413a3afa75f;
wire [fgallag_WDTH-1:0]         Ieb72df81e325eda4d80a237454fa9dbd;
wire [fgallag_WDTH-1:0]         Ia4979ed96ea3e7332635e1f1a14d9ed4;
reg  [fgallag_WDTH-1:0]         Id3662bbe1b5191995d1656045fe6b6a6;
wire [fgallag_WDTH-1:0]         If70e7ed8d4989cd75d37af1dc5d185ed;
wire [fgallag_WDTH-1:0]         I11a094c5fa993419d19f6361157d6ad0;
reg  [fgallag_WDTH-1:0]         Idf922fab93bc2357ac1f66f73f3ead0b;
wire [fgallag_WDTH-1:0]         Ifc99661bc592c2c43bae53db10c8d472;
wire [fgallag_WDTH-1:0]         I38007605c51aa852477e1901bdd292f0;
reg  [fgallag_WDTH-1:0]         I780371393ef898aa144c5bc36e74c654;
wire [fgallag_WDTH-1:0]         Ic8860cc8d323e5a4c68233109ed70512;
wire [fgallag_WDTH-1:0]         Icae30bad38ea69b85fa826ad52e25a51;
reg  [fgallag_WDTH-1:0]         I79696cd10cffa4c0181a2089da6b3262;
wire [fgallag_WDTH-1:0]         I439288f09536ca87fa0feb5f6436716e;
wire [fgallag_WDTH-1:0]         I1afd8ef52cb1eef06769b7a27c95fa03;
reg  [fgallag_WDTH-1:0]         I073155ab0359a13b77f730653dcfc08d;
wire [fgallag_WDTH-1:0]         I66c4beb8fe2d9f363c8e153a12f216ca;
wire [fgallag_WDTH-1:0]         I9c5442889b71c19de290cf33fa393bd9;
reg  [fgallag_WDTH-1:0]         I1b44f781d81438654f69bb7fbdb94011;
wire [fgallag_WDTH-1:0]         Ib2a96d55b1f7bf9b89286de32e59fad3;
wire [fgallag_WDTH-1:0]         I772891870fc29b32eeed162f198217e9;
reg  [fgallag_WDTH-1:0]         Id68f1a0ec8ff80da3190fe517bd935e3;
wire [fgallag_WDTH-1:0]         I3028dabd706c9e5768eac56c66463955;
wire [fgallag_WDTH-1:0]         If4167812b028552487002b44bdae0caa;
reg  [fgallag_WDTH-1:0]         I3704464d41956032b779eebe27511815;
wire [fgallag_WDTH-1:0]         I265f3da3571d2ddb786b98ba3959823b;
wire [fgallag_WDTH-1:0]         I4d470ec03c4967c49989f59671d735bc;
reg  [fgallag_WDTH-1:0]         Ie6756ee9631791940ffc6fddb223b4d0;
wire [fgallag_WDTH-1:0]         If8d81c152d863660081339144b37a052;
wire [fgallag_WDTH-1:0]         Ia28efddccf0f15c926e3901002bf6c9f;
reg  [fgallag_WDTH-1:0]         I085151dfc2e773a7a485f5ef1b7cd6bd;
wire [fgallag_WDTH-1:0]         Ie9cba6422546d378655d0ef98ef974fb;
wire [fgallag_WDTH-1:0]         I1f3c6900aaf35b7e0cf71c04d917cb71;
reg  [fgallag_WDTH-1:0]         I2654e83fff153df7760c341f59a23396;
wire [fgallag_WDTH-1:0]         Iaddf6de71a6329eb536f54e3d18d43d6;
wire [fgallag_WDTH-1:0]         I8788a098d0d9b94af7b93f6b5ef0cce2;
reg  [fgallag_WDTH-1:0]         Iee3eec7a9d7a3a5c22281545ec143e50;
wire [fgallag_WDTH-1:0]         I280ed7bf157554fcad915f0e7fa12653;
wire [fgallag_WDTH-1:0]         I46a61c4cc712f8ffcf45f93d11f0e146;
reg  [fgallag_WDTH-1:0]         Ied2b9ca07a6d498abada30fb0726df24;
wire [fgallag_WDTH-1:0]         I0ca797b233dcdac8e390e1e41d99b196;
wire [fgallag_WDTH-1:0]         I2a826f08bf1fc30c125cdb9a93bea1b3;
reg  [fgallag_WDTH-1:0]         If95315702519e7a08386a870e599aab0;
wire [fgallag_WDTH-1:0]         I150792edd72cc07cf8242d787cb52056;
wire [fgallag_WDTH-1:0]         I2614ad9be5eee336ad67441c050bd366;
reg  [fgallag_WDTH-1:0]         I1091064aef7d915ba8fb6cbded069102;
wire [fgallag_WDTH-1:0]         I186c13747ff5a1ee6e562ad9e5faabd9;
wire [fgallag_WDTH-1:0]         Iecd35290f27c4375873e964f2db90ba9;
reg  [fgallag_WDTH-1:0]         I40685c7d2c8be12698f734ec6213b5b4;
wire [fgallag_WDTH-1:0]         I6fb8240f8c68b71cafe4c2c43ac7db33;
wire [fgallag_WDTH-1:0]         I9b90edd08194934b456cf88beedf8785;
reg  [fgallag_WDTH-1:0]         Icc7775fe34c162006b93662530fd4944;
wire [fgallag_WDTH-1:0]         I166f5cab59c2a66117f2287d2b11c096;
wire [fgallag_WDTH-1:0]         I7db63c5bb5e53cbc83051b5c80c1a19c;
reg  [fgallag_WDTH-1:0]         I2e6f1a5695ad23b8ca282b344832ee8e;
wire [fgallag_WDTH-1:0]         Ie896986a747c1cd8ccad7117125c6e0d;
wire [fgallag_WDTH-1:0]         Iaec5353d68ad9092c0fb74683f876213;
reg  [fgallag_WDTH-1:0]         I016ce894bebdaa7e56af9deb1ccfb3f5;
wire [fgallag_WDTH-1:0]         I0c829f14ef188ff7ae1417e28903f2b3;
wire [fgallag_WDTH-1:0]         Iec7f88e1ed763c1f55c90b39870875c2;
reg  [fgallag_WDTH-1:0]         Iad2dd0815c1107160992e5070632f76c;
wire [fgallag_WDTH-1:0]         I3591d4f320f8401ef8ad8f92d2d89bf6;
wire [fgallag_WDTH-1:0]         I32f96b4803590ac0f86d2178cac9e4a8;
reg  [fgallag_WDTH-1:0]         Iefaba2acd282081b9a0a98ed057ca85e;
wire [fgallag_WDTH-1:0]         I3816895f23a1381e42aaeb64dd158fda;
wire [fgallag_WDTH-1:0]         Idc0fc3de3b05c5beebbf24649662f02e;
reg  [fgallag_WDTH-1:0]         Id4ef94eb8d5db8810bca4c9d669f0b7f;
wire [fgallag_WDTH-1:0]         Ic9c34a36b2fde9649064680904ec9150;
wire [fgallag_WDTH-1:0]         I9d54e626fd0b2e435b117ae6b5d5e194;
reg  [fgallag_WDTH-1:0]         I04e845e6a5ed71978b636593dd749b12;
wire [fgallag_WDTH-1:0]         If7eb75eccc5a6384c80d99b64d534fca;
wire [fgallag_WDTH-1:0]         Id5cff86905cde551a008a19305e87f94;
reg  [fgallag_WDTH-1:0]         I0b2760b437be2cb79382f8d6a7b8969e;
wire [fgallag_WDTH-1:0]         Ib788a897a1d1b86b2c16caade11846ee;
wire [fgallag_WDTH-1:0]         I3837a2e882da18f37f074b51cf5cbf85;
reg  [fgallag_WDTH-1:0]         I1b0fdaeebe5fee6fbb2e13aac5e233a1;
wire [fgallag_WDTH-1:0]         I6a5fec9dad124f6d8c5574bcc2643ede;
wire [fgallag_WDTH-1:0]         Ib584dc3e5dd346562062794c0f1c5f9e;
reg  [fgallag_WDTH-1:0]         Iee872d17e4a28075be0ad7086c3acc91;
wire [fgallag_WDTH-1:0]         I3936f324b08bea1bc5f8bcd12437b161;
wire [fgallag_WDTH-1:0]         I20ac1027f7da12ad62120cd3b0603c7e;
reg  [fgallag_WDTH-1:0]         I87656ddd4ef8f1ae36c7566d5e7892d8;
wire [fgallag_WDTH-1:0]         I1a59337d4da3e3ad1a738a9c3b56ef8c;
wire [fgallag_WDTH-1:0]         I8adacef11a4f33ff1ccea285fd1a8b74;
reg  [fgallag_WDTH-1:0]         I865cd0535644db7f17db1180c85f1744;
wire [fgallag_WDTH-1:0]         Ic3e3b4cba05d80c0ceaa6e25a906a602;
wire [fgallag_WDTH-1:0]         Ie2ad82bbff584541911e13b90a5d15a0;
reg  [fgallag_WDTH-1:0]         I71d46741fa94df65e1bdf6abff53d2ba;
wire [fgallag_WDTH-1:0]         Ife0830e12b8bbb5aa0b8c2c0e4191e59;
wire [fgallag_WDTH-1:0]         If6243c5fc2ec9a15eecf227b234434d1;
reg  [fgallag_WDTH-1:0]         Ic223d7941250d739ce9bb0ae5013646e;
wire [fgallag_WDTH-1:0]         I95eaa4ac5199ebbb06f780d1376062ec;
wire [fgallag_WDTH-1:0]         I41f34c28805f2653586d89312f73237f;
reg  [fgallag_WDTH-1:0]         I1ef9b548b943a1f2012b91c7e0b445f2;
wire [fgallag_WDTH-1:0]         Ib40ccfdb9ea28f333a7cc67f2446c923;
wire [fgallag_WDTH-1:0]         Ie2031e8a9632f0b98f617232f7c462e6;
reg  [fgallag_WDTH-1:0]         I88b6d7894d82ff394e89c7471c80dd5b;
wire [fgallag_WDTH-1:0]         I507515355429e697cd5496809aa03cfb;
wire [fgallag_WDTH-1:0]         I9d706a29e764935ac3cabdac4e95af1d;
reg  [fgallag_WDTH-1:0]         Ia5fc7e1f991f30042b848888a546534b;
wire [fgallag_WDTH-1:0]         I6bcc3a323e67f95eb4bf28a0704d3c50;
wire [fgallag_WDTH-1:0]         I7a2e1620640d2060cbb0a1bef5eb79c0;
reg  [fgallag_WDTH-1:0]         If699df4c8261ebce5c5d1aebe062cd61;
wire [fgallag_WDTH-1:0]         I55e3a2566ef3ac257021a294376be634;
wire [fgallag_WDTH-1:0]         I2795513c5d99dc8e09be4bebb4d12944;
reg  [fgallag_WDTH-1:0]         I19338369553e96bb2476d80fe84dec3e;
wire [fgallag_WDTH-1:0]         I40f10dc3289ea8a59f593f62066aaff8;
wire [fgallag_WDTH-1:0]         I03cb6aeff54e7e9e2ee809f8bea621bc;
reg  [fgallag_WDTH-1:0]         I9844ff02042cbc04dd5f4179908bbb2d;
wire [fgallag_WDTH-1:0]         Ieeabde5600d81208346ebd50d4a95d83;
wire [fgallag_WDTH-1:0]         I78c43fed329002e5ab9a0e429fb3b769;
reg  [fgallag_WDTH-1:0]         I89cc6a060b714985b24f724adc782e7b;
wire [fgallag_WDTH-1:0]         Ibb9220dcdd6d7fc2b6d6ca5f4cc93a8b;
wire [fgallag_WDTH-1:0]         I639755c3c20317c18359e96fce8e2f2e;
reg  [fgallag_WDTH-1:0]         I39d94ce7fbe37a74404e0043060441ed;
wire [fgallag_WDTH-1:0]         I05a3aebc90966144a6809e460d6ceda1;
wire [fgallag_WDTH-1:0]         I68c7cb0d5275b576e4021c8aedda4646;
reg  [fgallag_WDTH-1:0]         I0a1c9a8d59dbcffd6847f3a65107c407;
wire [fgallag_WDTH-1:0]         I7e3150622eb318e94f99b36016ac7d2f;
wire [fgallag_WDTH-1:0]         I2bd974f363231ecfaa9ef8d018a02936;
reg  [fgallag_WDTH-1:0]         I2328556c467a9e639f2b6ba1d0cb99b7;
wire [fgallag_WDTH-1:0]         Ifb146b2073d447377a1b21fe21baa4da;
wire [fgallag_WDTH-1:0]         I675d5b900c6a4bbdb8f14db50b873893;
reg  [fgallag_WDTH-1:0]         I5c9d75d6431d69db1abe412e591000a7;
wire [fgallag_WDTH-1:0]         Ifa5048ac43025e9cdf3f3436c37bb835;
wire [fgallag_WDTH-1:0]         I36b68c4fcf7a2adafce004ec0e231209;
reg  [fgallag_WDTH-1:0]         I8dc3dcdefc85b6ff8ecfa09cfc7e69fa;
wire [fgallag_WDTH-1:0]         I837ba4049e4973924e51d642f7f481ad;
wire [fgallag_WDTH-1:0]         Iea5c378e0635e3bb31343988c4dc6259;
reg  [fgallag_WDTH-1:0]         I69f6c909ea6b207c200b154e00e13a05;
wire [fgallag_WDTH-1:0]         I2910e5e74ca008b7e5502d787cb88a6d;
wire [fgallag_WDTH-1:0]         I2edf197a22f055871ed9b54f9e1a874a;
reg  [fgallag_WDTH-1:0]         Id365c9f8f7f97c777bd5da0ce9490511;
wire [fgallag_WDTH-1:0]         Ia24816d601e29172628cad0c364b47e9;
wire [fgallag_WDTH-1:0]         Ie80e559352812ffe4d9cf6006af19e85;
reg  [fgallag_WDTH-1:0]         Idf0206d2ad2bdef7db1d30a2d715cc6a;
wire [fgallag_WDTH-1:0]         I8f99af880f329241cfc9616ff9859091;
wire [fgallag_WDTH-1:0]         Id2f23da93344ae523d495478dd559ded;
reg  [fgallag_WDTH-1:0]         I07d1c54431eed887554a136f15f86d22;
wire [fgallag_WDTH-1:0]         Iea7c2970a7d80c55c1a6d6933c6c81c9;
wire [fgallag_WDTH-1:0]         If18e431ab87f137467f6f87e40b9c27e;
reg  [fgallag_WDTH-1:0]         Ic16809a3c82787ed88819fc9e9613f85;
wire [fgallag_WDTH-1:0]         I75a12697a4ee6de46fc098b0f02b8349;
wire [fgallag_WDTH-1:0]         I3f5b5d6b646070d84f2fb963f3824ce1;
reg  [fgallag_WDTH-1:0]         I1613ae89442495e703a52e65b8a0bf9f;
wire [fgallag_WDTH-1:0]         I623d1f0b6829caf5dc0f0eab0ca47f74;
wire [fgallag_WDTH-1:0]         Ie964e5a463904ac52c4529ffb3ebaf65;
reg  [fgallag_WDTH-1:0]         I6089da825af433e847c0b1bb9ff7d373;
wire [fgallag_WDTH-1:0]         Ieabf207f10f7df1e9059f1e953d7b399;
wire [fgallag_WDTH-1:0]         Ia74858d5df6a76635e6ba60d0b1a63ea;
reg  [fgallag_WDTH-1:0]         I6aa7fccf4e225fa70063fd24dab74e6b;
wire [fgallag_WDTH-1:0]         I1399b55530e343bd85606e7c7529d453;
wire [fgallag_WDTH-1:0]         Id9c69999bee621002fa9b387aa809dc5;
reg  [fgallag_WDTH-1:0]         Ibe2a5f680405f233256b6fd806b72ae5;
wire [fgallag_WDTH-1:0]         I39ee898ed8a8af64552e1aa145437310;
wire [fgallag_WDTH-1:0]         Ie9e8ae352a1699484f85ae1e7b7f9246;
reg  [fgallag_WDTH-1:0]         I662d408ffd8fb9f249e531a167161429;
wire [fgallag_WDTH-1:0]         I0af241f9f65af3bff2bb0d69977bb0c6;
wire [fgallag_WDTH-1:0]         I5a006c73dcb7807d5943857199cc3535;
reg  [fgallag_WDTH-1:0]         Ie95b8a5c2da6c0877d49c646c194f5b7;
wire [fgallag_WDTH-1:0]         I9de68705b5430023d2eb5554370bb188;
wire [fgallag_WDTH-1:0]         Idfb53869ea5692adddb6f7452d44effa;
reg  [fgallag_WDTH-1:0]         If940f33461f5e297e158db54f6aad610;
wire [fgallag_WDTH-1:0]         Icdf7ba01c4813abe3cfa760f2d8d5c84;
wire [fgallag_WDTH-1:0]         I0d11a8980f8fd7aadc8e48e62a653aa6;
reg  [fgallag_WDTH-1:0]         I54aa9d4c6333d94970eae97aeb3603fa;
wire [fgallag_WDTH-1:0]         Ia6b995eb6bbaad8a638c80d587d45ab9;
wire [fgallag_WDTH-1:0]         Ib843721cd2106b7e5cc21812aeb374eb;
reg  [fgallag_WDTH-1:0]         Ib82fc62720e6346e1c05cc33d596447e;
wire [fgallag_WDTH-1:0]         I75c2987dcebc9cdca578aeebec96fccc;
wire [fgallag_WDTH-1:0]         I400d30374ae90fa066db0f5a29195e4e;
reg  [fgallag_WDTH-1:0]         I24873624848b61f313865e10e77e35c6;
wire [fgallag_WDTH-1:0]         I6fab90e9a0f606d7c26346c89c6f1d47;
wire [fgallag_WDTH-1:0]         I49316949f603c233556dfe520b9e1a61;
reg  [fgallag_WDTH-1:0]         Icc3915d8325c22fc172f731553798fef;
wire [fgallag_WDTH-1:0]         Iab2f70a1d3093b3194e9047a8fe8e487;
wire [fgallag_WDTH-1:0]         I57c335ac00303b6df3bb5bc5a1b1bcb6;
reg  [fgallag_WDTH-1:0]         I93b9837e63103431a0fdaf319a465c90;
wire [fgallag_WDTH-1:0]         Ic84b6224be8eb8eefc9ad9bcc2280291;
wire [fgallag_WDTH-1:0]         I177fce9af9d7a8e9e9dfe423c8abe225;
reg  [fgallag_WDTH-1:0]         I91237af3aa2af551dbbc626bb701215e;
wire [fgallag_WDTH-1:0]         I64a0e60fdcc93d84606774196b2b7598;
wire [fgallag_WDTH-1:0]         I335535f77c13df799b6e5f9613607a9b;
reg  [fgallag_WDTH-1:0]         Ib254d9701567f642d3586641edf85128;
wire [fgallag_WDTH-1:0]         Iaa6a4f3826d87e43dd3213dc5083184b;
wire [fgallag_WDTH-1:0]         Icbe54351ad1360193ea28dc76e073f23;
reg  [fgallag_WDTH-1:0]         I25c50067a62d2b3599d15f12f89d384e;
wire [fgallag_WDTH-1:0]         I94fd5b790a9dceab1b4b3f1b5e30a0d9;
wire [fgallag_WDTH-1:0]         I812a6ce8adb2ef9a2a9eb7e7e8cc96f1;
reg  [fgallag_WDTH-1:0]         I238be7f0e4a209a6b4201a024c8aed82;
wire [fgallag_WDTH-1:0]         I9c8c1d22021bbe798b1863ae1dfc3965;
wire [fgallag_WDTH-1:0]         I87a99623e8305e331ca590dc62df5252;
reg  [fgallag_WDTH-1:0]         I233f5ddadd45c0df2108ea6c1d634f3c;
wire [fgallag_WDTH-1:0]         I870366e9c3b29c1683a7528f4b5d5329;
wire [fgallag_WDTH-1:0]         I130df8a2e7e3e33055f2f2997e6d5716;
reg  [fgallag_WDTH-1:0]         I87a320ddaa1478146ff6e519dc65c40a;
wire [fgallag_WDTH-1:0]         I066db3b79f8b4581f96567d943a7e7db;
wire [fgallag_WDTH-1:0]         I07ee1ac328d24e8fa9862659903fd379;
reg  [fgallag_WDTH-1:0]         Ibf03d6940c0a38bef038a28b6a7b625d;
wire [fgallag_WDTH-1:0]         Iabd6f58c4760c939dfd58e4f426bcab9;
wire [fgallag_WDTH-1:0]         Idd74d5e61d5397193aaf3cdb96dbc84b;
reg  [fgallag_WDTH-1:0]         I90942470e2057e50ce4f5745ed68b81c;
wire [fgallag_WDTH-1:0]         Ia3505661cb9b7eacbd47774346d12f5b;
wire [fgallag_WDTH-1:0]         Id74f690142fb1e4a04fa3dca841979a6;
reg  [fgallag_WDTH-1:0]         I77fbc3f3b65962b610e39f4b085ecb7e;
wire [fgallag_WDTH-1:0]         I4e7245fc882e3e284d8c152c8998b028;
wire [fgallag_WDTH-1:0]         I8327851510864c943e64c3d22b456152;
reg  [fgallag_WDTH-1:0]         I701845efaf1b02aefa381d4f6b45c401;
wire [fgallag_WDTH-1:0]         Ibe962754759204890883a6de0993a64b;
wire [fgallag_WDTH-1:0]         I4f37cf4b922e288365376a45753c4a38;
reg  [fgallag_WDTH-1:0]         Id446ddfd713c6e1592c562cfb123ea8b;
wire [fgallag_WDTH-1:0]         Id2ef1e193163adc702763541f37fec4d;
wire [fgallag_WDTH-1:0]         If50168d2535d752dd95301bfe723db9a;
reg  [fgallag_WDTH-1:0]         If4f752779d27392e7536565d425bce25;
wire [fgallag_WDTH-1:0]         I8a925721cf106d4e6ca1f69bbc2f53d4;
wire [fgallag_WDTH-1:0]         I6eb5641a21e34b4ced1cf124c3f23646;
reg  [fgallag_WDTH-1:0]         If112169057d6293326a56443ac3cf517;
wire [fgallag_WDTH-1:0]         Ib97671e4daa1b606aa01c5e8f753a9e8;
wire [fgallag_WDTH-1:0]         I94da98c2f9e0c8be8ab8f23a2a10095b;
reg  [fgallag_WDTH-1:0]         I78f727f8d85b5d7f0ffa57f02538f939;
wire [fgallag_WDTH-1:0]         Icdd0962fd06355a7dcbb491543eb9cb6;
wire [fgallag_WDTH-1:0]         I339ec0bef37cb2e72e8e8795686da0c4;
reg  [fgallag_WDTH-1:0]         I01ec629f60c17c2251f977205234cd44;
wire [fgallag_WDTH-1:0]         I003f9dc1b83f386f070b0a2e8c7ce4f4;
wire [fgallag_WDTH-1:0]         If7c621d8183ce83092644a1d80d6c77b;
reg  [fgallag_WDTH-1:0]         I23f774adb64807c0edaa9941c75651b6;
wire [fgallag_WDTH-1:0]         I66e8ad34c764833f038cff700a237fcb;
wire [fgallag_WDTH-1:0]         Icb4d6012447eb0d6bfa8e8b3f88f0ff9;
reg  [fgallag_WDTH-1:0]         I2361ef4fd70e4c05b25289d0845564c4;
wire [fgallag_WDTH-1:0]         I614bddda696787a552e28cfaa81a3aa3;
wire [fgallag_WDTH-1:0]         If7c3b54bc0cce4eecf8f55fcf4a5a588;
reg  [fgallag_WDTH-1:0]         Ic3067b434ca17be7bad595e1f9b822c5;
wire [fgallag_WDTH-1:0]         I38c22e6b7c066be10ec1f8929dbf88f9;
wire [fgallag_WDTH-1:0]         I1ffe02eedf41df8b947a285adc220fea;
reg  [fgallag_WDTH-1:0]         I3546ddbae9c9db4517802db56cee35f0;
wire [fgallag_WDTH-1:0]         I245816ec4a0392af2cfa4b44a4e93610;
wire [fgallag_WDTH-1:0]         Icd8c721f78cfbefbf25c2e094927401a;
reg  [fgallag_WDTH-1:0]         I35e91092ed503831ed818f36a1ce1537;
wire [fgallag_WDTH-1:0]         I83253182662d56779685c9742f55789f;
wire [fgallag_WDTH-1:0]         Ie139a6a80ab0051c5d951103b1554338;
reg  [fgallag_WDTH-1:0]         I973f185cf29e13193abf0108d4faa9d1;
wire [fgallag_WDTH-1:0]         I963a4391dba3d12756b89dda1e962c3f;
wire [fgallag_WDTH-1:0]         I993fd34b89fe9b0af3348cdd91ecf025;
reg  [fgallag_WDTH-1:0]         Iee58b0442a6cccf0990ebb551b47fa92;
wire [fgallag_WDTH-1:0]         Ie959690f46f82cbb15ae0cee69f3135f;
wire [fgallag_WDTH-1:0]         Ib5d321981c2997b3635fd0b342993d38;
reg  [fgallag_WDTH-1:0]         I2cb3207a5c1b25386ac7eb532955f260;
wire [fgallag_WDTH-1:0]         Ic475c578935fa69db2b1c834539750af;
wire [fgallag_WDTH-1:0]         If1660e858bdb3b0c8a4c1f93f4fe037a;
reg  [fgallag_WDTH-1:0]         Icd4f07bc30c66f7f5b431ed97e7ac7b6;
wire [fgallag_WDTH-1:0]         I4f9bc0f2aeafb89fbaa0d0af7dbda06a;
wire [fgallag_WDTH-1:0]         I7d9ab0daacce00542083a30a35297207;
reg  [fgallag_WDTH-1:0]         Ifec6f3a1e10144acb320d5d502ed1ea3;
wire [fgallag_WDTH-1:0]         I393fa73117dcbf1fb1b74ea1fc7e6c99;
wire [fgallag_WDTH-1:0]         I9761f2282bcb9637892cf898b928126c;
reg  [fgallag_WDTH-1:0]         Ic87bff64a597e6d02583041b552328ee;
wire [fgallag_WDTH-1:0]         I95836c571386b3b6de07c9195932fe22;
wire [fgallag_WDTH-1:0]         I25de2ab105b6cdb0e30ca97822109fbd;
reg  [fgallag_WDTH-1:0]         I489f21ef8243ef8caa1c29f034c3e2ac;
wire [fgallag_WDTH-1:0]         I6dd6f9abc962974c292d22f17a21a936;
wire [fgallag_WDTH-1:0]         I23c14408deedeecba4753f182549adf7;
reg  [fgallag_WDTH-1:0]         I773901563077961acada85962209d68a;
wire [fgallag_WDTH-1:0]         I9f9e6bc8d2cc6e41813d42ffcd5cff01;
wire [fgallag_WDTH-1:0]         Id208387ab734f8ccfaf1567e6b00a4a6;
reg  [fgallag_WDTH-1:0]         Ifbd176fe3e78bc2dc2e0e77ba3ccd2d0;
wire [fgallag_WDTH-1:0]         I2ba75ccf97b5caf5aa676a9e3c42a366;
wire [fgallag_WDTH-1:0]         I54e43b8da49648867403cf839e87a9ec;
reg  [fgallag_WDTH-1:0]         I53f68a4cb81c71ee7bd6f61171b7478d;
wire [fgallag_WDTH-1:0]         I006699f0e016e7022b2706751965c42c;
wire [fgallag_WDTH-1:0]         I66c8b8649e7997b7e4c9c17f7c0b17b7;
reg  [fgallag_WDTH-1:0]         I7568ec59f1359bedce86dbc6af50df71;
wire [fgallag_WDTH-1:0]         I66d5992f4f39337782cfbbb9fec3b2c8;
wire [fgallag_WDTH-1:0]         I9a0093065fb4cf517f1e7b75b3080b1c;
reg  [fgallag_WDTH-1:0]         Id2bf82d6bf0a201f80a58357038a0992;
wire [fgallag_WDTH-1:0]         Ie5f503c91ddf6eff2b9645e6e3c22b2e;
wire [fgallag_WDTH-1:0]         I72d18b26784448b5514e66251bb19ebd;
reg  [fgallag_WDTH-1:0]         I22442354ca2b77306f25839ce6124699;
wire [fgallag_WDTH-1:0]         Ieb7e6a2425e93a2b96a94f0e2c4442c3;
wire [fgallag_WDTH-1:0]         Icec022a0de167257d08e0b2beb6ba8f5;
reg  [fgallag_WDTH-1:0]         I71a5c2876a07d8edd001ef2d108e59c1;
wire [fgallag_WDTH-1:0]         I4a0483f2d2585cd44fe35191d7cd88b1;
wire [fgallag_WDTH-1:0]         I3d8a7850f0080b0d6068d58837e3294f;
reg  [fgallag_WDTH-1:0]         Iaf333aa6b135927cf1ad1f76298ccd63;
wire [fgallag_WDTH-1:0]         I00e8b3cde14889fcb0b40dc5582a58f9;
wire [fgallag_WDTH-1:0]         I26b947511e25e51f1bb9728c169e7e64;
reg  [fgallag_WDTH-1:0]         Ia71cfd8cf9bea4e600ea204e41271c7d;
wire [fgallag_WDTH-1:0]         Ib53dbb62231f729a278d2afa3acffdbf;
wire [fgallag_WDTH-1:0]         I8baf26027cc707ae93b6c74e2af5f207;
reg  [fgallag_WDTH-1:0]         I164b032929ac2b8cf1a6672859639a30;
wire [fgallag_WDTH-1:0]         I5503d6011d58dfa4e1ec524eb1875c7d;
wire [fgallag_WDTH-1:0]         I9902253554855a3d12ceaf47f6cc5569;
reg  [fgallag_WDTH-1:0]         I2ef0447f5c64fd5c65e23c16069a62ef;
wire [fgallag_WDTH-1:0]         Id86fbda00d923c29c99b4a9fe52d513a;
wire [fgallag_WDTH-1:0]         I81ab0ce0526dd851c51d5d42f807e62d;
reg  [fgallag_WDTH-1:0]         Ide7008ee7f1fba156dc6145b3505e553;
wire [fgallag_WDTH-1:0]         I3ba6e9f7d7fa98ad776299f8cd8a8363;
wire [fgallag_WDTH-1:0]         I51dc4acb242b33bb123f8b106aafbc93;
reg  [fgallag_WDTH-1:0]         I129a7ced6bc6f48f20fa552e2519925c;
wire [fgallag_WDTH-1:0]         I67b512efbaf9c063a4ac75cb97a8abdb;
wire [fgallag_WDTH-1:0]         I32ca8b2806bf397557167b133d1411ab;
reg  [fgallag_WDTH-1:0]         I67123cf825352e52cf0158060ad69a13;
wire [fgallag_WDTH-1:0]         If5f5eecf512463544c8b2419c0a58779;
wire [fgallag_WDTH-1:0]         I5c39fac168568808f33fc6be5eec66a7;
reg  [fgallag_WDTH-1:0]         I09923d784a9f9625a37221f639537941;
wire [fgallag_WDTH-1:0]         I81cdc8b54bc7f98798713985e8f4553e;
wire [fgallag_WDTH-1:0]         If355236b8b8375ad095cc46a373ad4d6;
reg  [fgallag_WDTH-1:0]         I5947be93fdb18bf0ad341fb826c9e6d7;
wire [fgallag_WDTH-1:0]         I35bb2eb0cb589f694001ba1509cbf7f8;
wire [fgallag_WDTH-1:0]         I31fad95729e24c7724a73285e966684f;
reg  [fgallag_WDTH-1:0]         I08621ee033cd49702ad08af4d31eb999;
wire [fgallag_WDTH-1:0]         I3bf8f19c98c78f8e1c315e75a533bb1c;
wire [fgallag_WDTH-1:0]         I0415d9d3687656d7a07ea2c12ba505d1;
reg  [fgallag_WDTH-1:0]         Id5eca60b22d3835119571fe4b1a03479;
wire [fgallag_WDTH-1:0]         I71cbdcd6e3a873851e9084bc9dcd99bd;
wire [fgallag_WDTH-1:0]         Id54f584cdc590112180e9000e1d015a1;
reg  [fgallag_WDTH-1:0]         I7267ba2b9cb511a48a3a7044e854f7da;
wire [fgallag_WDTH-1:0]         Iebad2e3d84bae3d4807badae823aec52;
wire [fgallag_WDTH-1:0]         If9930e999d72a139c345aeb1c33e51c1;
reg  [fgallag_WDTH-1:0]         I5893fa21ec8bbdcea9677cc12fc4057a;
wire [fgallag_WDTH-1:0]         I054f07cdf6a44100034c7e2fb438055f;
wire [fgallag_WDTH-1:0]         I28e9624edb8f59290eba51c87f2a88cc;
reg  [fgallag_WDTH-1:0]         I564896fe01ec799a0fbe790473753559;
wire [fgallag_WDTH-1:0]         If3b82307d1ad78e262f76ba9b711e1a6;
wire [fgallag_WDTH-1:0]         Ie6c99d8fe1a105832500bf8a722c82c7;
reg  [fgallag_WDTH-1:0]         If279ab7c515c4039c8272b913c2fa107;
wire [fgallag_WDTH-1:0]         I0f40c8301521c136b3ede2cc9e8352a3;
wire [fgallag_WDTH-1:0]         I24307c47884babba3b0a16a1791c674f;
reg  [fgallag_WDTH-1:0]         Ib61705ff5820f531eb17c40ed05f6ec3;
wire [fgallag_WDTH-1:0]         I3615a34cbf1646a7cd0f1da43d62faa5;
wire [fgallag_WDTH-1:0]         I2951bad4b57a2ad6715844998c491ec7;
reg  [fgallag_WDTH-1:0]         I50149e5de41ca2998c4e8cc4b19e166b;
wire [fgallag_WDTH-1:0]         I0bbd697ad8d3877570ab9e200e66164a;
wire [fgallag_WDTH-1:0]         Ie0149abcf22aeff58be4cb418f477239;
reg  [fgallag_WDTH-1:0]         Id40cac3272643f3f91b73c6aa1740f3b;
wire [fgallag_WDTH-1:0]         I298f7389a7fd8e927b7e3354f0d32344;
wire [fgallag_WDTH-1:0]         If8ec8dc5888438922c6074ff23eb42c7;
reg  [fgallag_WDTH-1:0]         Ic63eee2d700493c41ee2d186ff7111b9;
wire [fgallag_WDTH-1:0]         I9960d39fce3c5b9945965dedac46dfed;
wire [fgallag_WDTH-1:0]         If969c721b9636b840193a85d8946fc32;
reg  [fgallag_WDTH-1:0]         I51de42598e0df4a76cf7b02c61ae9550;
wire [fgallag_WDTH-1:0]         I02f48e93599dc91bb24a144a0ef1a933;
wire [fgallag_WDTH-1:0]         Id6dec5f563e485414043770af559ec76;
reg  [fgallag_WDTH-1:0]         Ia89a1a58f6327ee3c105cae860942171;
wire [fgallag_WDTH-1:0]         I7e31af1959a0374af6c2767e4837c566;
wire [fgallag_WDTH-1:0]         I79ae237d2105b50c92b8507272bcbd4e;
reg  [fgallag_WDTH-1:0]         Ib149a5872e31cd5df77b66298b4aad12;
wire [fgallag_WDTH-1:0]         I8d18e2ecaf2bda4a0ba47d9782e9917a;
wire [fgallag_WDTH-1:0]         I9ea4ebd1f6cea81da598f16b5a7c31f4;
reg  [fgallag_WDTH-1:0]         Iaa16c14572ad0442eb3c58a97bef5ada;
wire [fgallag_WDTH-1:0]         Id0a13655f967dfd3000b8dcf4a57f555;
wire [fgallag_WDTH-1:0]         Id7b8f8df1818623e7a9e897e019a09e7;
reg  [fgallag_WDTH-1:0]         I88d5d48e05b1c9a6d8060f58917e3834;
wire [fgallag_WDTH-1:0]         Ibf384c0b998b5a5f7808c54292c6b844;
wire [fgallag_WDTH-1:0]         Ia5e1a46c7d21e79ef859b788b27ee3d1;
reg  [fgallag_WDTH-1:0]         I4269e18c2df4d39c683ffb7d01a08322;
wire [fgallag_WDTH-1:0]         I58b8202ae510e96b4f6ae334f3b282c6;
wire [fgallag_WDTH-1:0]         If5b0270fa354f64b8b58e5f02353daa4;
reg  [fgallag_WDTH-1:0]         Ia29017fa9327fdaa7c10b2797f8aa6ec;
wire [fgallag_WDTH-1:0]         Icbc75d6e4d0bcc42cdf813529b017e0e;
wire [fgallag_WDTH-1:0]         Ie800c32198a9d6181225f2274b301d9d;
reg  [fgallag_WDTH-1:0]         Ia142ac799256541fe33f898a6a31dd71;
wire [fgallag_WDTH-1:0]         I6fa1835a8e7f8ea435c4515b1c059cc9;
wire [fgallag_WDTH-1:0]         Id596782860b623f79a8fd0e83712d9d0;
reg  [fgallag_WDTH-1:0]         I4c039794243933a9bb7ad6db7eda6a87;
wire [fgallag_WDTH-1:0]         Id3984a3dd1009c9c76347b9843f27b25;
wire [fgallag_WDTH-1:0]         If5a41054200c97e01b9132f7c7ff9793;
reg  [fgallag_WDTH-1:0]         I0debb3ed4f9540c162cd525588e0ae3f;
wire [fgallag_WDTH-1:0]         Id5fd757abdc0b2e1b1d4c5dab96ee08a;
wire [fgallag_WDTH-1:0]         I2cf304c8f8efef74593929b1bea0bf91;
reg  [fgallag_WDTH-1:0]         I681eed68ee814fb18fd794207d9266e1;
wire [fgallag_WDTH-1:0]         I98ab1b82b2991b4cb3bec530711bdc43;
wire [fgallag_WDTH-1:0]         Id0b597aa1dc456b83d4e38147c97a9fb;
reg  [fgallag_WDTH-1:0]         Ic260784b8910f5a0483afee9b68efb31;
wire [fgallag_WDTH-1:0]         I610d0ed6f55a4906aac1be5823358392;
wire [fgallag_WDTH-1:0]         I318a691d3ffd634a1c5c362d5b3a8c34;
reg  [fgallag_WDTH-1:0]         I22cd2d30a7684002cacca4deae4c95a0;
wire [fgallag_WDTH-1:0]         I2ed0ad73f73f9f4e1b7ec38af320ee4d;
wire [fgallag_WDTH-1:0]         I881c34f97e2d2f4765cf3cd7cde53c7f;
reg  [fgallag_WDTH-1:0]         I136b4136d582f9fad21f90297cfafea3;
wire [fgallag_WDTH-1:0]         I3dfc4dd447cd1f4e40506f516c106861;
wire [fgallag_WDTH-1:0]         I922d1ac78df6c82308d2028527f8f56c;
reg  [fgallag_WDTH-1:0]         Id8d6be9677d3b0ceca26b3b671757c2c;
wire [fgallag_WDTH-1:0]         Idfeea354b3f9ca8c671851fd90f4e1bc;
wire [fgallag_WDTH-1:0]         I49dbef91e0572ad9296838e769edf0c3;
reg  [fgallag_WDTH-1:0]         I6a93f928c104ea211dcc8a461506327d;
wire [fgallag_WDTH-1:0]         I415d8306edb869fc838eb518aad75168;
wire [fgallag_WDTH-1:0]         I8819e4519e4930d300f5536af5d62a94;
reg  [fgallag_WDTH-1:0]         I240da147648bec33195a5f5c273fc6f4;
wire [fgallag_WDTH-1:0]         I1dc6b2aef1bb326c3d5c19f97a2e1d4f;
wire [fgallag_WDTH-1:0]         I4779a6c85288e6dba977cedd1cd3cb6b;
reg  [fgallag_WDTH-1:0]         I55494d0e8454e3cbb4158559e0d29984;
wire [fgallag_WDTH-1:0]         Ie2f47a06ca4b6d5823cbbe099f5de0f0;
wire [fgallag_WDTH-1:0]         I934d36f3afd37afdaad46c93f45a044c;
reg  [fgallag_WDTH-1:0]         Ied3cc579b3cf126081acf8e1117007cf;
wire [fgallag_WDTH-1:0]         I55b7a58384e50ade254c3c8934c290f6;
wire [fgallag_WDTH-1:0]         I2667428380ad21221430252aa00402bf;
reg  [fgallag_WDTH-1:0]         I76140bdc374dd6031097575fd231b468;
wire [fgallag_WDTH-1:0]         I53bf5dca5911aec50866be5a720d4aa2;
wire [fgallag_WDTH-1:0]         I257185648f29565e2259890a6a70583a;
reg  [fgallag_WDTH-1:0]         I650345d21e5c2e7a9bf1810630161089;
wire [fgallag_WDTH-1:0]         Ie57f78d4c002e69e0e92b25bad752d3f;
wire [fgallag_WDTH-1:0]         I49a61c916eb52d0bfd08700d087d379a;
reg  [fgallag_WDTH-1:0]         Ie852635f073dc918e7b1075ffad46f24;
wire [fgallag_WDTH-1:0]         I2ac511a908c9973254672fd38cabccd3;
wire [fgallag_WDTH-1:0]         If180a1b31f53c672e4f05b2aeca3caba;
reg  [fgallag_WDTH-1:0]         I9ec80c14eb5f0f305e1a9e6107a6001e;
wire [fgallag_WDTH-1:0]         I8f06d78dd2e6be736f4e4f41fadf130d;
wire [fgallag_WDTH-1:0]         I335057378d9ae46b1e1442fd341fabad;
reg  [fgallag_WDTH-1:0]         I80ba56447ab19b33610c23105b0b1637;
wire [fgallag_WDTH-1:0]         I65450e396e33720967b7a6271e3a70e1;
wire [fgallag_WDTH-1:0]         I3027f4cba09ab3eee29cf9b34ed27ae4;
reg  [fgallag_WDTH-1:0]         Ib9132d9fa7180c3fcbacb7c570d6b0f2;
wire [fgallag_WDTH-1:0]         I876c6361d2164d03cad2ffc8bf920ac0;
wire [fgallag_WDTH-1:0]         I9ac1c5487994b853d666af93d35c82cc;
reg  [fgallag_WDTH-1:0]         I01621f113f636a9caf9b5ca0bb20ef77;
wire [fgallag_WDTH-1:0]         Id3b8e1157a3e9eea4d210f466740f673;
wire [fgallag_WDTH-1:0]         I099f1e1b4eb55718dd73dff7efc16ae9;
reg  [fgallag_WDTH-1:0]         I3eeddb549c6e1f07469c0e0dca68be92;
wire [fgallag_WDTH-1:0]         I6973de59fb6014d7c4bf5b982cddc4d8;
wire [fgallag_WDTH-1:0]         Ie9ebb06f41fbc042867ee14d8f4090f2;
reg  [fgallag_WDTH-1:0]         Ibe664dd203ed4162abcd36eb8d57bfa6;
wire [fgallag_WDTH-1:0]         I26cb99c4cc37be5f52dfeeca60d5d102;
wire [fgallag_WDTH-1:0]         I2647305e100a9fb38fbf290f12778d49;
reg  [fgallag_WDTH-1:0]         Ia66176893fe306ecfb415d948c50486d;
wire [fgallag_WDTH-1:0]         Ie9835b1d512d9c9c4f2801956fbf13cb;
wire [fgallag_WDTH-1:0]         Iae4b5e5348101abc4640c84686ddad69;
reg  [fgallag_WDTH-1:0]         I8bd4210dcbfc1956381b460fd9ef789b;
wire [fgallag_WDTH-1:0]         I89057e4e979b903ae1f10f9dd2f196fe;
wire [fgallag_WDTH-1:0]         Ibeba1d51f76197f960672ea90dabfb75;
reg  [fgallag_WDTH-1:0]         I1ba6328ea9cb7cebcce47d5407d0eae7;
wire [fgallag_WDTH-1:0]         If1299e6b34cd1f2239d64ade23f33f01;
wire [fgallag_WDTH-1:0]         I83ebb6a41c9d866a8ff3fe3fa0b5321f;
reg  [fgallag_WDTH-1:0]         I9e79c17bd782bb7981b4a3623baf96a1;
wire [fgallag_WDTH-1:0]         I3f106ef1876021bb3cc5866d2b5698f4;
wire [fgallag_WDTH-1:0]         Iedc551659ac328435c906b5748c9790f;
reg  [fgallag_WDTH-1:0]         I7c6f64d73ff9c6e7f2ed69713e056a2b;
wire [fgallag_WDTH-1:0]         If6cb9fec3dc380f1c4894bccfa35b33c;
wire [fgallag_WDTH-1:0]         I95e1540f2a2eadf6fb80e3519a1d9d5c;
reg  [fgallag_WDTH-1:0]         I00b962a9bf04b62244591051d2dfdbbd;
wire [fgallag_WDTH-1:0]         I313980f8406e9f26d5eaa53270a23b9e;
wire [fgallag_WDTH-1:0]         I3587e6334c7c3f23bee5675353bbeaba;
reg  [fgallag_WDTH-1:0]         I3a660b57588325989319701026f658e6;
wire [fgallag_WDTH-1:0]         I792b5aea212da69a9c18f5723e820432;
wire [fgallag_WDTH-1:0]         I4e71cbc9773ff4abc24804d39a64abf8;
reg  [fgallag_WDTH-1:0]         Ibae27cccf3f64e8653c1e244e940e421;
wire [fgallag_WDTH-1:0]         I98f245ec9b667dc065c9494c00ecdf88;
wire [fgallag_WDTH-1:0]         I884dc79c03a585814e9d058ef7669ed8;
reg  [fgallag_WDTH-1:0]         I27b89a5001312b2aa48fe385d8a52063;
wire [fgallag_WDTH-1:0]         I15254b39b6e136520a9497d8684f9d94;
wire [fgallag_WDTH-1:0]         I0b2b9b8f1d6c6d5c6c5a8bd883d3ea5c;
reg  [fgallag_WDTH-1:0]         Ic6a7476db711a812d146331c562ca7c9;
wire [fgallag_WDTH-1:0]         I6c8312a9d655f143a0b65d91907ce533;
wire [fgallag_WDTH-1:0]         I645a63009d5be827b30fa02df646c872;
reg  [fgallag_WDTH-1:0]         I01ca07fe91b5f1edf87300b3583e77c5;
wire [fgallag_WDTH-1:0]         Ie6df2f89b05947f6be3b64e3b4f23df3;
wire [fgallag_WDTH-1:0]         If4630c847d9890c2b93acbaa6c9bd392;
reg  [fgallag_WDTH-1:0]         I6da707fd74249175d1f68dccb66390c0;
wire [fgallag_WDTH-1:0]         Ia71232b0b468b729fa1262957cbe9faa;
wire [fgallag_WDTH-1:0]         I49c56ae29a27e764325a9dcacb99f907;
reg  [fgallag_WDTH-1:0]         I0ae62aae426b75b06d95c46baf33f08e;
wire [fgallag_WDTH-1:0]         If75d8d882c6afc3df62096486b8e5b80;
wire [fgallag_WDTH-1:0]         Ie5272faa6aabb6e8d0720cdb7ec98358;
reg  [fgallag_WDTH-1:0]         Iec512b5870f295a50921e7e0289a7d35;
wire [fgallag_WDTH-1:0]         I7ed551b891500784c827992eb53f9ef9;
wire [fgallag_WDTH-1:0]         I92779ca466dbced9070a774d84439921;
reg  [fgallag_WDTH-1:0]         I3aac84acd9d78070472b1cbc745c80a7;
wire [fgallag_WDTH-1:0]         I5b5a24fd7116acd8ad2161513848c6a2;
wire [fgallag_WDTH-1:0]         I037e8ab38d779544d25ca5a4bfadeade;
reg  [fgallag_WDTH-1:0]         Ibbb900f56de318bf6e65b49791835ef4;
wire [fgallag_WDTH-1:0]         Id7055f4e578533dbd25d0505f8e47f34;
wire [fgallag_WDTH-1:0]         I3001e26d13b0cca9bc53d24324ac44d4;
reg  [fgallag_WDTH-1:0]         I2c2ac1e722fba72c759f1d37b88a9a10;
wire [fgallag_WDTH-1:0]         I9c78f3a2aa3986718caf8e70d4d939d4;
wire [fgallag_WDTH-1:0]         I933465899e56523ce1c470cad8dbd229;
reg  [fgallag_WDTH-1:0]         Ida0a18f1b79aff4ddf0e8f7e27794674;
wire [fgallag_WDTH-1:0]         I2def789e23f8ea0edee6f58200144096;
wire [fgallag_WDTH-1:0]         Id8b135f08d0464f9e308e25b8df2eb1d;
reg  [fgallag_WDTH-1:0]         I9f2029db42c5a968b370587c958c8929;
wire [fgallag_WDTH-1:0]         I319c2cb3a815a6347511f0c398876a3c;
wire [fgallag_WDTH-1:0]         I938596dee81ba14870ee4acfabce5e7b;
reg  [fgallag_WDTH-1:0]         If5755f4f61a89d91a91188c17ff5dc5a;
wire [fgallag_WDTH-1:0]         I0603434655e30a66d4e00b2bc2c878c0;
wire [fgallag_WDTH-1:0]         I61599f00ae7d6964dd40c96edefd6f67;
reg  [fgallag_WDTH-1:0]         I4419d97c3174ee4610eb6ee9c06cb256;
wire [fgallag_WDTH-1:0]         Ia6f16190b83b661f68a7a217bb356bdc;
wire [fgallag_WDTH-1:0]         Ic847a85de8e8ba2df520b737ea004374;
reg  [fgallag_WDTH-1:0]         Ia964f83676273055e20a2f63c8fffa0d;
wire [fgallag_WDTH-1:0]         I68fc61dbee0900bd66be7c7f5aaf8825;
wire [fgallag_WDTH-1:0]         Ifb0f088bf5bbf1884e1f27ed9808c273;
reg  [fgallag_WDTH-1:0]         Iab4fbc811e87df1d1f5821ea732b6a93;
wire [fgallag_WDTH-1:0]         I4ddd7ecf84b4ee4a4b6290f3d362f190;
wire [fgallag_WDTH-1:0]         I8705aa11e5ada7ec6e5431292d83fc54;
reg  [fgallag_WDTH-1:0]         I4fbefbb10724b0844c95e85495d4a87f;
wire [fgallag_WDTH-1:0]         I8e60b67eb6a187737de2717ebb95cf6c;
wire [fgallag_WDTH-1:0]         Ieaa7babedd5bfa1c8e1eb50d62ad9682;
reg  [fgallag_WDTH-1:0]         I717217d0b5a526f04c7f5ab0835dd5c7;
wire [fgallag_WDTH-1:0]         I7e17264500cb48d228c20542c40169cb;
wire [fgallag_WDTH-1:0]         I9eb9f7a6fe5932b574084bb18ce44e78;
reg  [fgallag_WDTH-1:0]         I235937b643e8f2848116dc76c43f47a7;
wire [fgallag_WDTH-1:0]         I6bddfc7b277ff042899fb2acd5625c5e;
wire [fgallag_WDTH-1:0]         Ic4b80e5673ad931188a2edfa1119e139;
reg  [fgallag_WDTH-1:0]         I7481f17d659cce5b4c72a68a9f6be67f;
wire [fgallag_WDTH-1:0]         I6daafbc7b14e2736b2a4e29c5f6fc5ff;
wire [fgallag_WDTH-1:0]         I5cdaf1ff24d7fb2bb4411b63a0a4488a;
reg  [fgallag_WDTH-1:0]         I5715c21c80992a61bff8aabc3f80415b;
wire [fgallag_WDTH-1:0]         I29df797d4c3ebd64fb088660bf89e922;
wire [fgallag_WDTH-1:0]         I7db6dcc03117fef703f20919a3c2ee89;
reg  [fgallag_WDTH-1:0]         I434e3216a615eb46be5c26ef914b9cd2;
wire [fgallag_WDTH-1:0]         I9418cc6766916bf1afc1f8a01feaad4e;
wire [fgallag_WDTH-1:0]         I3d2a8a166ccade50e320baaa68b40954;
reg  [fgallag_WDTH-1:0]         I918326ac0a744d234d74e2c08cf41eb4;
wire [fgallag_WDTH-1:0]         I90e1a5b43e93c02512a76c5cab15c5ad;
wire [fgallag_WDTH-1:0]         I3356737fddf6440f36fde442d29bb860;
reg  [fgallag_WDTH-1:0]         I966706d314f4c0a7ec842dd699d34926;
wire [fgallag_WDTH-1:0]         I26977fe4cdb2f9714fae2f12ca4a809b;
wire [fgallag_WDTH-1:0]         I13d6fc4a99a3a9989e655c417552fdb1;
reg  [fgallag_WDTH-1:0]         I5a7d246d88ef12e999f4bdee40e5a585;
wire [fgallag_WDTH-1:0]         I59775b68e199902c38d62e28cff01393;
wire [fgallag_WDTH-1:0]         I8a508ec5f2c2aaa05b632f422e67394f;
reg  [fgallag_WDTH-1:0]         Ic2dfaf65c4e17a8dcd55f766c314d6ef;
wire [fgallag_WDTH-1:0]         I9470ef82dad13754d8d061b5fd00a667;
wire [fgallag_WDTH-1:0]         I451fd82336efc778a51debf10f7cf325;
reg  [fgallag_WDTH-1:0]         I151831ba6bd0e162275c84815e3c0f12;
wire [fgallag_WDTH-1:0]         I62eb7a176351be84d086ce3c463214e8;
wire [fgallag_WDTH-1:0]         I76637de9be7c2c0dd0c324b4327a6184;
reg  [fgallag_WDTH-1:0]         I5a8f1675234ebed14d719344b530bbd7;
wire [fgallag_WDTH-1:0]         I106eb0d8f9ea92cda7bec4fe4aed6409;
wire [fgallag_WDTH-1:0]         I6e6d24ccb985ade6f058ce459592dfb0;
reg  [fgallag_WDTH-1:0]         I95dce76a8d0e729d40fb3f573cfc06ad;
wire [fgallag_WDTH-1:0]         Id0c12bc1a2139e57ea40c3254f30de7b;
wire [fgallag_WDTH-1:0]         If379a7696fdd0afebcb8ca169bb8f34a;
reg  [fgallag_WDTH-1:0]         I6c26c7918254426c18f2e747c91438c5;
wire [fgallag_WDTH-1:0]         Ib809a6099992799ce0235f22ce798c9a;
wire [fgallag_WDTH-1:0]         Idbd1062a6090858034185f1d5d503adf;
reg  [fgallag_WDTH-1:0]         I0414ead2472e42da8a271cb0bd1debf4;
wire [fgallag_WDTH-1:0]         I1a9be3897e044e9b24ac330ef3a20419;
wire [fgallag_WDTH-1:0]         Iea3c638b692d2540c1c8c81a6308673d;
reg  [fgallag_WDTH-1:0]         Ic6a6f5090470a76ddb7315c022ddc104;
wire [fgallag_WDTH-1:0]         I6e87b3400b7ddab94faf11c3910fa534;
wire [fgallag_WDTH-1:0]         Icd9e1d048d56d5d8557f80329bc6ffcc;
reg  [fgallag_WDTH-1:0]         I2a00ee56a5aa639f45eb3b1bdcffe81c;
wire [fgallag_WDTH-1:0]         I51e0ff0f52ca609663781545174b763d;
wire [fgallag_WDTH-1:0]         I6f0de2d570fa0245666c834b823e545b;
reg  [fgallag_WDTH-1:0]         Ibceb2b824cd4bc10bb06ee8adc693bd1;
wire [fgallag_WDTH-1:0]         I5c523df1fb2161ab4efd1c9b3e6b7aef;
wire [fgallag_WDTH-1:0]         Ief41e2502056d029a0c8bea8c052700c;
reg  [fgallag_WDTH-1:0]         Ia8b9f373fe68ac4cbca35e04376e3cca;
wire [fgallag_WDTH-1:0]         Ia307e5901694783f7761cdf724b767d0;
wire [fgallag_WDTH-1:0]         I7cd5df0d2845c7ed9f336a7940c7256e;
reg  [fgallag_WDTH-1:0]         I5d1a89e85f6609b469e73e15aeffcbc4;
wire [fgallag_WDTH-1:0]         Ia47164e8ba831b85e696e30ff59ceab1;
wire [fgallag_WDTH-1:0]         I5471bcc8bf4f4d0fab46d549b43113ef;
reg  [fgallag_WDTH-1:0]         I677fe06bad241bc8dd6a65a97f6db520;
wire [fgallag_WDTH-1:0]         Ic217af0cb9728801034fdcb273a577fc;
wire [fgallag_WDTH-1:0]         I599b8e0677efc1541283c2d7bf84809f;
reg  [fgallag_WDTH-1:0]         If3c0f892fd71eb0ed8d1f70b4b33450b;
wire [fgallag_WDTH-1:0]         Id5c8ea61025914f6e5a9b5eab9269261;
wire [fgallag_WDTH-1:0]         I4e4829b24a42e96e5c8399156aa61786;
reg  [fgallag_WDTH-1:0]         Ic65f0f75f56bf85122a89cdf07e98152;
wire [fgallag_WDTH-1:0]         I924ef8499a83579e3449bbac0994775e;
wire [fgallag_WDTH-1:0]         I1cda8d902f71f780775c85f38f9e799e;
reg  [fgallag_WDTH-1:0]         I41d22bafaf58e4a6de04640864653a16;
wire [fgallag_WDTH-1:0]         Ia8da4833c93e9ef6188709e7082092de;
wire [fgallag_WDTH-1:0]         Ic0b2c3e49d55853bc705021e5c0a2b06;
reg  [fgallag_WDTH-1:0]         I06a46b86f6edede0f5f72658a19910b7;
wire [fgallag_WDTH-1:0]         Icd8516e6bf231bce29ebefbc7c97bff7;
wire [fgallag_WDTH-1:0]         I6235ba2f129cfbcff36b368a39312bd7;
reg  [fgallag_WDTH-1:0]         I8591d0399594adacfeb006c5195c2c71;
wire [fgallag_WDTH-1:0]         I76c6762c515d0c9de1d777c0868b20af;
wire [fgallag_WDTH-1:0]         I6804a691f5de298ab553ee66c3e9610c;
reg  [fgallag_WDTH-1:0]         Id90588b5f82cd32e801fbea04d24e4a5;
wire [fgallag_WDTH-1:0]         If5da296bcf91d370f8341fc402eed6df;
wire [fgallag_WDTH-1:0]         I973825f628679f8bbaf0650136e7259b;
reg  [fgallag_WDTH-1:0]         Ib642d757fae818cd6d713ffb6ce18fc1;
wire [fgallag_WDTH-1:0]         I64673b4b013682f9ce54925853c06ca4;
wire [fgallag_WDTH-1:0]         Ibfa3babbd7909dfada58a7f579281b8c;
reg  [fgallag_WDTH-1:0]         Id76bff2a12cf792e52ccc463647334c0;
wire [fgallag_WDTH-1:0]         Iabfccf7b60f9be4e3714ad753cd8922a;
wire [fgallag_WDTH-1:0]         I0aa6569579526ac14e0d55caa4cef2a7;
reg  [fgallag_WDTH-1:0]         I92ffa890ed6d83d4fc543504e4d421c1;
wire [fgallag_WDTH-1:0]         I73ab1f85232818929b1b2e9d343584a3;
wire [fgallag_WDTH-1:0]         I87c99b1e08ca19dea7ffbfa15ecc2db9;
reg  [fgallag_WDTH-1:0]         Ifc4a65edeaf630b3d29437bcd6c20121;
wire [fgallag_WDTH-1:0]         I06f989f65e614903ffba3594e8112235;
wire [fgallag_WDTH-1:0]         I40ba1533f32b981c4e937b2e48f38ea0;
reg  [fgallag_WDTH-1:0]         Id57a11f56fc223501a9b68b8b05ebd3e;
wire [fgallag_WDTH-1:0]         I0391247480cb6bd6bda2c59dcf8f7607;
wire [fgallag_WDTH-1:0]         I83483243e11dd867b1eea10b6ef0dbd2;
reg  [fgallag_WDTH-1:0]         I522ba8bfc1949337e8befe82cc1e86e6;
wire [fgallag_WDTH-1:0]         Iee114a92d2238e4b8fcdfa79c4c99d6a;
wire [fgallag_WDTH-1:0]         I8265d9994495dbe871b565be6710b428;
reg  [fgallag_WDTH-1:0]         I7153e27c44ebbc2f04e9ba03cf09b5e1;
wire [fgallag_WDTH-1:0]         Ida429b8e252b80b45435af1c6522f783;
wire [fgallag_WDTH-1:0]         I3d4ee0ad8461c2ac5128adc9c231f465;
reg  [fgallag_WDTH-1:0]         Id15e4b4f186ec863f12a54acd8ef8963;
wire [fgallag_WDTH-1:0]         Id3849d43e39d78fd2428109bf9677e0d;
wire [fgallag_WDTH-1:0]         Ib609900664dc10ef97873cccb161c320;
reg  [fgallag_WDTH-1:0]         I95c77eec7575cd7aa93a36f31ea635a2;
wire [fgallag_WDTH-1:0]         I5e51799e585f3dbef5e64908bcfc3e7a;
wire [fgallag_WDTH-1:0]         If8b44d90a4ef1715e9144255d606a27e;
reg  [fgallag_WDTH-1:0]         I3c8114dbe0658cc2889c787f1366abfa;
wire [fgallag_WDTH-1:0]         I6d12e4545b8befb8d09545ea00c8ea96;
wire [fgallag_WDTH-1:0]         I06715db3159c94a5913c05e9827cddd1;
reg  [fgallag_WDTH-1:0]         Ieacf971e9e10fb73c7df9f1da8372f30;
wire [fgallag_WDTH-1:0]         I98d04e6bae91796784a864c5bed637cb;
wire [fgallag_WDTH-1:0]         Ia295ba836438cd4e7c1b03b4261949ed;
reg  [fgallag_WDTH-1:0]         I35de1b03ea865f2c6381ce73e03dc220;
wire [fgallag_WDTH-1:0]         I83b3247bed67d1e2ed488d5b7812851d;
wire [fgallag_WDTH-1:0]         I5f9c502cdffe77bb7e298a9bfdd325b1;
reg  [fgallag_WDTH-1:0]         Idec12e02904ea98c7580919584f2dba1;
wire [fgallag_WDTH-1:0]         I868021f44830a9d81c4ba3dad804f889;
wire [fgallag_WDTH-1:0]         I3f13e4887f4982583fe615807c42d121;
reg  [fgallag_WDTH-1:0]         Ia370c83631a2c1bbf39c7264deafafb5;
wire [fgallag_WDTH-1:0]         I685e59e3865058f29978a8cc2f1b6c7c;
wire [fgallag_WDTH-1:0]         Ie1a491c10dad8dfd4b0fe42977d625b6;
reg  [fgallag_WDTH-1:0]         I05b4a07dfc0d2695eae34bea4c1c6565;
wire [fgallag_WDTH-1:0]         I5a76dd9f4a2078dee81102a9f205ca53;
wire [fgallag_WDTH-1:0]         Id2334d193c70ad43e5b7cdcd923e364a;
reg  [fgallag_WDTH-1:0]         If1ecdc27e3419dd1434e403f237c2b58;
wire [fgallag_WDTH-1:0]         Ice3bd7a4bbf0705a3dc1f89c5ceca084;
wire [fgallag_WDTH-1:0]         I621999a98b66cc50cf7732668af444e0;
reg  [fgallag_WDTH-1:0]         I039c552777d0fb40bebcdd2d4a3394c2;
wire [fgallag_WDTH-1:0]         I5f741a3213cecdf58440120c2ea78e87;
wire [fgallag_WDTH-1:0]         I8c5fe32c1860a2beb9c14634c62a95aa;
reg  [fgallag_WDTH-1:0]         Iaa52fb63184514b6d754bcc896235150;
wire [fgallag_WDTH-1:0]         Idad89ade7f96091abfea876b3af0d5b4;
wire [fgallag_WDTH-1:0]         I5cc33aeefc2bbf0d777b4b59bcba7ec4;
reg  [fgallag_WDTH-1:0]         Ied9781e625c1fa8741853dd6b8b3a9e7;
wire [fgallag_WDTH-1:0]         Ie0ab4b7c79196195db0971e7c7a85adb;
wire [fgallag_WDTH-1:0]         I5a2f74df4050f2898061471586f3fb63;
reg  [fgallag_WDTH-1:0]         I767272262e9d2e85dba1aa93f578f25c;
wire [fgallag_WDTH-1:0]         I0093585d710940feaa8ebdc5fb000806;
wire [fgallag_WDTH-1:0]         I54c68d66f2692522fdd982a31ff0b3a8;
reg  [fgallag_WDTH-1:0]         Ib3b4cd6d8ab17869a2278552c02635c8;
wire [fgallag_WDTH-1:0]         I76a0b74bb633743ac56cf4a0d52f80c0;
wire [fgallag_WDTH-1:0]         I98b0bc583105e551a5c1c7a8b6de61e1;
reg  [fgallag_WDTH-1:0]         Ie7a5cb2ecb3fce35825785b9bca6b3bd;
wire [fgallag_WDTH-1:0]         I11931fd13219c1ae615d164a8f4130f9;
wire [fgallag_WDTH-1:0]         I3ca304e8b6c5440935c6944b64ddde65;
reg  [fgallag_WDTH-1:0]         Ib9a0f8efd3dad427f247ce90fdfb94a4;
wire [fgallag_WDTH-1:0]         I6de7a344ae1574e551c7c10a1773d880;
wire [fgallag_WDTH-1:0]         I33c7b994472de0942347e9b06ed9f59c;
reg  [fgallag_WDTH-1:0]         I69a221a1bd95a588aa74b9bed0357762;
wire [fgallag_WDTH-1:0]         I4920b0740cb56988ba4fc10b86195cdd;
wire [fgallag_WDTH-1:0]         Id5395616ea942f63477bffe5c17560e3;
reg  [fgallag_WDTH-1:0]         I64f125cf2ca6a6da8a9cdae9e246c24a;
wire [fgallag_WDTH-1:0]         I37d27fda03770ad37a1fbad835c076c3;
wire [fgallag_WDTH-1:0]         If90e3127bcb3ed51a225ce72afb0a793;
reg  [fgallag_WDTH-1:0]         Ifac9dd60dd6c543aa94b39c599f0819a;
wire [fgallag_WDTH-1:0]         Ib868fcb71300c09a49719e0b0459ca06;
wire [fgallag_WDTH-1:0]         Ia6ff80807e320ef75fbdad7c86add89d;
reg  [fgallag_WDTH-1:0]         Icf062382a1e462571569ccee75b0a3ee;
wire [fgallag_WDTH-1:0]         I2c67e89b58d7f998c43c68d857fa2381;
wire [fgallag_WDTH-1:0]         If8a6eb502f55f58090ffd901b27086c2;
reg  [fgallag_WDTH-1:0]         Ieed8b94295bed265961c4f52c3379914;
wire [fgallag_WDTH-1:0]         Idb770d9fc630f77beca27c3182279001;
wire [fgallag_WDTH-1:0]         If10a93a95dd1f3e7117e64ae2915bcd5;
reg  [fgallag_WDTH-1:0]         I165eabcdde76821fdc308ff7a8c6d2ea;
wire [fgallag_WDTH-1:0]         I6ab74c183d97a5df7a336c6c66c66e2e;
wire [fgallag_WDTH-1:0]         Id86eeb13a357d077460584e1941e74a7;
reg  [fgallag_WDTH-1:0]         I8b3542a6d64d6a7ebba4124bc6702f3e;
wire [fgallag_WDTH-1:0]         Ic4fc6d6a69dccb796d208aba87ec002c;
wire [fgallag_WDTH-1:0]         I5d7e70c0e768f5868bf9fa07111036e7;
reg  [fgallag_WDTH-1:0]         I7b68afec199be705d766c169f1ece981;
wire [fgallag_WDTH-1:0]         I450cd05f0109ad62ae4ca7f540ac7505;
wire [fgallag_WDTH-1:0]         I48f780aaedbd67e6342d9e0232635ac8;
reg  [fgallag_WDTH-1:0]         I4b6c8226ef2bc20dbd31d242bdb98b8c;
wire [fgallag_WDTH-1:0]         Ia6f1bdee90a01ee3f3e59eec00689d50;
wire [fgallag_WDTH-1:0]         Ia9a47dd6aa0313a806147f2c4a91df0b;
reg  [fgallag_WDTH-1:0]         Ic3b4a86f22caf5b6103d52b6c9d2a991;
wire [fgallag_WDTH-1:0]         I33193403a8d72dcd02e87ae03b668e09;
wire [fgallag_WDTH-1:0]         Id0a9c8069c91546ee6dcdcca1dbddd61;
reg  [fgallag_WDTH-1:0]         Ia37592b207086f63e2d94e3d7d26c740;
wire [fgallag_WDTH-1:0]         I5208f3202b32a30c4abaca4c617d3b3b;
wire [fgallag_WDTH-1:0]         I3e30cc2747c9a7dd9c4fcd144f640552;
reg  [fgallag_WDTH-1:0]         Id0d786026e3ab0ddbffbc20e4d409857;
wire [fgallag_WDTH-1:0]         Ib607167c806dd831aaed4a42b9cf4349;
wire [fgallag_WDTH-1:0]         Ia4433ae2b484d7bfff269cb336831628;
reg  [fgallag_WDTH-1:0]         I333837f976cfc7f90ab0a6dcd8c1ce79;
wire [fgallag_WDTH-1:0]         I42b87e52c168abb775c1e1e5ddfc1958;
wire [fgallag_WDTH-1:0]         I7aef236fed5567b77c8a3f5c22e3bff3;
reg  [fgallag_WDTH-1:0]         Id115b4708a49dcfd167e79ef6993e371;
wire [fgallag_WDTH-1:0]         Ifc4e50801a1606717efd57bd5ac6f41f;
wire [fgallag_WDTH-1:0]         Iff3859ddd94ff25ba5a08a367baf602b;
reg  [fgallag_WDTH-1:0]         I666da645400344644e848ee6f7592d3c;
wire [fgallag_WDTH-1:0]         I5e7282e9a35cead2f4d1d9860d45852c;
wire [fgallag_WDTH-1:0]         I4c0c110a6f362969bce6db69cb1c0bfc;
reg  [fgallag_WDTH-1:0]         Ibafeadd691eee03f855ed657c01022c9;
wire [fgallag_WDTH-1:0]         I8503b90594f3d4b492cca9cf154fc3d3;
wire [fgallag_WDTH-1:0]         I51225282195bed9916ae55ae7887c1d2;
reg  [fgallag_WDTH-1:0]         I10ec5c43a3fb65273053063001307280;
wire [fgallag_WDTH-1:0]         I95010cdf08c373916ab02e3794afa77a;
wire [fgallag_WDTH-1:0]         I58380b8eb6332c81366215b1dd60cea5;
reg  [fgallag_WDTH-1:0]         I05c778eb3588bdaccf714ba456f534c2;
wire [fgallag_WDTH-1:0]         I832fdc71e665ad2acac2576188e0d65b;
wire [fgallag_WDTH-1:0]         I55df86c0751564116c4f1a65de2ac9fa;
reg  [fgallag_WDTH-1:0]         Icd11e8d97a6ac6c0a73e8adee1f98c4e;
wire [fgallag_WDTH-1:0]         Ic21a6f1abcecf14acaf2aa23b7dcdb6b;
wire [fgallag_WDTH-1:0]         I0bc0390d7c9b369ebc92e9547b87b9df;
reg  [fgallag_WDTH-1:0]         If07c2223d4262e22cca9b77c3ed5ee01;
wire [fgallag_WDTH-1:0]         I49847c8c979d9ed82be80f62552e97bf;
wire [fgallag_WDTH-1:0]         Icfe3de1a8dc46c883a65345392921c50;
reg  [fgallag_WDTH-1:0]         If0c8ce0ff66fe2806448f1c819d58ec8;
wire [fgallag_WDTH-1:0]         I7a2bfe5efbe1d0dc222bff675c621485;
wire [fgallag_WDTH-1:0]         I4c0e5a2ba1c2b42970f41699d5ddcb9a;
reg  [fgallag_WDTH-1:0]         Iccdc2371dfd9fda3e506adc2b1681ba3;
wire [fgallag_WDTH-1:0]         Ie0d874ce4b0713de7d087396a1879c54;
wire [fgallag_WDTH-1:0]         Ib81161d68b741b2656196d7284209d58;
reg  [fgallag_WDTH-1:0]         I26e61dca9d045c4661b97afe346152c8;
wire [fgallag_WDTH-1:0]         Iaf4c12394552f42e476b70f6c75003d7;
wire [fgallag_WDTH-1:0]         Ib98bf53c446dcc7920b842d29191fe0a;
reg  [fgallag_WDTH-1:0]         Id488d650b86f5def0668f4a1ef841b6a;
wire [fgallag_WDTH-1:0]         I64d7f4a0df87ce07ce49350610122f79;
wire [fgallag_WDTH-1:0]         I31c34cf26a3890305171a6beca791fa3;
reg  [fgallag_WDTH-1:0]         I479365266255d2228ecd86c350e8d38b;
wire [fgallag_WDTH-1:0]         If51795ea140bec96fdefbc52291801b5;
wire [fgallag_WDTH-1:0]         Idc436d6b98d48c479d762c31bb55e071;
reg  [fgallag_WDTH-1:0]         I08d9c488fd85db45344e649699196263;
wire [fgallag_WDTH-1:0]         Ib0a0f80cb818018b2fe0fd4597325bb4;
wire [fgallag_WDTH-1:0]         I49300b5a8d4f2ce3ef7238f75a2800a9;
reg  [fgallag_WDTH-1:0]         Icde86d0ead44385b07e9a29057417417;
wire [fgallag_WDTH-1:0]         If01a65e097f026a816133c34d73ccff1;
wire [fgallag_WDTH-1:0]         I4c1b051c518c4fa2e042e11cae60de02;
reg  [fgallag_WDTH-1:0]         I21feecd24d912ef3d0aec0e375958f3f;
wire [fgallag_WDTH-1:0]         Ida9ed61c543afde2257053443d133119;
wire [fgallag_WDTH-1:0]         I3ccb0a4c235cd79c6c11271aa1aeb8af;
reg  [fgallag_WDTH-1:0]         I59f419b3bc183a5fe743be3878fac587;
wire [fgallag_WDTH-1:0]         I983a5656d68192a7a3d5a78f17f12ff0;
wire [fgallag_WDTH-1:0]         I8a2e9aba30b284e87bdbb6e91a30d9a6;
reg  [fgallag_WDTH-1:0]         Ib0804d8bdda49ecd0024300eed52be53;
wire [fgallag_WDTH-1:0]         I315445ad2d762b66f94a75d76fbfb839;
wire [fgallag_WDTH-1:0]         I29d269323cfbc900f3868dde96e8da48;
reg  [fgallag_WDTH-1:0]         I37b0efdee34647a5111d698a5a80f367;
wire [fgallag_WDTH-1:0]         I7a97a8fe65e56b0a80c242e13e70db09;
wire [fgallag_WDTH-1:0]         I39a53ef95ccd9c8b1b85e3214af441f3;
reg  [fgallag_WDTH-1:0]         Id382a04e94d0749d0858041bdc5861be;
wire [fgallag_WDTH-1:0]         I2243095f420e4d996f1c69c965932778;
wire [fgallag_WDTH-1:0]         Id64ff7aeff6f73342f863be760a32a16;
reg  [fgallag_WDTH-1:0]         I368be992a21201268c41506396dcdcf6;
wire [fgallag_WDTH-1:0]         I0154a19f9adb43089080304978256c09;
wire [fgallag_WDTH-1:0]         I083900fbd062835b505165f1da19e228;
reg  [fgallag_WDTH-1:0]         I603a008893b5196d9f273b47a9d63144;
wire [fgallag_WDTH-1:0]         Ib8bdc3b41b3cc7132c43833802115880;
wire [fgallag_WDTH-1:0]         I7cf9dee91f849e28b2b2b38d2df00dfd;
reg  [fgallag_WDTH-1:0]         Ie70d3a768bc09ddff6ac68aaba7d9f2c;
wire [fgallag_WDTH-1:0]         I167586906b601ffc473a5b856b213f2b;
wire [fgallag_WDTH-1:0]         If54b33370dcdf69c464c92dab1248828;
reg  [fgallag_WDTH-1:0]         Ifb8bd837ada3d8ed5116db29da82d2a9;
wire [fgallag_WDTH-1:0]         I094a6ac91aacfdd2f8de8a0d776f732b;
wire [fgallag_WDTH-1:0]         I79c5230097571dcdf6ec2a15d633cdba;
reg  [fgallag_WDTH-1:0]         I978b93d46e20cb3eda70e5a976d62348;
wire [fgallag_WDTH-1:0]         I9d4437c250c28653bbccdea6af8b6280;
wire [fgallag_WDTH-1:0]         I71efb4b4bb9b37a4e9b717282c5fbb03;
reg  [fgallag_WDTH-1:0]         Ib404040d4fb58f47f245184c3be01789;
wire [fgallag_WDTH-1:0]         I4afab82ea1a6ad0a36fea0692de1d106;
wire [fgallag_WDTH-1:0]         I0cc336baadd473b40a866cb2944eb719;
reg  [fgallag_WDTH-1:0]         I9c664265c53ebffaad097b70ff3cbbce;
wire [fgallag_WDTH-1:0]         I864d41b77a51fda97ea7017ed18b5fea;
wire [fgallag_WDTH-1:0]         I42d8c11aefc92acf389d12e26217e867;
reg  [fgallag_WDTH-1:0]         I781306c6b1ce0741d9c2fa06865f7a19;
wire [fgallag_WDTH-1:0]         I758ee12b430cda151b452699eb2039dc;
wire [fgallag_WDTH-1:0]         I40412ee4da7bae7c7745064488928be1;
reg  [fgallag_WDTH-1:0]         I16fa2e3dc0b3eddbc72811b51d6ac8ed;
wire [fgallag_WDTH-1:0]         I134cd61326b70030c027a3821d98a994;
wire [fgallag_WDTH-1:0]         I7f6fc13ef5b20f9f1646a608b63f6f77;
reg  [fgallag_WDTH-1:0]         Ia6f232495726806d01b702b0e248b2f2;
wire [fgallag_WDTH-1:0]         I99951d295b9065614c103b3e43fa255c;
wire [fgallag_WDTH-1:0]         Iddd6e6676bf1c96936bb1dbecf6fd805;
reg  [fgallag_WDTH-1:0]         I66b3734060600caa45d699508c5083d2;
wire [fgallag_WDTH-1:0]         I31a4e4f3eac271c84b36c84d7de338fd;
wire [fgallag_WDTH-1:0]         Id0a701ba3adbf20de140020b675cc363;
reg  [fgallag_WDTH-1:0]         I85fae6b23d086235a94a0162e2fb5310;
wire [fgallag_WDTH-1:0]         Id36c36d2b2dd9a79f9887c9950b385c3;
wire [fgallag_WDTH-1:0]         I7e8db4d3310c345d7ada4c2fe05cf9b6;
reg  [fgallag_WDTH-1:0]         I8d6443d1be42203cb834345ae7e5aff5;
wire [fgallag_WDTH-1:0]         I59455b0e53bac4fe6b1cbf609cb03da5;
wire [fgallag_WDTH-1:0]         I3fba42f5d091f0b7a5d8b4d099f72284;
reg  [fgallag_WDTH-1:0]         I717332b7f76e9caf9351f1aa69b72a12;
wire [fgallag_WDTH-1:0]         Ifd633f2ea91cb88aaa2a0bf5579ed1e0;
wire [fgallag_WDTH-1:0]         Ia12c6ec292c6e9fdf58fe58a2af18a53;
reg  [fgallag_WDTH-1:0]         Ieebd34db071409288f489129b70ab599;
wire [fgallag_WDTH-1:0]         I87218b174c1db735ac153604b5ff3e15;
wire [fgallag_WDTH-1:0]         I37448ddc452e005ec974628ade793433;
reg  [fgallag_WDTH-1:0]         I917c874137d64a9a495335c8f8ef5374;
wire [fgallag_WDTH-1:0]         I4608c92d52306432c114f31b9ba6dd69;
wire [fgallag_WDTH-1:0]         I4dee5017c9b71edda82d50b867879afd;
reg  [fgallag_WDTH-1:0]         I15fb4fb838d4a614c468f7d49261bda3;
wire [fgallag_WDTH-1:0]         Iba3f6cde40827d82bc32078344b9bd81;
wire [fgallag_WDTH-1:0]         I2115d9af1cbecde8b5e89c70e582de00;
reg  [fgallag_WDTH-1:0]         I2eb093d2a38ba8cf4be47d1d7f54ecc4;
wire [fgallag_WDTH-1:0]         Ib987bde3ee5a0256d0b8b3aa7357cdb2;
wire [fgallag_WDTH-1:0]         I0e2c6c08e1bcd629678ff57f6bf23be5;
reg  [fgallag_WDTH-1:0]         I8f9affdc5cda0fecc35dd15fc5aeb244;
wire [fgallag_WDTH-1:0]         I3c33a2bfaa82172457b15f4f621eefee;
wire [fgallag_WDTH-1:0]         I00a3c15421af76c65865ff21d2598055;
reg  [fgallag_WDTH-1:0]         I615a443d49d1479338d033d2a2cab51f;
wire [fgallag_WDTH-1:0]         I7ce33eb337b6cacaea13f748061e338a;
wire [fgallag_WDTH-1:0]         I9fa21fd04ffc0a7dc281717e599fd443;
reg  [fgallag_WDTH-1:0]         I0635a3270a9653ca0f23c116fd5b2f97;
wire [fgallag_WDTH-1:0]         I7a8c5be75d87552ca717a87d1a832d21;
wire [fgallag_WDTH-1:0]         I66231fd914db4a60705f1d6de751077d;
reg  [fgallag_WDTH-1:0]         I93a7c75ebce8fbf4c613b4d11dc98b72;
wire [fgallag_WDTH-1:0]         Id9c9cebf44647040da33567d815c261f;
wire [fgallag_WDTH-1:0]         I1142cf230d2632a5972a95316f2fa15f;
reg  [fgallag_WDTH-1:0]         I39334aa9d55bcc001ece37ce2a6c329c;
wire [fgallag_WDTH-1:0]         I6c522c28a0dc265facb1f21ebe51c564;
wire [fgallag_WDTH-1:0]         Ibe1b4cc79b063aafddadcfdb5bc4a694;
reg  [fgallag_WDTH-1:0]         I07e328d23da9383a296ecb03679ec74b;
wire [fgallag_WDTH-1:0]         I86c367b0fd4548d5edfb8863f454653e;
wire [fgallag_WDTH-1:0]         I5371e6575d8bdc6f72cb08beca627fec;
reg  [fgallag_WDTH-1:0]         I8a6e1eace6152af5c98c415804cb60fa;
wire [fgallag_WDTH-1:0]         I800271efe85fcbaee8fe733190e90f6d;
wire [fgallag_WDTH-1:0]         I5e78e43fbf13f79a885bb3cee615d926;
reg  [fgallag_WDTH-1:0]         I6ed4d6c350e8691b3a12ab51419cfa65;
wire [fgallag_WDTH-1:0]         Ia5172996abb4a6bc50046d36ec033c7f;
wire [fgallag_WDTH-1:0]         I735298e3ea4442615df21b3699c94a7d;
reg  [fgallag_WDTH-1:0]         Ie2b9ed680dac51ac866cb830ca17ef84;
wire [fgallag_WDTH-1:0]         Ibe20363746d437eef2c85360425739d1;
wire [fgallag_WDTH-1:0]         I1f2f072bb15b57b5437572b156499e12;
reg  [fgallag_WDTH-1:0]         Ie439b520bbb0c8b29a5ecea167acb1c9;
wire [fgallag_WDTH-1:0]         Iee695b22e8a55479dfcbaa68f5c8b6c9;
wire [fgallag_WDTH-1:0]         I0344e18f3a5fe97467ba8e6641562f92;
reg  [fgallag_WDTH-1:0]         I9f8ef3295578acf5b0a42d074a15a70b;
wire [fgallag_WDTH-1:0]         I7cdb0bf6c7195df38d701768e655af70;
wire [fgallag_WDTH-1:0]         I8aedaf42a56212b44d820d704945cb99;
reg  [fgallag_WDTH-1:0]         Ief01b06341d489e36ee344fd52084ccf;
wire [fgallag_WDTH-1:0]         I1057373671fd4cfba6696f8e88a2d740;
wire [fgallag_WDTH-1:0]         If267b8451ce8bfd1c33273a9c5d08233;
reg  [fgallag_WDTH-1:0]         I3b72a085b104e17dca3d8b2824f84e97;
wire [fgallag_WDTH-1:0]         I7dd9da64c1516e6ae1b703defc4cdc55;
wire [fgallag_WDTH-1:0]         Ie90356409910181f0ffbfdbfea6a47b2;
reg  [fgallag_WDTH-1:0]         I5e1f41e23887493db1d723e1e2cbd996;
wire [fgallag_WDTH-1:0]         I58bf5f51208a98b2448e2b4fad3f63ac;
wire [fgallag_WDTH-1:0]         I43a2d55679515c4766a6e7c19c3ba1e0;
reg  [fgallag_WDTH-1:0]         I0e6f4c7bdc39bd22833f3d9fcfa55f1d;
wire [fgallag_WDTH-1:0]         Icb8281c05ea7168d39d6012a1d622e15;
wire [fgallag_WDTH-1:0]         I2b1e17eeb208749a9c320187e98f3c50;
reg  [fgallag_WDTH-1:0]         Ie346802a8898b4b075be289e062b462c;
wire [fgallag_WDTH-1:0]         I5b16ad2952938bc64f6c9f5ff1ab5a0b;
wire [fgallag_WDTH-1:0]         Ib9c8fc92cd361858e4fb1ddc6dcab191;
reg  [fgallag_WDTH-1:0]         I82ea6f21706a97166ef11af548e80392;
wire [fgallag_WDTH-1:0]         I5d5790b480d08bf6c957f26e24467b9a;
wire [fgallag_WDTH-1:0]         I7ef5a40bcc9976da690ae85ee866b2d0;
reg  [fgallag_WDTH-1:0]         I5f38764f6ecc2dcd1fdd5316102f1f82;
wire [fgallag_WDTH-1:0]         Ieb32ca618265eed3419f01907f48527d;
wire [fgallag_WDTH-1:0]         Ia52b8e11416781165d713f38018047d6;
reg  [fgallag_WDTH-1:0]         Id4034bf7a0e92a6c92d0187e00d3df99;
wire [fgallag_WDTH-1:0]         Ief90415b272ce5707ba28a8470132f5e;
wire [fgallag_WDTH-1:0]         Ibb05d1616c4b57cdf6a268fe16bb9ef9;
reg  [fgallag_WDTH-1:0]         I44692fd63388c57268ea9035a7e4c3ef;
wire [fgallag_WDTH-1:0]         I386c79f4301dea9a37c9ce283e8050e4;
wire [fgallag_WDTH-1:0]         I3be04ed5b262f461ad65b860adc6c601;
reg  [fgallag_WDTH-1:0]         I0c2892a34e5236f1366959eadfd83825;
wire [fgallag_WDTH-1:0]         I0d113fab9d7095f8d1693fec58b7c5a6;
wire [fgallag_WDTH-1:0]         I0bcc8dd8d2adfb33dace6c005377ef97;
reg  [fgallag_WDTH-1:0]         Iccef2754044e7066e191bc5e1a3805f1;
wire [fgallag_WDTH-1:0]         I2bbbe9e5d322d9cee76903fa813765ae;
wire [fgallag_WDTH-1:0]         Iad8fd338d5a105b6fe3a3a021f96f317;
reg  [fgallag_WDTH-1:0]         I8ace46f1c56cfb3f4773324e0f8cae58;
wire [fgallag_WDTH-1:0]         If5317506b6ab92c946af745a65b9e86a;
wire [fgallag_WDTH-1:0]         I46f7c02eeea9f5a0058da869a84e57d4;
reg  [fgallag_WDTH-1:0]         I94ec0139bd827ef5dce2c5ee9eb9aded;
wire [fgallag_WDTH-1:0]         Ib61ddb3ef6c7239bfc720b1761cc0221;
wire [fgallag_WDTH-1:0]         Ie8e3dd32f3ccf581400d8dd0fd5daea7;
reg  [fgallag_WDTH-1:0]         Ied62b116607c549ff5918d5b95e2118f;
wire [fgallag_WDTH-1:0]         I70d669976b271b2319d60114c468cae5;
wire [fgallag_WDTH-1:0]         Ic23bbefb8e8e80ac5df4ef8a50aa5c83;
reg  [fgallag_WDTH-1:0]         I9efa5796297bc922bc5fe17f8319a515;
wire [fgallag_WDTH-1:0]         I96cb81892e2d1737d6cb25522ea2d9e4;
wire [fgallag_WDTH-1:0]         I7c56e54d472bc2301521ecb93aed0ea2;
reg  [fgallag_WDTH-1:0]         Ifa6908d8fda29713d7c1bbaa69b72b53;
wire [fgallag_WDTH-1:0]         I6c87926b040d4006c2294c516a3c46fd;
wire [fgallag_WDTH-1:0]         I4979d09a4bf88992a280e598841f5e50;
reg  [fgallag_WDTH-1:0]         Ieb46857229186ce0391cddb2d30f434e;
wire [fgallag_WDTH-1:0]         I549670efc854cdc29bad1d9bc03e9f5e;
wire [fgallag_WDTH-1:0]         I15264bbbe49fff9c53b8066414264010;
reg  [fgallag_WDTH-1:0]         I67fa03f808026b38ca5b4e71e21588bf;
wire [fgallag_WDTH-1:0]         If54c0c169048bb3e8a1423a58aed0e70;
wire [fgallag_WDTH-1:0]         I32293d41086053c7055fa40ce224631e;
reg  [fgallag_WDTH-1:0]         I70938dfe09b0da9d87dafed6af3fa05c;
wire [fgallag_WDTH-1:0]         I5c956f39031611db595fbc34e6edad65;
wire [fgallag_WDTH-1:0]         I4bd0008f9e9598e9f60a0aa8c2aa2da5;
reg  [fgallag_WDTH-1:0]         Iff30a4e14b6282e9ef92e7f58230b516;
wire [fgallag_WDTH-1:0]         I86851725f5d424c4636f9f41e5a7c7e9;
wire [fgallag_WDTH-1:0]         I584861d31ee7ff0efc61b192c64bca32;
reg  [fgallag_WDTH-1:0]         I43e0faf8070869ab0528a7a4a5cdc103;
wire [fgallag_WDTH-1:0]         Ibec300322cef05615c818b163f8a1fef;
wire [fgallag_WDTH-1:0]         I64f092a873fee78a333072d8c5bbddf8;
reg  [fgallag_WDTH-1:0]         Ib2f0333fac7701ae4a5589d54005b8f3;
wire [fgallag_WDTH-1:0]         I09cc443ecf3811a8a672c4aec1f7d6d4;
wire [fgallag_WDTH-1:0]         Idd6f95a4386cbea3c1533683854a4c75;
reg  [fgallag_WDTH-1:0]         Ie4e1491da700923e81b2c1a246e528b1;
wire [fgallag_WDTH-1:0]         Iaaf5b9288b4eb557d56908bf072cc642;
wire [fgallag_WDTH-1:0]         I32710d1855b18d6c70f6e23a0a440a69;
reg  [fgallag_WDTH-1:0]         Ie8602467de2ece2013878a6b8d3129a1;
wire [fgallag_WDTH-1:0]         Ib224ff2bea17f6e694b10bc7cfdb898d;
wire [fgallag_WDTH-1:0]         I32cc6023f28c6dee2b4b097f1fe890d6;
reg  [fgallag_WDTH-1:0]         I85c93c62f79b1703cb6928f96737cf27;
wire [fgallag_WDTH-1:0]         Ide7d6472bf33f8dcf5c6397c7d7fb733;
wire [fgallag_WDTH-1:0]         Id91b5daa1685f0e3d492f0c3c8306f8e;
reg  [fgallag_WDTH-1:0]         I3dc816ee6c2a818b32f6d4e1228704bf;
wire [fgallag_WDTH-1:0]         Ie6193636ea1cba8b71e1d0d5f2e3c1b2;
wire [fgallag_WDTH-1:0]         Icfdd224aa430648d4afe7b224340b91d;
reg  [fgallag_WDTH-1:0]         Id34d83701e815c01359bc5cd1b9c993c;
wire [fgallag_WDTH-1:0]         Id631b0a4de889a3c3eff4df79367d3d4;
wire [fgallag_WDTH-1:0]         Icbcaa7780b1ad02e07cbbc871b0c2729;
reg  [fgallag_WDTH-1:0]         I0a20e3e26261ba558d681346649cf0b3;
wire [fgallag_WDTH-1:0]         I93d80b8bfb77e7af4d9ac734f26c4e62;
wire [fgallag_WDTH-1:0]         I587b0b57b4f95e8533842965674d1416;
reg  [fgallag_WDTH-1:0]         I331c6e8dbe2ea1e2232f82766926d0e6;
wire [fgallag_WDTH-1:0]         I7fba5fee37c5912e7f635feb8c111b3a;
wire [fgallag_WDTH-1:0]         I1188961bb659f61f0749a27f4ee5c62d;
reg  [fgallag_WDTH-1:0]         Ie27046fd2751357e4a81dc62086f00be;
wire [fgallag_WDTH-1:0]         I22c14ad43399d8a1aee258826a71f50e;
wire [fgallag_WDTH-1:0]         I4ed124c919ba9e29d61a5f771b554ead;
reg  [fgallag_WDTH-1:0]         I0897ceba8201bc14a49ab30318183875;
wire [fgallag_WDTH-1:0]         I3bdc4806c5c09de9a7de8d3601c57bfe;
wire [fgallag_WDTH-1:0]         I735b52f16a8beb195d3e7332f39a1c86;
reg  [fgallag_WDTH-1:0]         Ie7b15aa8ce2492bfb433894efeb967f3;
wire [fgallag_WDTH-1:0]         Id451569510e0d1bbba9002c2b27bb3d4;
wire [fgallag_WDTH-1:0]         I626977a5bbbdb2da503472e8fe6c9569;
reg  [fgallag_WDTH-1:0]         I255add08e982f701508a98db221e617d;
wire [fgallag_WDTH-1:0]         I16753a377bced0688797a464157d847b;
wire [fgallag_WDTH-1:0]         I8f2450ac5c97afe557d068ee5760b527;
reg  [fgallag_WDTH-1:0]         If7ca4919fa1449f38777f742ee1fb875;
wire [fgallag_WDTH-1:0]         I76fd17f22401b66bfc0a6239a0518157;
wire [fgallag_WDTH-1:0]         I13834193a9eb2706cdc680b303efbcf4;
reg  [fgallag_WDTH-1:0]         I24cafcb5b9825321c54e84827a662fdc;
wire [fgallag_WDTH-1:0]         Ie56f8b245ab7833b6939cfea43a99874;
wire [fgallag_WDTH-1:0]         I798a185688b52e59c92b42161b3da7e7;
reg  [fgallag_WDTH-1:0]         I3ede71cb7cb39774aedb9889240a2462;
wire [fgallag_WDTH-1:0]         I668f8103700f044c7764f2281a5b457e;
wire [fgallag_WDTH-1:0]         Ib695cf55b921ed43db22362a28761714;
reg  [fgallag_WDTH-1:0]         I24da9598a6840d3ba7b12fe4f638219b;
wire [fgallag_WDTH-1:0]         Ib75c0ca4f8b59afc2fdd7793bff7ad16;
wire [fgallag_WDTH-1:0]         I1dd0afb6f1a979176d01ab7d37f39bed;
reg  [fgallag_WDTH-1:0]         I0358ca8833007cec4ce5047db32ab7a3;
wire [fgallag_WDTH-1:0]         I3d39fa04d24aa69d19a2db8da00eb0d3;
wire [fgallag_WDTH-1:0]         I559878eee7f3bee345a0f0e891dd2c05;
reg  [fgallag_WDTH-1:0]         I85b5354463c1c15f91ed67292da912c1;
wire [fgallag_WDTH-1:0]         I284b4ccbcb23293efe64fa45b2e0ad98;
wire [fgallag_WDTH-1:0]         I6c688b7c6f01ae353117029f80487ec4;
reg  [fgallag_WDTH-1:0]         Ie93731739ace44811198d0fd95b04a6a;
wire [fgallag_WDTH-1:0]         I689ac029a268fe244a8793367c900602;
wire [fgallag_WDTH-1:0]         I62ad8f36d1e0b80d0d04a326d80e1729;
reg  [fgallag_WDTH-1:0]         I464926faf4e005ad491b0bf93a365e07;
wire [fgallag_WDTH-1:0]         If53dace3e8a7be2524d711de84855015;
wire [fgallag_WDTH-1:0]         Icf1eb32cfc4a48f7e53c180aa94f5833;
reg  [fgallag_WDTH-1:0]         Icdaaccfead6f2d5ac2ce19caf1104d57;
wire [fgallag_WDTH-1:0]         Ie3fe635b63e13732c17ae2076b807b4d;
wire [fgallag_WDTH-1:0]         I8bdfadcfa5cb308e6e254d42997340fd;
reg  [fgallag_WDTH-1:0]         I916d6f9429f2b0cc1bd6fb900484cde5;
wire [fgallag_WDTH-1:0]         I1e196a61113d4db7b51f3d6b18c33da3;
wire [fgallag_WDTH-1:0]         I6ceae370fa59e601566286b127dec684;
reg  [fgallag_WDTH-1:0]         I0142f9b3d361a0d88522f1c5f54aca84;
wire [fgallag_WDTH-1:0]         Ic80e494400a5d7dcfdbf96424391e596;
wire [fgallag_WDTH-1:0]         Ifcf5bef8ae2998f0bd3d270e98acc1c5;
reg  [fgallag_WDTH-1:0]         Ie6871983b4f81b5321519647e628bd0e;
wire [fgallag_WDTH-1:0]         I69d20a7aaf2c66ed9b41fdeff0d5c6ec;
wire [fgallag_WDTH-1:0]         Ic1c8e5992501f0e04191fe6dadd2d56c;
reg  [fgallag_WDTH-1:0]         I17d7be125df22153fc1ed051d4e0770a;
wire [fgallag_WDTH-1:0]         I19b667bdb053ebd555aaa540d3a76f95;
wire [fgallag_WDTH-1:0]         I3f88a35a94c77ca32f3b58c4b509b21c;
reg  [fgallag_WDTH-1:0]         I50b13959e06243e54fad2088eaf65aa7;
wire [fgallag_WDTH-1:0]         Ifc3d9cc420aa1274fed24b38c4d9fd8a;
wire [fgallag_WDTH-1:0]         Ib875be40a1b73b1583cfc9cfec760e31;
reg  [fgallag_WDTH-1:0]         I7a423d609b492f73d5a322849b4b1cce;
wire [fgallag_WDTH-1:0]         Ie8a6ed15370edd38bfc92290bf7bb55a;
wire [fgallag_WDTH-1:0]         I15eae5f35300569305dc03e24d1cdd7f;
reg  [fgallag_WDTH-1:0]         Iefec67e214d1868670a34a7297d4a1c8;
wire [fgallag_WDTH-1:0]         Ife5a1b49d4b0342f06ef83750ab914d4;
wire [fgallag_WDTH-1:0]         Idffbcb47f4a04fc71d1406e46f4ab6c4;
reg  [fgallag_WDTH-1:0]         Iae7da7fdc002b635ce4285d6916d8156;
wire [fgallag_WDTH-1:0]         I9906c49536062867b98ed290e49bbe50;
wire [fgallag_WDTH-1:0]         Ifaf09d72a75fd4f9948e997b8a8388f4;
reg  [fgallag_WDTH-1:0]         Ic561e44b2caeae84df6720f1afa3e8f6;
wire [fgallag_WDTH-1:0]         I41be66295070bec696e91d0f9efdc233;
wire [fgallag_WDTH-1:0]         I661c1624e4d13ba49efc3fb608ba84ed;
reg  [fgallag_WDTH-1:0]         I5be062f5b52e104ca67e615ce75a7c80;
wire [fgallag_WDTH-1:0]         I4838b956d8a597e78bef9a0fce82542e;
wire [fgallag_WDTH-1:0]         Iaa8bf572a01757f5e9321e6ff7364d7e;
reg  [fgallag_WDTH-1:0]         Iecdde23e34c34ee0055be41f44959a19;
wire [fgallag_WDTH-1:0]         Ia06cb40e9a3341f34625c5804e02c07f;
wire [fgallag_WDTH-1:0]         I7ef389b5ce4bdcca7fab9e9ec2bfa3a9;
reg  [fgallag_WDTH-1:0]         Ibe09be9cad0e56d5403868d072d7d628;
wire [fgallag_WDTH-1:0]         I4eaad70758412eab097822b2feda7a57;
wire [fgallag_WDTH-1:0]         I4e7823ff42f8f44a21778dc4b3633a67;
reg  [fgallag_WDTH-1:0]         I464e1f3c13acaf466afb354a9b35ba0a;
wire [fgallag_WDTH-1:0]         If89e1da3daa6fd3090781723173b140b;
wire [fgallag_WDTH-1:0]         Icf5823b64f3a9b7d2656656b61724bcd;
reg  [fgallag_WDTH-1:0]         I160a465c22073a53510e8a4c489c3321;
wire [fgallag_WDTH-1:0]         I9ac67c519fd5a55d0ffb727389781492;
wire [fgallag_WDTH-1:0]         If77f93c61b38d10360f7dd382686d91c;
reg  [fgallag_WDTH-1:0]         I9e86d3e49827861b24f4fbeb308ad3a4;
wire [fgallag_WDTH-1:0]         I73799799e5469ae887dec9b46c9c965d;
wire [fgallag_WDTH-1:0]         Iede699ff40abf5838b54678df24ff29d;
reg  [fgallag_WDTH-1:0]         Ib96b7d796e20967e89a47e01bf424e59;
wire [fgallag_WDTH-1:0]         I7ebd7c3f0617cf500deeb8c152c09af2;
wire [fgallag_WDTH-1:0]         Ia1c9e86b6112a18e7aa613315343e696;
reg  [fgallag_WDTH-1:0]         I565e666f6ba14b4c25e0dd402a3266e1;
wire [fgallag_WDTH-1:0]         I2ee7d4f522ba17ca941c67079309c398;
wire [fgallag_WDTH-1:0]         Iad94272a2a302f4b6b963e71ccd64ccb;
reg  [fgallag_WDTH-1:0]         I97e8bac5becd5128bc70f3bb48f73e6c;
wire [fgallag_WDTH-1:0]         I62d13683ba05cfc27d9ae9a82fb04689;
wire [fgallag_WDTH-1:0]         If4d54d2b483d85b0c4f31db721b14323;
reg  [fgallag_WDTH-1:0]         Iced39475c6e5e3d8f36d2a5c5a80f146;
wire [fgallag_WDTH-1:0]         Ic06032eaed49f01d3d5513b2d145eaaf;
wire [fgallag_WDTH-1:0]         Ia3b12887d984da936d88d657090f8972;
reg  [fgallag_WDTH-1:0]         Idcbd423c2b963c1f693dea2ddf428195;
wire [fgallag_WDTH-1:0]         Idba6350812d3c90bee79636db48257e2;
wire [fgallag_WDTH-1:0]         Ib23dbfa64e4a9364e0c1dbbc6b2ff001;
reg  [fgallag_WDTH-1:0]         If1640e294bdcc51ee12fca5b3a33be6d;
wire [fgallag_WDTH-1:0]         I6e7ed391604c7e0ff7cca99d5aeddc9f;
wire [fgallag_WDTH-1:0]         Ic8d47dcabda3b23d4451e609395c4698;
reg  [fgallag_WDTH-1:0]         I4754c6c355e632d2ed1336b5a88c3b46;
wire [fgallag_WDTH-1:0]         Ib78d45cc282f110ed3ddaeb706a0fc12;
wire [fgallag_WDTH-1:0]         I5d4903ecdf83967c7f60d876bcd0b215;
reg  [fgallag_WDTH-1:0]         I1634d703ad5d6e58a97b13ef957bdbec;
wire [fgallag_WDTH-1:0]         I0f5d081f9846ad888eac13d4916f5b8c;
wire [fgallag_WDTH-1:0]         Ief11c4434035425db82902c38e47be48;
reg  [fgallag_WDTH-1:0]         I804e1e6a01edeb780b0159ecae707b71;
wire [fgallag_WDTH-1:0]         I607bdd63c3ee70e2721de3f994d2923e;
wire [fgallag_WDTH-1:0]         I1c3a6173bb59263a31998a5a69aaa38c;
reg  [fgallag_WDTH-1:0]         Iea3c0f3c3c3017fe87a3b01647189fe0;
wire [fgallag_WDTH-1:0]         I5453775d628c6c01c088278b6e090ddf;
wire [fgallag_WDTH-1:0]         I2d77f481539c1258b61c2a6ca7208455;
reg  [fgallag_WDTH-1:0]         I756b7d7e6bd3e71afa472e7e4727264a;
wire [fgallag_WDTH-1:0]         Iff51257cd95c2f3a38c64ae872317410;
wire [fgallag_WDTH-1:0]         Ie88dbc3340cd953d819e7fa12d1fe3fb;
reg  [fgallag_WDTH-1:0]         Ifbeae0a2acf80eda6ffd050d3bb07eb3;
wire [fgallag_WDTH-1:0]         Ie5faf4f522c8d24bc2d3725be57453e3;
wire [fgallag_WDTH-1:0]         Icad54aaa6f380f2808749db56b76a959;
reg  [fgallag_WDTH-1:0]         I990ab4dcb70ee860c2c40f306ef314d3;
wire [fgallag_WDTH-1:0]         I7952b4b62af35c930dcffe35b1629100;
wire [fgallag_WDTH-1:0]         If41dd08de4b2e28dae0404832fa0edd4;
reg  [fgallag_WDTH-1:0]         Ib131087ea9ccc4bd161c3f9ac2c72303;
wire [fgallag_WDTH-1:0]         I47337a0b371f749c3f7f5118362c2301;
wire [fgallag_WDTH-1:0]         I161c799aa59a0d82ca4db2b7b0293fdc;
reg  [fgallag_WDTH-1:0]         I9a967ac9d11583faaa783984229aeb2c;
wire [fgallag_WDTH-1:0]         I21ea597751b3243936aea7c07cc90f70;
wire [fgallag_WDTH-1:0]         I911555064a463cd6a7ebdb4de801b8fb;
reg  [fgallag_WDTH-1:0]         Ib9921dfcf121e5f4ac4d8be83a868210;
wire [fgallag_WDTH-1:0]         Ibdce05e98adef0314000dba3c482ace6;
wire [fgallag_WDTH-1:0]         Ib2fce59707fcc6d804b748678d3fa03a;
reg  [fgallag_WDTH-1:0]         If22d8fd45caed08b2c7cee8b7349700f;
wire [fgallag_WDTH-1:0]         If0dbc84f59311eeabfb57b5fd0c3b632;
wire [fgallag_WDTH-1:0]         I5d40a4f6c096b4962285bee680a366c0;
reg  [fgallag_WDTH-1:0]         Iabf029e67c7f827faf17b6518cd1bfa3;
wire [fgallag_WDTH-1:0]         I74f2e7798a8383b78a5e7b816c2370af;
wire [fgallag_WDTH-1:0]         I692db6abe25b064802b76618cfd8d151;
reg  [fgallag_WDTH-1:0]         Iaeab83001c6285630e3404ae67227f46;
wire [fgallag_WDTH-1:0]         I58ee302a3a1faa2b44d9052bffbc2a03;
wire [fgallag_WDTH-1:0]         I396539ceb8b33c1dfe096f71954586e7;
reg  [fgallag_WDTH-1:0]         I53ac6d02d2bfc9aca9469148753070a7;
wire [fgallag_WDTH-1:0]         I979a71fc0942bf62c06405bb63a717c5;
wire [fgallag_WDTH-1:0]         I4335c153299e851249a1492c14987447;
reg  [fgallag_WDTH-1:0]         I61992979f60b26d313efd1dc23bb54ab;
wire [fgallag_WDTH-1:0]         I30be0ac758b5a0fbacb1c51a36ca8a73;
wire [fgallag_WDTH-1:0]         I5d81087b001624992357f909d2d7e9e2;
reg  [fgallag_WDTH-1:0]         I8b46b3f0835310114208963de7ac8e97;
wire [fgallag_WDTH-1:0]         I9c50e0a8a01aaed98ae54530d5c76ba1;
wire [fgallag_WDTH-1:0]         I2b8539d21de88ded1152a26741003b99;
reg  [fgallag_WDTH-1:0]         Icda26ba6f5c7f77a80776b2c1bbc975d;
wire [fgallag_WDTH-1:0]         I0daac80ebeec26e428328344a398ce57;
wire [fgallag_WDTH-1:0]         Ib5f0b838019cb6c583e7aae384a7ffba;
reg  [fgallag_WDTH-1:0]         I0863565b3ae88137a2384750436f9e19;
wire [fgallag_WDTH-1:0]         I6739f13ea431943bb5bacb4a05140063;
wire [fgallag_WDTH-1:0]         Iee7fb9e4ff68c15395c13083bb14e8af;
reg  [fgallag_WDTH-1:0]         Id646110f8d09cd47dc7695e05f73efc6;
wire [fgallag_WDTH-1:0]         Ifa0e560fe6445b006ab74096a807b90f;
wire [fgallag_WDTH-1:0]         I18176a5b74de8d98a21cbbbfd35b0bdd;
reg  [fgallag_WDTH-1:0]         I5999eef2304e579a3d47e4f15ba336e1;
wire [fgallag_WDTH-1:0]         I9595c0fd77d6a0610eb859dcd2b67d1d;
wire [fgallag_WDTH-1:0]         I033c58d2361a232bcfa2eda4ac665761;
reg  [fgallag_WDTH-1:0]         Idd302bdc6ff8368a6b73d53bbc8f8425;
wire [fgallag_WDTH-1:0]         I6f3e685e70fa700b52bec62d0aed942c;
wire [fgallag_WDTH-1:0]         I0ddecbd9a2e867e3bf8a447434f626a1;



reg                              I92cb615e2c439914e72ce001256518e4;
wire [MAX_SUM_WDTH_L-1:0]        Iea07d1adf9016a29cffd61d183e268d0;
reg                              Iad799775eb657f8973e6dfcf70a9875c;
wire [MAX_SUM_WDTH_L-1:0]        If92db65b39a83e1c699e4cc6d7f9e57b;
reg                              Ifb064c69c7110c014593149ae69c75fb;
wire [MAX_SUM_WDTH_L-1:0]        I8f2986bc015fcc64ac5e5395ac6dd851;
reg                              I7f7b30f2acbb8e31f50b58096b738254;
wire [MAX_SUM_WDTH_L-1:0]        I355725a804e0df68b4acf96ca98f2448;
reg                              Iefe4099ff7e457f6b9fefc83e176c1a0;
wire [MAX_SUM_WDTH_L-1:0]        I78212ae965ab2dcb2eed0b060d6b253f;
reg                              Icddb43f9b760a4597a0bb637fb405616;
wire [MAX_SUM_WDTH_L-1:0]        I0b56aa7a1b7549c91dddd3a06ecbaacf;
reg                              Ic76e72b434b47c10ebac3fac4ea50bde;
wire [MAX_SUM_WDTH_L-1:0]        I71412803cc5229025487255aec62ec4f;
reg                              I9eb87e62d23bc87d7cd82c0f329f247f;
wire [MAX_SUM_WDTH_L-1:0]        I32fcb28a27356bc6f403528836ea4c1f;
reg                              I2eac5b39c6f485c9ae0bd341f894633d;
wire [MAX_SUM_WDTH_L-1:0]        Iad354d876cb9fc72fc0143e6f7da9357;
reg                              I76992221b1edff5684c482df7ac4693d;
wire [MAX_SUM_WDTH_L-1:0]        If6e745bb85abba7282dae1f6f701225e;
reg                              Iada5bc4a51dc1bf57bb9cca11326bdff;
wire [MAX_SUM_WDTH_L-1:0]        I93bb43c1b89d4c70a57bdc019d64fd22;
reg                              I364ed3f83c49626bc3b939e53524d9c7;
wire [MAX_SUM_WDTH_L-1:0]        I7a2e554d07bbea291f2cfc18694fca3a;
reg                              Ic2b000c3b2ca3beff2d427caab04701a;
wire [MAX_SUM_WDTH_L-1:0]        I3e59b2419c7dd1553b792d536208514e;
reg                              I8e873fb2321eea82bb590a92411e2e2c;
wire [MAX_SUM_WDTH_L-1:0]        I46894c6526983bf1ce4b503159131b41;
reg                              If4cb744ee52b6ae793431cd038069b57;
wire [MAX_SUM_WDTH_L-1:0]        I6404d0df952b5bf8292c753e4c6f35d8;
reg                              I7741e239c16828889d488cc87647c154;
wire [MAX_SUM_WDTH_L-1:0]        I8522c402e654d007abffcb0e904af5e6;
reg                              I7979161aa1e2262ebea862004c387697;
wire [MAX_SUM_WDTH_L-1:0]        I5ed85845c39337c37791f16e718069b4;
reg                              Ic62fc602da3d16fe13d03a49a21269d0;
wire [MAX_SUM_WDTH_L-1:0]        I89013d61c1ea8da8b1c6071cc21c316f;
reg                              I94009bb7239be96243902ab0f0abea7e;
wire [MAX_SUM_WDTH_L-1:0]        I4102100fa5f1dd299af0190862efcc42;
reg                              Iae7b72abf4d3c536330a229e3836b441;
wire [MAX_SUM_WDTH_L-1:0]        I4939f69abb1eac56d5021e06406a93b5;
reg                              Ie5d9cc18b2dd300132470f206452ff17;
wire [MAX_SUM_WDTH_L-1:0]        Iadbd245bf842aebb456417579a3e6296;
reg                              I7c791c854d0bc28e8dd787545f8fbda0;
wire [MAX_SUM_WDTH_L-1:0]        Ifc8ece44a4e68c3117eda9e65f3084d2;
reg                              I5b177dd5c14ad082516b47f550875682;
wire [MAX_SUM_WDTH_L-1:0]        I91679dfab57a372eddc7f9b94a231edb;
reg                              I55e4ad2d71a29ad63b4999d64ac0dc4f;
wire [MAX_SUM_WDTH_L-1:0]        I2213c1a2b831f421707a261f5a58b1b1;
reg                              I59c5da6338f431a626c86a065a355c35;
wire [MAX_SUM_WDTH_L-1:0]        Ic53b875b2ddcba11406eb2ca39354757;
reg                              Ia098bbeda8b755ece6b88eac83d03e55;
wire [MAX_SUM_WDTH_L-1:0]        I634484f00590216c0f74f975c9c83400;
reg                              Ie7470dd75b54d14038de19e4d3043ba9;
wire [MAX_SUM_WDTH_L-1:0]        Ib3b1db2d8b669988c887ed780e439b26;
reg                              Ie95662d4faf6b5a4cd5ecfa41697b983;
wire [MAX_SUM_WDTH_L-1:0]        I735db8b0ee0ec98e4cce0030b11508da;
reg                              Ia1b617e3d141263b51e58c5ef0bd7a89;
wire [MAX_SUM_WDTH_L-1:0]        If1607e907e626902ee26d15020a64c21;
reg                              If9a5d830e3ade0fd96b98f5949f165f0;
wire [MAX_SUM_WDTH_L-1:0]        I081b38dbb37d4c14a6a9fd3fefa13daa;
reg                              Id3de87169c440f95d406693ef77cacd6;
wire [MAX_SUM_WDTH_L-1:0]        Ibac5e7b6d4bf5cd6926358318f0c418f;
reg                              I3751f191f5009322acb7c9be4f8d7129;
wire [MAX_SUM_WDTH_L-1:0]        Iadfc60386481092ae85cc148a2c40abb;
reg                              Ic1927bb3335f6a28c0816eba12d3975e;
wire [MAX_SUM_WDTH_L-1:0]        Ie0ee5445c56a5f9b41640b57422206de;
reg                              Ia659126b51468cfef48c97a135a71500;
wire [MAX_SUM_WDTH_L-1:0]        Ie5f8620371236cb11c9e88c16b509ee8;
reg                              I3c3c22bf63e55a81ae91b1dd1ef615a0;
wire [MAX_SUM_WDTH_L-1:0]        I8d7c1fe2e33bbd45379b0325a3c5e989;
reg                              Ia62832d325f86160285c4d1a790a32cb;
wire [MAX_SUM_WDTH_L-1:0]        I4fbdc4ee57a3be42b62d9bd43078d6ef;
reg                              I83c7d177eec2dad0a924557cdc91ba77;
wire [MAX_SUM_WDTH_L-1:0]        I5510b88bfd65811b3200adf4ef975b48;
reg                              I7050adb9d06f767549b7f35c4679e391;
wire [MAX_SUM_WDTH_L-1:0]        Ib57ef2f577cca54713c16717cbbd1ce9;
reg                              I04aacd95d9e44657f616e01c9053f0fb;
wire [MAX_SUM_WDTH_L-1:0]        I15943aa74e9fbbaebdc0d54eb6a3bffa;
reg                              I2ff317d57f59747c4524ef4278d51092;
wire [MAX_SUM_WDTH_L-1:0]        I6ac24c46319a787daa5c545de8c6eeea;
reg                              I8bd2a9d90074500698b302cb8db7f03a;
wire [MAX_SUM_WDTH_L-1:0]        I52403a0454e5fa002e79eaab7ea497bd;
reg                              I3b8cdfb1440732ce98cd1676e05a2af1;
wire [MAX_SUM_WDTH_L-1:0]        I634f0ce28934600a1a31ab0d8e59b4a9;
reg                              I671de3d408b5b783541663c7f1e3a6fa;
wire [MAX_SUM_WDTH_L-1:0]        I7103aa739616a39c03e675ea0efb0335;
reg                              I446857735e680cae93a24dccb59b1924;
wire [MAX_SUM_WDTH_L-1:0]        I0296d01fd3f9a269a617efd4beea9b8b;
reg                              I77b05a8aa92c66a235195a66dc13c0cc;
wire [MAX_SUM_WDTH_L-1:0]        I065a81ba25962785215583e7ece27661;
reg                              Ie92110d19f4886cdfcfacd0920c06a4e;
wire [MAX_SUM_WDTH_L-1:0]        I631a3300cb6685f47da7781940ec5d27;
reg                              I36ba87b69b5b9dd919319230f697dfad;
wire [MAX_SUM_WDTH_L-1:0]        I8bbe1a2ace8f51aa22cca5d9fc66f136;
reg                              Id20e72ac258d1d1b6cdca1e6c9e3596d;
wire [MAX_SUM_WDTH_L-1:0]        I38c3e3e136acb79c8a0ff850bcc55f16;
reg                              Ifc34f5d6b7a7d0533439794958959856;
wire [MAX_SUM_WDTH_L-1:0]        I35b2c7e9cdc53a98913e1c16a3a47b37;
reg                              I849ee5d34760be03d4285185136aa52e;
wire [MAX_SUM_WDTH_L-1:0]        Ib1a2b31d49ae476e2f1fb9acba2d5af0;
reg                              Ia3559d98eb372b7307f30ad1f7c4c7cd;
wire [MAX_SUM_WDTH_L-1:0]        Ic72f41f9bbf470aee3c9b9b8787b31c3;
reg                              I7332e088bbff69db19c62685e033d26a;
wire [MAX_SUM_WDTH_L-1:0]        I3ea4c33a9419820ed54460eb64134dff;
reg                              I44daa5992b00e7af19adbee70bf01f2b;
wire [MAX_SUM_WDTH_L-1:0]        Ia0d940e16c8cbd4f7544f5a5cd7d83b2;
reg                              Ie517386cb5832e406fefc5e85eb2e7d1;
wire [MAX_SUM_WDTH_L-1:0]        I4a8abfa0896ce414d9b98093ef84455f;
reg                              I9b096ce09467c10f448496fda13987d2;
wire [MAX_SUM_WDTH_L-1:0]        I680be647bf2a62e0ee9b5d379dc87b4f;
reg                              If1c0a3726041f70e508d68cbf6e40e04;
wire [MAX_SUM_WDTH_L-1:0]        If4d75f83299a21802b6fbe136913489f;
reg                              Iaf36ce8598a29573979c683a5e2cf9fd;
wire [MAX_SUM_WDTH_L-1:0]        Ibddfda6413e3dd2f483c3174ea836b6a;
reg                              Ice82cfe55a5f226746e59e5c8beb46be;
wire [MAX_SUM_WDTH_L-1:0]        I33bddb0adcc2af7b12a83bf843036385;
reg                              Iea1297491d1dfe98f395d8c73808a893;
wire [MAX_SUM_WDTH_L-1:0]        I529f92b82248efe2cf64f7da0ec8283c;
reg                              If43dd31198c8a0da6fabd194cf13bb70;
wire [MAX_SUM_WDTH_L-1:0]        I2f34af0036985cd94ade9cc905bec065;
reg                              Ibeb8c72b90b50c6897224ca1a792fa56;
wire [MAX_SUM_WDTH_L-1:0]        Ia1a0d8d7dfd6e877f15cce773f85f5b7;
reg                              I8e87530a131b5a73cad6df68b9e4967f;
wire [MAX_SUM_WDTH_L-1:0]        I5dd29fd1a73df5662d2b636e7285bad9;
reg                              Idf8d15c7bd7705b9aafbda09c3a5b46c;
wire [MAX_SUM_WDTH_L-1:0]        Ide530e6f4622c8a7b101b6dce9650e42;
reg                              I2aea17846a53e2eb2968581ee2c48226;
wire [MAX_SUM_WDTH_L-1:0]        Ibaf00a6780325882067a79f0c4d693d2;
reg                              I169d8f2bb5fde5b202b4239b7a7f1ed5;
wire [MAX_SUM_WDTH_L-1:0]        I16e3559c63ebfed83d6698fc9a9cd93a;
reg                              I40a223380fb4414a3f26a08cb90025ec;
wire [MAX_SUM_WDTH_L-1:0]        I9747a02384abb1c2dd1f52b3a5a999cc;
reg                              Ie117f6ec475f5d6444998af151ce4e69;
wire [MAX_SUM_WDTH_L-1:0]        Iceb7a1d4c23806b8f5824016779ad129;
reg                              If7f3174da35dd39af7f4792aaa649bf1;
wire [MAX_SUM_WDTH_L-1:0]        I40ef50004a60ae58aedc49eb5e6797c9;
reg                              I719a892ad54e63b217c7271741b29cc5;
wire [MAX_SUM_WDTH_L-1:0]        I753f92da60980736440aba814a156f1e;
reg                              I4acf6d84471cd237f65c9b2391b7a20c;
wire [MAX_SUM_WDTH_L-1:0]        I4ac79b67a8904b95f7912d24af420585;
reg                              I7a387a1f887c32e9d0f8e89912a8618c;
wire [MAX_SUM_WDTH_L-1:0]        Iad44c932cfa5c249c5e59f8c706173a8;
reg                              Ib862ac63c230ccde7fae0e62f9d047fe;
wire [MAX_SUM_WDTH_L-1:0]        I10f14b6433498e3b9e9bf021b60115e8;
reg                              I8f1a8a22637d37c3692e808d5eb3d543;
wire [MAX_SUM_WDTH_L-1:0]        I96008f47b9f134c9c4274cfcfb28e550;
reg                              I6f420c64640dfb0c001f57df7e3b4504;
wire [MAX_SUM_WDTH_L-1:0]        Id0344146d1a53d418add6d2b185377dd;
reg                              I3600031716c2b4e21c9f577d34e033dc;
wire [MAX_SUM_WDTH_L-1:0]        I1eede74f12d37331b399eb7136bc621f;
reg                              I002820a37fa7c6c504c487df4368e2cf;
wire [MAX_SUM_WDTH_L-1:0]        I3e4754acc31d99bc71525789bdee0c1a;
reg                              I8a4c1f23212ff846400651b100add502;
wire [MAX_SUM_WDTH_L-1:0]        I11c1fc94a3bd6dffa17e1571cc6ae97c;
reg                              Ice1ce5b4c30841dd92268559ebadafcf;
wire [MAX_SUM_WDTH_L-1:0]        I5395ee57418c31e11cf847f0f514ec19;
reg                              I3eeeb1949945032d6c1759875426b733;
wire [MAX_SUM_WDTH_L-1:0]        Iff125392fa39afebae1637a19c4e23ec;
reg                              I384d5377ee6b8f7eb2db23a2e444ddbc;
wire [MAX_SUM_WDTH_L-1:0]        Ia6308e16fae5428f4ab6560f5b21479a;
reg                              I30d615203b697787ead37394953925cc;
wire [MAX_SUM_WDTH_L-1:0]        I5ea02b5349cd4d99ccbcb6b26f0cfdd7;
reg                              Ib16548d471f0a4f4625852ea04335dcc;
wire [MAX_SUM_WDTH_L-1:0]        I21de4f6194dec9e3c401934db92c25e7;
reg                              I0987c561670b7b2b6683303c1be39561;
wire [MAX_SUM_WDTH_L-1:0]        I57d0920119f8901bd4dea2d5f8fb5d90;
reg                              I2bdf4736022e5da7294a0e851006a124;
wire [MAX_SUM_WDTH_L-1:0]        I89537301987d6da0dbe6cff3caab3ff4;
reg                              Ic6fd9592d2ffcb8f4ca83c6f0bd19975;
wire [MAX_SUM_WDTH_L-1:0]        Iaf0bbbe791bb71d0f557dc71caa5fb87;
reg                              I14bf11ad80890227e47fda26ae1b9c24;
wire [MAX_SUM_WDTH_L-1:0]        Ic7ff9cde71054c1ee9eef81eabdd7061;
reg                              I8ca17b6cf35e1b1f8f601604575d3f27;
wire [MAX_SUM_WDTH_L-1:0]        I88c10c47ae424fbdcb852fbf1e94127c;
reg                              I275cd09649a750edb8ae8313e4e1e279;
wire [MAX_SUM_WDTH_L-1:0]        Icd2e75e47cab1d539ba9ff1b6e1d7155;
reg                              I7d6a6026eb3c4d06e682523424f9628f;
wire [MAX_SUM_WDTH_L-1:0]        I37e6bc7aff363ed0ed1f84b23c5f3e34;
reg                              Ia0c192e590d8c914555b434ce5a634a8;
wire [MAX_SUM_WDTH_L-1:0]        I733605337bf6972630c089d32fd7f98f;
reg                              Ic98c8641d2022080297c54ff2539e75d;
wire [MAX_SUM_WDTH_L-1:0]        Idcb1d8bbdeaed6768c2a418c3048e6ee;
reg                              I87f34821cd0b58f8855b25c75f2dd32d;
wire [MAX_SUM_WDTH_L-1:0]        Ia89da2f1890524ad3519ab403dd0686c;
reg                              I87211ac14d832ad3205d47fb83cf256a;
wire [MAX_SUM_WDTH_L-1:0]        Ie33a780b0221084898c9fc5b237b244a;
reg                              Ib81431cfb3b281555fa7e5b4582a2524;
wire [MAX_SUM_WDTH_L-1:0]        Iabbd1668e0014df518ede5216232834c;
reg                              I835b902949c2c4c09b757d4d35574a76;
wire [MAX_SUM_WDTH_L-1:0]        Ibd89458312687610aa166a9538968851;
reg                              I8510240df7dc41f85ad58a39868a1fd7;
wire [MAX_SUM_WDTH_L-1:0]        Icbaf92a8e9875bcb19a1d074779a9ea5;
reg                              I1b6abc8fbab3849b285e9f88a4fe867b;
wire [MAX_SUM_WDTH_L-1:0]        I80f3c8559da8e97bc5397bb8b621a0bd;
reg                              Ied638fee34f8baed4154b0b72e43a21e;
wire [MAX_SUM_WDTH_L-1:0]        I7a0eada108891aba06cecab5071232c9;
reg                              I14fa7aebb608d4a3d67176ba27d34d9a;
wire [MAX_SUM_WDTH_L-1:0]        Ie21a2c9b22e7bf8425fb5c0f33e5f4f7;
reg                              Iad90879acba3fc2101829549264960f3;
wire [MAX_SUM_WDTH_L-1:0]        Iaa5b2807e5cc2403c5787eeb3d10ca6b;
reg                              Ife0952b85f14a960007b67646b0cd969;
wire [MAX_SUM_WDTH_L-1:0]        I6da2b3a481ee71b85f3087b36b399288;
reg                              If876ca6a14ffb4323503ed46666bc25f;
wire [MAX_SUM_WDTH_L-1:0]        I11094e852295755925c3c61f1df81643;
reg                              If2dfcbf493b761fb5d7c622e739b23f3;
wire [MAX_SUM_WDTH_L-1:0]        I9c633aa620cca127b0ff8cf882178e76;
reg                              I2c8f4a147b363d9c5ef0e080d9a9ed40;
wire [MAX_SUM_WDTH_L-1:0]        I694d471fd353eb54aae08a2afa7b645a;
reg                              I485f9d1104a965d5d035feef912a2ca8;
wire [MAX_SUM_WDTH_L-1:0]        I816704585ad393f685731104ad3ec64f;
reg                              I10fca5f2cbf5e2bc3433c0dda579a051;
wire [MAX_SUM_WDTH_L-1:0]        I85d95015a9ce27a18ccbf73bbbcdbd70;
reg                              If8572800d5d80cc92dd917b60447b63b;
wire [MAX_SUM_WDTH_L-1:0]        I992e7c551b4aa818606c3465d33eb798;
reg                              I24645082ef16129eed1c574f5fc601ca;
wire [MAX_SUM_WDTH_L-1:0]        I2ead0e9941e2280309ab53535b1e1ac1;
reg                              I207a0f6184a0b3be71766a8b47ea5535;
wire [MAX_SUM_WDTH_L-1:0]        I56873feb8418005b5661c7382f2dbeec;
reg                              I5cac08dabbb6de3b01c821d4db93a8e3;
wire [MAX_SUM_WDTH_L-1:0]        Ib6ea4a822da2ea32e0abf6cf8a33d295;
reg                              Ibe6b8c57d7ff47b6fdad5fadf1f6b841;
wire [MAX_SUM_WDTH_L-1:0]        Id1659ccdeaea3e59eb2d3f65a65ebd05;
reg                              I477326720157df2503149125a43ee987;
wire [MAX_SUM_WDTH_L-1:0]        Ic2171967791a0329f3e39fc19d0a6bc8;
reg                              I2c741a5fed7d88e9bdd6b7459feac649;
wire [MAX_SUM_WDTH_L-1:0]        I7d5041a6796c00188f74936d283defe6;
reg                              I17a6511072c7fb4846be5844decf17d6;
wire [MAX_SUM_WDTH_L-1:0]        Iba7608ee0a01af103e022bcaf564bf6b;
reg                              I5ebc3047985651f4b9a957d502a97e95;
wire [MAX_SUM_WDTH_L-1:0]        Iedbe9d0e48bd36064f59faea51afddb9;
reg                              Ifa09fc1b009d073d5a9973b430c63469;
wire [MAX_SUM_WDTH_L-1:0]        Ic3871325d57b310c95ca02fcaca529eb;
reg                              Ie6212a29c7c6b035cfff4c869f945b68;
wire [MAX_SUM_WDTH_L-1:0]        I42f9b1f8ef24ad56c10086852678b456;
reg                              If343015b4815b01dae88bbb6f2017b3d;
wire [MAX_SUM_WDTH_L-1:0]        I3ed5d0fca86f35b3d4b4a89c6147d0cd;
reg                              Ia0116a3cebf94318ed5b287960957ad6;
wire [MAX_SUM_WDTH_L-1:0]        Ib0126fb335e32793c400a97c5a4a337c;
reg                              Id75c23e80cdf25d883806ed20d4ae783;
wire [MAX_SUM_WDTH_L-1:0]        I20590d8fb97ec0b2164ffe17826136a7;
reg                              I1b43f29e0ddb72467befd6f3a9c1c829;
wire [MAX_SUM_WDTH_L-1:0]        I3c128efc9f80c9b8334bf7b61de71b43;
reg                              I3fd0fa3b774d30a267d61e9427d09f3f;
wire [MAX_SUM_WDTH_L-1:0]        Ic7147944f8835e26b9838fdbdc18ca41;
reg                              I2eb08ebaa07a1004638cdd61a7209b7d;
wire [MAX_SUM_WDTH_L-1:0]        I698b1dbc9d8664d1c86c7a763d97b3b7;
reg                              I258c45897919cec5c6acaddee7f3a41b;
wire [MAX_SUM_WDTH_L-1:0]        I508bbade361787127e1a2e8687ec884c;
reg                              Ib42d37576e3aff3d205f1f8822cc58b5;
wire [MAX_SUM_WDTH_L-1:0]        I2afeb2a7b199c0c6738938f156ae4274;
reg                              I1c2ee281cd47a8414851c5e1c758ea65;
wire [MAX_SUM_WDTH_L-1:0]        I86255756ddd1f88b74e070b19f8c3bfa;
reg                              Ie644d131c4f2c603e8e64c5581fdf822;
wire [MAX_SUM_WDTH_L-1:0]        I7d4924388dc5373ad7936dca76797473;
reg                              I9b76f0121a3f7e887e7121db50024ab4;
wire [MAX_SUM_WDTH_L-1:0]        Ie317e5ea2ca4ba2060d0f491290af96f;
reg                              I9eaf4e9ebe07717503ff69b51f0e1905;
wire [MAX_SUM_WDTH_L-1:0]        I56ea52c50a188ec47e48740839a031c9;
reg                              Icb0841ecf142687c3aa23e68f01c927c;
wire [MAX_SUM_WDTH_L-1:0]        Id9b9a8fe43992ec0793845715dd2226c;
reg                              Ie8c0fac00a9de74870e59cbf9e87a39b;
wire [MAX_SUM_WDTH_L-1:0]        I93b69bfb228db4b569a6772179d603be;
reg                              Iae5d6faac1f5685cb1d400ee2b1d85e0;
wire [MAX_SUM_WDTH_L-1:0]        I71afab29cdb962e1f1ca21b61dfb50c6;
reg                              Ib62b02ddf0f57bee49838d19783ef6c3;
wire [MAX_SUM_WDTH_L-1:0]        I9905e2686b350e8a6e7f790563a91294;
reg                              Ibd59d0e5a062f149bd0e91ba76985a13;
wire [MAX_SUM_WDTH_L-1:0]        I524e78ae6a4204e17ba4532dba047d4b;
reg                              I876fdba97e755b74532f7ab191fbac14;
wire [MAX_SUM_WDTH_L-1:0]        I71228fe4188ab1d9796081184a422094;
reg                              I8edf1a08ef943f06ee28771c6e140e28;
wire [MAX_SUM_WDTH_L-1:0]        Ie19b39200436b0bfca13502ad36c21b9;
reg                              I7e12ad8a8ef857e02f4563b2f3a7f0ca;
wire [MAX_SUM_WDTH_L-1:0]        If6657f90c84ca5e2ba08ec705f34be03;
reg                              I17b3a9df6752da6cc987e902e6bbad48;
wire [MAX_SUM_WDTH_L-1:0]        I60ec7459bbe99fce295406bee1f2af46;
reg                              I487496233a32f657171b3789590d0522;
wire [MAX_SUM_WDTH_L-1:0]        I29ab844f80c105d247c5c15faa35863c;
reg                              Ie34534dfd435b3d1cf35e82ca71e83ba;
wire [MAX_SUM_WDTH_L-1:0]        I856fa68463aa5ef1ae53442699d38b33;
reg                              I0e8679271ba733bb87c44b6b9f0b6ed2;
wire [MAX_SUM_WDTH_L-1:0]        Ic3d00a27f15f8983a120395082854d6b;
reg                              Ic14760b65c6fe150c3c48e64389a41d8;
wire [MAX_SUM_WDTH_L-1:0]        I6b1d01c3cb8fb51e43cdb788b89816be;
reg                              Ied6c684cdd280b41ffab93a026d27282;
wire [MAX_SUM_WDTH_L-1:0]        Ib74a56900c1f8b159ad381f61acee801;
reg                              Id0f4dbb72da33748d8baf723c5a32567;
wire [MAX_SUM_WDTH_L-1:0]        Ia5eba52d169755c507b9e0094e467fab;
reg                              Ib0bb71b1f8829347b3a9a7543f9dd964;
wire [MAX_SUM_WDTH_L-1:0]        I0899e8fec1a7209cd94757c0b2f87c9a;
reg                              I47cbb92d2284aef7b9e56e88f0ba6f7e;
wire [MAX_SUM_WDTH_L-1:0]        I08ece7cd684e593e02321612b7a88cee;
reg                              Ic69094123b75ae36e3e54f179a9f2cb5;
wire [MAX_SUM_WDTH_L-1:0]        I691c84d81c60a462e28e2b2bae3ea845;
reg                              I07abbbd75d91018ac53f53e64cffafb9;
wire [MAX_SUM_WDTH_L-1:0]        I58dc9cce6384160c0a85c6efb3319cdb;
reg                              Ib02268d5048c7c8e83118070e927453f;
wire [MAX_SUM_WDTH_L-1:0]        I56bf74b5890ec67090f499afdc0a9c88;
reg                              Idc2a9c6dd8d2aa912548c918c8a488f4;
wire [MAX_SUM_WDTH_L-1:0]        Ibaf2f1f8bda2f6b932dc30f8369c0e1f;
reg                              I5ad7eb9d3ce7c712515254f892d1670d;
wire [MAX_SUM_WDTH_L-1:0]        Id9364a29fd79b52d0442e18dc0227854;
reg                              Ife25829fb3c5023b7d69bbaadf9cf77e;
wire [MAX_SUM_WDTH_L-1:0]        Ica3a41ace27f7d94377981079952f4f7;
reg                              I8b2a79aa4ac88e6b4ca8188a7852022e;
wire [MAX_SUM_WDTH_L-1:0]        Ib57795a63d642a73456324bab41384b6;
reg                              I081e2595b18f306a74d070203447ecf6;
wire [MAX_SUM_WDTH_L-1:0]        Iabf572c97b48c6a7dcc19e56676e3a82;
reg                              I68b152a599887c0039dd9d45c528c219;
wire [MAX_SUM_WDTH_L-1:0]        Iefd370d0df1a93639af482f78a1e8706;
reg                              Id051f1d5454802e0eb37e22248efe8ca;
wire [MAX_SUM_WDTH_L-1:0]        I995d2809ffaf0ecda6a004d01cb9c8c4;
reg                              Ic4c6f707f461cebbc4c93f2ba664ae7b;
wire [MAX_SUM_WDTH_L-1:0]        I4e8ebc46bc068c3f9889d970db131112;
reg                              Ia538dadbd6ae3711740595a18c89b65d;
wire [MAX_SUM_WDTH_L-1:0]        I7b561638da1b4a45ff59be81243e4471;
reg                              Ie7d9730b191781c78391141d95d4f8bd;
wire [MAX_SUM_WDTH_L-1:0]        If0a3b88a66a816b25f17ced5d0e8f775;
reg                              I12f2f886517647044cc251861721bbb9;
wire [MAX_SUM_WDTH_L-1:0]        I0374ada4fe50717f2158468b7ad205d4;
reg                              I615053b36a1851a06125e2ed5ec7f880;
wire [MAX_SUM_WDTH_L-1:0]        I357137b41bb91e0659b1ac6ead9b5c12;
reg                              Ifbc6aa14cd448bbe416897a3671ba857;
wire [MAX_SUM_WDTH_L-1:0]        I5d70bc64cf7b3d3ef4180e082e533237;
reg                              Ie596289582a73e37f78f4ca4cab21e3c;
wire [MAX_SUM_WDTH_L-1:0]        I7d9ad929660cd212387d893266b681da;
reg                              Ifad8c7bacf72583f91be27fbe5b7a1e1;
wire [MAX_SUM_WDTH_L-1:0]        I34be4b353cf75603301372840c2f91c2;
reg                              Ie74c72742807ae4243748fd27d80d626;
wire [MAX_SUM_WDTH_L-1:0]        I14834fc8e6489775359bcecf5a37ff4d;
reg                              Ie7a68c2b368a295f95571bc4a109b9f1;
wire [MAX_SUM_WDTH_L-1:0]        I633a74e4dfa841c9fd13dbb6564c8493;
reg                              Id88a7edf897eea1b4a137141789a04f5;
wire [MAX_SUM_WDTH_L-1:0]        I157bd468200e63385583b9045758d81e;
reg                              Ib13436ad16a37d656d6b1ee95b9aee20;
wire [MAX_SUM_WDTH_L-1:0]        I918c46173eebc5b2a95e041cfd91d958;
reg                              Idc07dc30c0a957e474546ac7a60df38f;
wire [MAX_SUM_WDTH_L-1:0]        I4f8792c18bd07b23e82bbc44b4ca947f;
reg                              I595665d8128bb87ab62741d7ac520a4b;
wire [MAX_SUM_WDTH_L-1:0]        I8d0a1ae4c47edf1f2b99d1175aaa7197;
reg                              I256050251d23250854ff337bef28e460;
wire [MAX_SUM_WDTH_L-1:0]        I734e601f5f9d568a44a48834559e04db;
reg                              I82f0e5a32d1bcd761a74f1f9ce8c88ba;
wire [MAX_SUM_WDTH_L-1:0]        Ie421da1dc5aaea57c50d0c7d9c5a2717;
reg                              I98febac90cccb5fc1f3d966b6e38c4d3;
wire [MAX_SUM_WDTH_L-1:0]        Ief5cbddfbfb98fce4812a676849b9a98;
reg                              Ib534288c2cf976b6ec85db743bc2a823;
wire [MAX_SUM_WDTH_L-1:0]        Id113cab2dd1949d32e3c1c15273185c8;
reg                              If988b82b86db1f4ff6d3695f7b0197e4;
wire [MAX_SUM_WDTH_L-1:0]        Icfe1a689e33b2b9aa9dba692d6d610b9;
reg                              I6ef260ef75e47b011a46ba2080ac3684;
wire [MAX_SUM_WDTH_L-1:0]        Ia4b671f3360f3ce55db0dc0e4d78ddbe;
reg                              Ifc1da524e7670772834d521a6fc4c96f;
wire [MAX_SUM_WDTH_L-1:0]        I60cbd4369e7ba9b6532f279e5c59084c;
reg                              I852d5295a32984af00c95f6d9389555e;
wire [MAX_SUM_WDTH_L-1:0]        Ifb6c65a00d9a2c31d8b1119b949828d8;
reg                              I3c0a621dbef864fd1f566bc2e47f32c6;
wire [MAX_SUM_WDTH_L-1:0]        I4a777f0dd62b19dd340ad31517c4e789;
reg                              Ic04828ba2db8239b093043c27476d345;
wire [MAX_SUM_WDTH_L-1:0]        Ib75747cb32130d44b338ed8c8af8ca11;
reg                              I319012bc6fe93d78de57bcace0caaef5;
wire [MAX_SUM_WDTH_L-1:0]        Ic7e35cf8d5cd230b94c40714f16e2418;
reg                              Ibb35bace971548c9fc98d773d1aff712;
wire [MAX_SUM_WDTH_L-1:0]        Ic51bb9184dfd103703cd0c6ad6edff4b;
reg                              I90023493600924a76d2192080cf6194e;
wire [MAX_SUM_WDTH_L-1:0]        I103f1449c78c47396d6a54dc1c810934;
reg                              Ia9f5ce4603af279bbd9b486b67016482;
wire [MAX_SUM_WDTH_L-1:0]        I56b3a97dc3037f0bb2eed93a9482c813;
reg                              I05721e06a1acdcc0571907c7d853f18c;
wire [MAX_SUM_WDTH_L-1:0]        I51e98035b35a35fdc52f5bab8f19c152;
reg                              Ibfcfd3151af0d82bfce293ada44059b3;
wire [MAX_SUM_WDTH_L-1:0]        Ia6a7f9beaceb08d81012f0e72171252f;
reg                              I9539fcc40d26b13015a864718b116d5b;
wire [MAX_SUM_WDTH_L-1:0]        I21b062856ced09cb9131c01b5e166f32;
reg                              I5490039998187a1a2efc3549e3dee7d6;
wire [MAX_SUM_WDTH_L-1:0]        I4f1221ce7880729fe584b42ef3afe6b2;
reg                              I2b97a79c90f6578c8b2f321f8d598cc8;
wire [MAX_SUM_WDTH_L-1:0]        Ie7f3f1d6cee7f02ae1b17740ed54c049;
reg                              I0c616f736879c28a5222de3d6f49a587;
wire [MAX_SUM_WDTH_L-1:0]        Ib196f5bcf9152703dc32c5101076600a;
reg                              I5590d801fd7fb496019d4c31b7c6d898;
wire [MAX_SUM_WDTH_L-1:0]        Ide9ef5a16d8fe32353c2c2a30e8ee3b0;
reg                              I27e1d2e0e980216b27b90ea48c061025;
wire [MAX_SUM_WDTH_L-1:0]        Iee6f2484a381bd42e441ff072ec582e4;
reg                              I474f6bd977f4197742d0bddb3bece684;
wire [MAX_SUM_WDTH_L-1:0]        I53121a39de0bcba91a4d0438be2ae958;
reg                              Iaa1e981134f5a5c02983c49562683bc5;
wire [MAX_SUM_WDTH_L-1:0]        Iff7950f24f0a6b0073942c37fff49d37;
reg                              Ib051eb1091a85f85a1e50007f1b27cab;
wire [MAX_SUM_WDTH_L-1:0]        Ide86f019e9573706c25bd8b4552396a8;
reg                              I6b5645cdde4b35a16fe3e91d90caaa4e;
wire [MAX_SUM_WDTH_L-1:0]        I2370042234b0e93bb66e44b97fca3e43;
reg                              I8850ab26807dcd55fefadf6310729ca7;
wire [MAX_SUM_WDTH_L-1:0]        If9efe7a1c359ec03014a52870ac13aec;
reg                              Ic5cb81c821716a8aabf8cc2283ff73ba;
wire [MAX_SUM_WDTH_L-1:0]        I6a6eb62960b616043415406ebfc21346;
reg                              I9a6923c6368526a53ef70e16471386ef;
wire [MAX_SUM_WDTH_L-1:0]        I06c7728ef64be8311f48d10d766d0c44;
reg                              I620b8ecdcaccc1ec80ebcf9fa6af0017;
wire [MAX_SUM_WDTH_L-1:0]        I9fe11f6c8147391aa4a5afd1a4e4f731;
reg                              I141cda06bae0c5666e3bc61c6fe5ad66;
wire [MAX_SUM_WDTH_L-1:0]        Id50edc56fce48130247fdbc42eeff9ea;
reg                              Ia9c273b32d0701c7f185ab2de9e57829;
wire [MAX_SUM_WDTH_L-1:0]        If3e5161254eb9056914c46263b865c10;
reg                              Ic3fb524ab434e80b3289c9241b65d224;
wire [MAX_SUM_WDTH_L-1:0]        I58703e8b6d04f8c69ac38f5fcfdc4efc;
reg                              I23c8b64e433af0bd00cef44e38df99f8;
wire [MAX_SUM_WDTH_L-1:0]        Ie1f41720e296ced1b74cb325b666d88f;
reg                              If6a5dc79c0f6ce348956286737a369d8;
wire [MAX_SUM_WDTH_L-1:0]        I5d5701435c96f1078e741921b56e3c65;
reg                              I34e6e9d2153e4a70ee36ab85e72d5318;
wire [MAX_SUM_WDTH_L-1:0]        Id96e744d9b10dcddd1ae0115ea57a76a;
reg                              Ifdabf743a8cb46b7053000ff48ea0c60;
wire [MAX_SUM_WDTH_L-1:0]        I0c0060fe260afa3cdc72f35ffb6938ff;
reg                              I22f5bb821a2571d1764978fd76c8f1d0;
wire [MAX_SUM_WDTH_L-1:0]        Iaec1f186cb4a65da21d41e637fc628f7;
reg                              I1b695aa715615662eff7065c742b0859;
wire [MAX_SUM_WDTH_L-1:0]        I9c15a6a5c0db11ede80ff6d04c9a56d8;
reg                              Iec91b3ca3b54010755d57f8b8ea4a544;
wire [MAX_SUM_WDTH_L-1:0]        I8922487573e02d684a3d71448c3828f5;
reg                              I06ad520cb02e46d34c45f207d42a9243;
wire [MAX_SUM_WDTH_L-1:0]        I47f17afcd5871fc3ac378316fd3d7ae9;
reg                              I9d18ff3465afd8cae63abba68487542e;
wire [MAX_SUM_WDTH_L-1:0]        Ia9642d79bb50567348083b4435c7d66d;
reg                              I914dedc1d5e5e21c9b8d07ec0ecc01f9;
wire [MAX_SUM_WDTH_L-1:0]        I2b2bd845428c49346ef8e94e95b618f8;
reg                              I3375fff5ee0d4b4b12c5a70fbdee59fe;
wire [MAX_SUM_WDTH_L-1:0]        Ib730fdb59198f23d1e590f6d6039e96a;
reg                              Ia8e304ca12c82e41cb8e4de7be199394;
wire [MAX_SUM_WDTH_L-1:0]        I644e83f0a7d432fba38ffb2d99088eca;
reg                              I3566f2779e860008b1a5d305366a07c9;
wire [MAX_SUM_WDTH_L-1:0]        I97f2b15ce0a74e68d5a4438111adcb0a;
reg                              Ie68b31360c12a83c6095254b6f14603c;
wire [MAX_SUM_WDTH_L-1:0]        I84c88b631bed5311cb6e99e58941149e;
reg                              I42ae0c42360c977b35429ce290516a6f;
wire [MAX_SUM_WDTH_L-1:0]        I45c5e6710240685bf54b73b0d7a64271;
reg                              Ibe01835305315fab50269c72ef849b61;
wire [MAX_SUM_WDTH_L-1:0]        I5827bc87b5db1801b7db16e1e61515db;
reg                              Id806a2df1c4519bbbe811791cb4072f9;
wire [MAX_SUM_WDTH_L-1:0]        I1c85c8f73ef80a6808c6aec0c8eca8ab;
reg                              Ifb70a30f8bade95f402e71f95fe6644b;
wire [MAX_SUM_WDTH_L-1:0]        Id13c99b7f7500c8195b54627efbc4232;
reg                              I592a495aecc800236c3470ff8e6adbb5;
wire [MAX_SUM_WDTH_L-1:0]        I4636821315d702a677dc93113872e647;
reg                              I1c8024aa9d81704d2dcf63e34853f8cf;
wire [MAX_SUM_WDTH_L-1:0]        I9c981b0614a29386ca5e8ebc06a17f15;
reg                              Ief03713f5cf37200373a20d42c7fc9eb;
wire [MAX_SUM_WDTH_L-1:0]        I4df3d4dac24877b14e6d361bafc1a800;
reg                              Ic3cb34aae74c5f1a870b3635f8a40764;
wire [MAX_SUM_WDTH_L-1:0]        I913d818403024510c55b65b56a38dd89;
reg                              Ifa3df8b249467cc1e827c69925ef415f;
wire [MAX_SUM_WDTH_L-1:0]        I57015930f5b09a6c6b030ed01dad2177;
reg                              Icf3ad912aaeaa0c5cd1ab0edb898d6e8;
wire [MAX_SUM_WDTH_L-1:0]        Ib54d55a70605119e37e9898b940ff636;
reg                              Ib774f380e3d7cfd1f5f064e93d8134b4;
wire [MAX_SUM_WDTH_L-1:0]        If7e146da4f3bd255b8457fd6902005f6;
reg                              Ic07c650e6e49892a41cfaf3a37471426;
wire [MAX_SUM_WDTH_L-1:0]        Ied00d87af99ae55144fdde41ebfc1357;
reg                              Ib1073489d63ea33d7f3892f4ff875358;
wire [MAX_SUM_WDTH_L-1:0]        I7774313f1ae5a2de98855aad572b3676;
reg                              I174b6c36f2af82f8047cc76543a3b4ee;
wire [MAX_SUM_WDTH_L-1:0]        I679baea452c3c6d04c53baa88edd8eb3;
reg                              I953b975a89adcc88039284970e9b3404;
wire [MAX_SUM_WDTH_L-1:0]        If4132b39ddb92aa02d8d0346fb0e6691;
reg                              If2b40d249c531e10cc22d1335f350441;
wire [MAX_SUM_WDTH_L-1:0]        Iba70e737d52e6812a67c159520e5192f;
reg                              I44ccc3ae897109dd51f9afeef93daca4;
wire [MAX_SUM_WDTH_L-1:0]        Ib9ceb8315f0cd848f861bab677c2c694;
reg                              Ie9236599cea94cfb603c6b977fdbb44a;
wire [MAX_SUM_WDTH_L-1:0]        I7846bc2cc11e08d05f7c853c4920d555;
reg                              I25f1ee9cee4d04bd8fec1fe601d016d7;
wire [MAX_SUM_WDTH_L-1:0]        I0865623d3350645e63fa6e6c9b78ac57;
reg                              I5ec1e530b9007a75a778af4d82ab427b;
wire [MAX_SUM_WDTH_L-1:0]        I0262b30a4efa9f1cfb11d1c3940de9e7;
reg                              I8a9e516aa824260998d10db758642bb0;
wire [MAX_SUM_WDTH_L-1:0]        I7a2e79d42779ad235bca6ce3757cf588;
reg                              I70dd1350d65155ee7b562f4c79024a3d;
wire [MAX_SUM_WDTH_L-1:0]        I09e9a3cd4c12d204f760758e873a177b;
reg                              Ic9146d8b3dd0c612073b70b8a8791e8c;
wire [MAX_SUM_WDTH_L-1:0]        I30b0b1d54912c1a41a02a25ab238bb54;
reg                              I857d3155df0b6dd704514b039c66fa97;
wire [MAX_SUM_WDTH_L-1:0]        I49fb0909ddf66fc0073e6400f1a07844;
reg                              Idc1b8aa2f81a7fbd87e4f5821d14bf01;
wire [MAX_SUM_WDTH_L-1:0]        I9938397dc94002481984f5b560fadc58;
reg                              I68b585571699a57bc6ba5e8955467119;
wire [MAX_SUM_WDTH_L-1:0]        I4378d139db4b710e3587aa72df22b70d;
reg                              Ib70e99c3acc76286a6811bcacc9284de;
wire [MAX_SUM_WDTH_L-1:0]        Ifa43d74fa91b7b9884969f575ef9ca8e;
reg                              Iee17ece482d04964d3c21a092ec955a4;
wire [MAX_SUM_WDTH_L-1:0]        I7c19a79f441ecbb73685db5a505e7479;
reg                              I5a247475beb737d470f03507e55f5b24;
wire [MAX_SUM_WDTH_L-1:0]        If2af8106efc1f7dd02c074af68278b3d;
reg                              I13b0c9578f7b6b3b7e6704d7b44079c4;
wire [MAX_SUM_WDTH_L-1:0]        I89a3f8d5f760d1a650f85814cbfdc017;
reg                              I41eff06fe1dea8be4613945de596d3ca;
wire [MAX_SUM_WDTH_L-1:0]        Ifae345c79662c3df3dff0fe68ad68746;
reg                              I08f22261d5713c0636d77c7938f592d6;
wire [MAX_SUM_WDTH_L-1:0]        I88a61cf72347d695489909d0819332ab;
reg                              I1c7e41b9cb1bdb6f649c88c0ed3f4100;
wire [MAX_SUM_WDTH_L-1:0]        I9aaa036a6158d11c235bdc8406d79f4c;
reg                              Idd59a5357d4c835379ed180ac0924bf1;
wire [MAX_SUM_WDTH_L-1:0]        Ie8df350430970b5f1229cda772440f85;
reg                              Ibe7e5c2cb9c50eca34a3859d13e83a92;
wire [MAX_SUM_WDTH_L-1:0]        I7d77ac9b64b2e8cae21c6e36947e3ca2;
reg                              Ibf5c141c5cc0a6a20c05b52bf8282476;
wire [MAX_SUM_WDTH_L-1:0]        Ic1faed76fca5a9ceb7db26c2f43623d9;
reg                              I0038305f94aaefe2cd1a243580d95932;
wire [MAX_SUM_WDTH_L-1:0]        I3ca2b9b77ed8d78a10aff42a07a53b07;
reg                              I5364deb983adc2ae505ed2b8c57f876d;
wire [MAX_SUM_WDTH_L-1:0]        I1f00849ea055a7893df386aed162a7b6;
reg                              Ifdb5589982db805a0416e1c01276249a;
wire [MAX_SUM_WDTH_L-1:0]        Iaf8a19fde3de660c3fa925593bebbe0c;
reg                              I8bb5522183b65583fda83067990b3e94;
wire [MAX_SUM_WDTH_L-1:0]        Icd1da43a4d95230e79dbd35a7ae41066;
reg                              I1e77fe6aeaba852aba34ed37dd53add6;
wire [MAX_SUM_WDTH_L-1:0]        Ice9079fb6e08d629f8c0c9ce332c8f11;
reg                              I9171019227f35760d02d0c8ce786f4d3;
wire [MAX_SUM_WDTH_L-1:0]        I15fafe2baba4d2f28037023a81ce0a81;
reg                              I6e92a48aaab94074a555efa9bd1e7243;
wire [MAX_SUM_WDTH_L-1:0]        If4d5b48882e9e628cf51ad2ac2f38c22;
reg                              I3bc094d67805664859fdcb66f1360e64;
wire [MAX_SUM_WDTH_L-1:0]        Id0eef1adba01447c14a6f005782dd9a2;
reg                              I2518ccf385b3b677d95983bc550282e8;
wire [MAX_SUM_WDTH_L-1:0]        I1d1a7c5928982c278d068ebd262254da;
reg                              I7547c56b32513ad45d775b4502596d9d;
wire [MAX_SUM_WDTH_L-1:0]        I6354a0e638340378124e4df7f3d145b8;
reg                              I013d84bfd582acc7accf07ec522961fa;
wire [MAX_SUM_WDTH_L-1:0]        I0236c912c6d684bf4862b725be9d5951;
reg                              I0ec27b590ee6dcdd9c1086105e3b6c23;
wire [MAX_SUM_WDTH_L-1:0]        I6f3be51d69b2b64a04e55b8946d5dd56;
reg                              I4cdc955fa9afc75c2c977de4ec540e1e;
wire [MAX_SUM_WDTH_L-1:0]        Icde3e6dbcf985682041f30903ad95572;
reg                              Ieefbb5d6f4ac1e586832c5c0f513c5a2;
wire [MAX_SUM_WDTH_L-1:0]        I46ee30b46020d91707689f3468f00e26;
reg                              Ic828cdd5dfde844df4c150921af2a443;
wire [MAX_SUM_WDTH_L-1:0]        I2605f078c1a9006c93855a9a2b0cf6b9;
reg                              Idf1ecab26889c4adcb835fda6b1cb368;
wire [MAX_SUM_WDTH_L-1:0]        I4d226dd2f0bfcdbea6a2e6a6613c1b64;
reg                              I00d3f14b20e1ea7d726533386e0eba27;
wire [MAX_SUM_WDTH_L-1:0]        I5c942076b173cf527e1be2ddb8560e84;
reg                              I7f720a18542528f0c9bfb14f699ff4da;
wire [MAX_SUM_WDTH_L-1:0]        Ic95191bccb18e26c10e56be395ca6b1a;
reg                              Ia98a6f01e4eb5bc74d50d350e79be426;
wire [MAX_SUM_WDTH_L-1:0]        Ia284f974dd8a526f31eb81ed71a06e94;
reg                              I182b43872d50de6f7afb700f178b160e;
wire [MAX_SUM_WDTH_L-1:0]        Icc93450a007cee4c0a42717ed7600528;
reg                              Ic9b72b2a91d951cf08cf54ed215ecaa8;
wire [MAX_SUM_WDTH_L-1:0]        I9ec9f389d0489908d497487e44c6edcd;
reg                              I93084ccf5b5e4efaee968b497bb2a775;
wire [MAX_SUM_WDTH_L-1:0]        If8a527cc7f06a9963a80a880d225d34c;
reg                              Id38852415486e6989b89a0d85ad6771b;
wire [MAX_SUM_WDTH_L-1:0]        I39ff4663007dbc89b403f3b08a69bb6c;
reg                              I17cf58ef5326978c62c03c56090a299f;
wire [MAX_SUM_WDTH_L-1:0]        I9590eb28a81c730b83b92ef7653e71a1;
reg                              Ie41ca18c7d11a47e274f9c33f75393ec;
wire [MAX_SUM_WDTH_L-1:0]        I2ba1acca919bddcc22a41a28d43a4e3e;
reg                              I7b80b4902fe98c10dd72c9eb082346e5;
wire [MAX_SUM_WDTH_L-1:0]        I62d8efd4227cb3dc88aa08b6585fafc8;
reg                              I20ffba20af04b99954bf719589e90d1a;
wire [MAX_SUM_WDTH_L-1:0]        I749e987266a20840bb8a4b1a2a2fc5b0;
reg                              If8fe5af7e5c3c97b5a713f6bcf919f1f;
wire [MAX_SUM_WDTH_L-1:0]        I7607af5d98e8070e3d15cee23cdf877e;
reg                              Idc5fb0f3a04ab32948e249e088a11b11;
wire [MAX_SUM_WDTH_L-1:0]        I2e11a697d7f17ac30302eadb500de72d;
reg                              Ia9f1e580e8f441394d719d52a7bad688;
wire [MAX_SUM_WDTH_L-1:0]        Ia0886ce792e062e22d0c224158cdfb7d;
reg                              I02849282dd1bd663fd39baccf41762f9;
wire [MAX_SUM_WDTH_L-1:0]        I6b3cd79aa87235ff174c0299b855dd3d;
reg                              Ie4cda4648f6ceb76b8fb74f290ab6439;
wire [MAX_SUM_WDTH_L-1:0]        Ie4ae993ddb776bdffec843db0def2f5c;
reg                              I24135210c23b2422a42c90ee25594191;
wire [MAX_SUM_WDTH_L-1:0]        I3ed2da9b53daac0852a06ad1acfad21b;
reg                              Ib08897f9216599042f7b97b137e07fe1;
wire [MAX_SUM_WDTH_L-1:0]        Idefa29d4d4e2a6e9147f84893520096f;
reg                              I51e14ece9ab6607f83e6ba27f3f046a9;
wire [MAX_SUM_WDTH_L-1:0]        Id1fbbe0594dae272856566522633bb3d;
reg                              I7a626ec321bf963a5401892a7e3891c7;
wire [MAX_SUM_WDTH_L-1:0]        I8070a3b7d8b1a7ae90c1a2d27aed09aa;
reg                              If76f04fe0baf171d7df2c0cd849aea2b;
wire [MAX_SUM_WDTH_L-1:0]        Ie88285ce2b9c71de02ebd62e8f44ca72;
reg                              Ia9c8cc5e3becf3d48feedec8fa2c93a4;
wire [MAX_SUM_WDTH_L-1:0]        Ica1997c6c569c1d1f45224fbaa4e6b59;
reg                              If3b77c41fabcdb283f2c6fdacaa5e9a4;
wire [MAX_SUM_WDTH_L-1:0]        Iaf08bcaaeb15bb0c971432f7f8b16d0a;
reg                              Ie5373b01a92f2ff85be8077cfef2175a;
wire [MAX_SUM_WDTH_L-1:0]        Idcb37cfc357cc088c775409fb9225b51;
reg                              I5109afc4dc91780e05704ea5e1399e3e;
wire [MAX_SUM_WDTH_L-1:0]        Ic419255414995e7168afb97b051fa64f;
reg                              I3e0b41bee4c76eb5f3340ad23bfa01ad;
wire [MAX_SUM_WDTH_L-1:0]        Iee6da3120d73373627b25ab7c0dedd28;
reg                              Ic0732810fd355d59a3168be896a0f9ac;
wire [MAX_SUM_WDTH_L-1:0]        I56fc99a22960232b305d6e683c66fcc7;
reg                              I220e32641265b46527ca61111f7ebf1b;
wire [MAX_SUM_WDTH_L-1:0]        I0a9a09b0ab43d2a0f1d1d01e13f0333c;
reg                              Ice59d2af73d0b0f2ae91a2ef0c2b7f04;
wire [MAX_SUM_WDTH_L-1:0]        Ibc73d07e0c97a6fcae791e04106cb082;
reg                              Ic308610ea8bb62ecb6094192e02dbdba;
wire [MAX_SUM_WDTH_L-1:0]        I224bbdf94ac86c5c376d1db4f4d4e060;
reg                              I33ee415d85e2bcd8f975d34b880f6ea7;
wire [MAX_SUM_WDTH_L-1:0]        I43f2b69c6b427de3095c44d4166b77cd;
reg                              Ie61f299252b8fecfd3e8634b64df5a90;
wire [MAX_SUM_WDTH_L-1:0]        I1e50c90010a3df1a8ce1cff811cc7a0c;
reg                              Icc67656ad2dd3fffae4e5abe02f8fff9;
wire [MAX_SUM_WDTH_L-1:0]        Ie1817cbf3a80dae435a5571dfbd2f5ad;
reg                              I0c47ccef4b55410286248884a7249703;
wire [MAX_SUM_WDTH_L-1:0]        I0052d562fb3182890c8828e52d437b11;
reg                              I94e4041b482064334fd0ed92b91bde89;
wire [MAX_SUM_WDTH_L-1:0]        I1eedecb1d8ff505c75be7787199afada;
reg                              I39d3bce4060032a81e6b6a1c1805cfe8;
wire [MAX_SUM_WDTH_L-1:0]        I7ef544597a185b1de63b4ffc4a1d44c2;
reg                              Ifb422c30663eb4824caa72326b238df6;
wire [MAX_SUM_WDTH_L-1:0]        Iadeedf3870f0b1eae98d0f7dbbeff04a;
reg                              I41ab6fb6ec6ef7ffff70e50f25f217b6;
wire [MAX_SUM_WDTH_L-1:0]        I70ae07db9b44d530be220f06401d3d3d;
reg                              I3ce10718a2211184999663c3c2493cc1;
wire [MAX_SUM_WDTH_L-1:0]        I7992ea31927b4f0e268462a3b0f18c5d;
reg                              I877e8d94236c3d8b0a31858a98fba5d6;
wire [MAX_SUM_WDTH_L-1:0]        Iadf927d18644a232ad1f1eba7db82934;
reg                              Iff2f1716cbd73b406d8f07c22dc79fc8;
wire [MAX_SUM_WDTH_L-1:0]        I2a9c673cdd7ded79e09ada38c0f47e6f;
reg                              Ibc48fabc172f27ebce18d0a9b5120dc5;
wire [MAX_SUM_WDTH_L-1:0]        Ia86740e870d8063f0266b68ad6d7481d;
reg                              Ie562ebb336e476a81f20a652d4cb20f1;
wire [MAX_SUM_WDTH_L-1:0]        I6627bcdbaa8afb115123777abd45435b;
reg                              Ib5ee5a6ffc45ed1fece0822dc4619b57;
wire [MAX_SUM_WDTH_L-1:0]        I96fe3eb633eff6958ac575b997460bb9;
reg                              I86ba73ee348f80e2f9891d2ebc8a02ed;
wire [MAX_SUM_WDTH_L-1:0]        Iefdcb71f2903b11f5cb0b8857f7a1727;
reg                              I1e96d5af3d0e3fdce39530dfd0131a7d;
wire [MAX_SUM_WDTH_L-1:0]        I2eb90278aaa54b9c8212b3b4af7c3617;
reg                              I38352b363fa37f6f822fbc1a39100968;
wire [MAX_SUM_WDTH_L-1:0]        I43493f70f0336453d77caf7f27503daa;
reg                              I4ba41864bb1d2130c6971e0b2903027a;
wire [MAX_SUM_WDTH_L-1:0]        I26a7fe395eb583258c1ac58aaaa3234a;
reg                              Ib68deeb7bec4ca3585d1a4dcbf8793f1;
wire [MAX_SUM_WDTH_L-1:0]        I21668ff77cf75570cae97f575cbcf644;
reg                              Ida3d808d100e0bba290f96ed9e744e65;
wire [MAX_SUM_WDTH_L-1:0]        Ie48be9e6b6fd63baa104d0a6a4561a1a;
reg                              I4d4901ff372f6820ca9c8c29cefa664a;
wire [MAX_SUM_WDTH_L-1:0]        I05370777439b01811fe7f750d2f724f4;
reg                              Ib99e1b93fb7fbda260d93eea3d24c3e9;
wire [MAX_SUM_WDTH_L-1:0]        Icdcd83341f6b5c404f91ec7e97d0550c;
reg                              I019e399a1cef87745e025a7d74e94db0;
wire [MAX_SUM_WDTH_L-1:0]        Ibba4e82d1510ddc16eb4ef64893cec02;
reg                              Ia8974083bfd064f2c27dcd421490fcfd;
wire [MAX_SUM_WDTH_L-1:0]        Ifb00ae47340bc99669c71da34cccc59e;
reg                              I8fd5787ebf758919e7cb75d7419441e8;
wire [MAX_SUM_WDTH_L-1:0]        I75a4cf2948bebc58e12bb039ed273ff2;
reg                              Id14074d5230885c38b89b09b130ecf68;
wire [MAX_SUM_WDTH_L-1:0]        I5a9fdec7d7ff99fe33ad6cd8afd9e059;
reg                              I86fefad34d3c864dd0e725133f303b4f;
wire [MAX_SUM_WDTH_L-1:0]        I47b1695a74e4d27389b97543415dcc67;
reg                              I1ca188bcdebbf41d84f7a5220bd1d195;
wire [MAX_SUM_WDTH_L-1:0]        Ieb38fa62119a5a77c060d6634e051298;
reg                              Ifc640243288c9b37b7eb9e00351b23f0;
wire [MAX_SUM_WDTH_L-1:0]        I3459d98131faef5a5040a03847890b55;
reg                              I3d149293f106ae8680c7f4702daa0bd6;
wire [MAX_SUM_WDTH_L-1:0]        Ie9b9221b2122087cd5f309570b6d31ca;
reg                              Ie232799bd6c4ec99e24c78f3ad798265;
wire [MAX_SUM_WDTH_L-1:0]        Id4451722e8e2393d627dcd0175dc9903;
reg                              Ifebcf64858d5e2d07ad7894d6182eb11;
wire [MAX_SUM_WDTH_L-1:0]        Ic10356f9069e3651b9c045c906e63512;
reg                              Ibab55499323660588ec82ebd07ab0572;
wire [MAX_SUM_WDTH_L-1:0]        Ic3a431f39c678b7175ed30fde1fa6424;
reg                              I89af7644c48a80d7d22f50b008d35841;
wire [MAX_SUM_WDTH_L-1:0]        Ib01cfd833a63500e03333f263805db3d;
reg                              I0152dc6e6a7acd72a2144623e63998ef;
wire [MAX_SUM_WDTH_L-1:0]        I0b7b4c0a8503c751229edfe0237cc903;
reg                              I951dedd7af44c3865a8f36888432d0c9;
wire [MAX_SUM_WDTH_L-1:0]        Iace01234164c8a9f7c98eeb83268745b;
reg                              I8188dd7cb03854c6f709de06ff785d91;
wire [MAX_SUM_WDTH_L-1:0]        Iace8b3b3a4c16763132b5aaa6b24212d;
reg                              I3b30b4ab00a49e10a75587aa324d6132;
wire [MAX_SUM_WDTH_L-1:0]        I80a89644e278e96b1cd1c4b7f764dc34;
reg                              Ie50aca688b3433fad7565998cb900155;
wire [MAX_SUM_WDTH_L-1:0]        Ia92d2276a8a23521ad1b88df7c27bc2e;
reg                              I3342fe0c5d3ee5021892d53eb45bde21;
wire [MAX_SUM_WDTH_L-1:0]        I39bbec42c442d1e8c818f46ad9c096a8;
reg                              I5134b762ac428bed07ce102d8927a418;
wire [MAX_SUM_WDTH_L-1:0]        I88f1b5c12759a5efb2d2ded8483c9ed2;
reg                              Ic14f948884da19a272a4760ffaab9ea9;
wire [MAX_SUM_WDTH_L-1:0]        Iaf4ae293c576af16f5f43a8b86c1aa3d;
reg                              I46e1047bca2b38e62b4de80d1d2249de;
wire [MAX_SUM_WDTH_L-1:0]        I68b575fcbc5321d4d26a22bcdbb506f6;
reg                              I866b30a63b3b5fb708934a1cbb0e1d9a;
wire [MAX_SUM_WDTH_L-1:0]        Idf600b93ee1018ecf969ed7944b6bc7b;
reg                              Iaddc1f2e822fd2fe9d9046d759a82cb4;
wire [MAX_SUM_WDTH_L-1:0]        I1cd93172cf5996bc870063aa642188a2;
reg                              If9285bf7611bcc5ea6432215c349e021;
wire [MAX_SUM_WDTH_L-1:0]        I4af080cb4e5cc525db95e5f401019e8c;
reg                              Id277f5f05551eeb5dec1701056330da1;
wire [MAX_SUM_WDTH_L-1:0]        I6fc8044eb226a14ff1a786ddc96d2414;
reg                              I9963d0b24763ed8038b1f3922b8f9548;
wire [MAX_SUM_WDTH_L-1:0]        I27fd0073dbcdee599fbe85cf48806efc;
reg                              Ia98de3691917dfb63bebdc3f8655c8be;
wire [MAX_SUM_WDTH_L-1:0]        Iaee6d725a8b2653eeac6d5acb91f8f36;
reg                              I0bce960fcc58938e6a1e01b912eabbf2;
wire [MAX_SUM_WDTH_L-1:0]        I4afdeba4fc2a12a6cbe3567a519367fc;
reg                              Ice5f7168aeb940d48093cc9df7cba36b;
wire [MAX_SUM_WDTH_L-1:0]        Ib42816335dd8475dcc78662c4c0786c1;
reg                              I859d795a7d141eb777c1f3c038203794;
wire [MAX_SUM_WDTH_L-1:0]        I343c9efe71164c01e9c7d599e032864a;
reg                              I0dccb8eaad52ce4d780696a8485420f1;
wire [MAX_SUM_WDTH_L-1:0]        I108c269ceec4adcff9afeda01101b838;
reg                              I6d4fc81ced37c159303c243af04d345e;
wire [MAX_SUM_WDTH_L-1:0]        I761983331fb6e3c6c437b3f1660f0b6b;
reg                              Iefdb8bd28839af9413a3906cbfe715e6;
wire [MAX_SUM_WDTH_L-1:0]        I70d32affde22f9dcb2d77430fca39069;
reg                              I0615acb0f7cf79b5f6ae8e91cb525dc9;
wire [MAX_SUM_WDTH_L-1:0]        Ic08e85346f61da036a15345a13ac12f0;
reg                              Ieed4c810a5bb69de112522dcf00b16ed;
wire [MAX_SUM_WDTH_L-1:0]        If5dfdadb3868ed5a495007362f7db648;
reg                              If533578cacb685a95afbb8e1c05d3c07;
wire [MAX_SUM_WDTH_L-1:0]        Ia1ee5579358b564de06c08ca418a9bf4;
reg                              Ia858ff5551286beffd4cf82f876d30ac;
wire [MAX_SUM_WDTH_L-1:0]        I9bb81dda8102b829441be46460eb8900;
reg                              I4c66570630a650fa7b9bec543f685487;
wire [MAX_SUM_WDTH_L-1:0]        I8eef6ca0a61a21882ea28b3d63735228;
reg                              If10f33385e236eaba56cbab8c2883399;
wire [MAX_SUM_WDTH_L-1:0]        I438522d92cce6f7010246424746ca255;
reg                              I7cb58e4c486e683faa4acad4756815d5;
wire [MAX_SUM_WDTH_L-1:0]        I92496f68b44a94565af28a2c28d6fbae;
reg                              I452e51cca9acec44e36e4efd21b43034;
wire [MAX_SUM_WDTH_L-1:0]        I66528f43f614f0edb715564eba3c77c1;
reg                              Ice0234f25de4ab1f03a3cb01a2d61dbf;
wire [MAX_SUM_WDTH_L-1:0]        I8cab9fba615b94fd4bb6934325be8ab8;
reg                              I12a18a1f8d4416e9bc8abee6ac3dacfc;
wire [MAX_SUM_WDTH_L-1:0]        I92d9fec22d36b1baac8bd78abfc1bbd5;
reg                              Id17ada8dae3f9810d1892d34f2288859;
wire [MAX_SUM_WDTH_L-1:0]        I4eadce87f47df6d8f0e4acd057de5a09;
reg                              Ia2c5fe53cb5b318fa63d09881609655f;
wire [MAX_SUM_WDTH_L-1:0]        I73203143fe37933c16fff873c1abf512;
reg                              I579c7926e7b78f4ffc606adc10522f53;
wire [MAX_SUM_WDTH_L-1:0]        Ibed2a63af723a7abf96dacf1951e5266;
reg                              Iffa06a336949f56f4e5a88a06d8b7e60;
wire [MAX_SUM_WDTH_L-1:0]        Id667c80003b5541de9f84d3b8709c828;
reg                              Iaf82668eb49248709540f2f529f1b3e4;
wire [MAX_SUM_WDTH_L-1:0]        I02cbb4255db2b21ea32140f9e9ddb36b;
reg                              I90b3708abdf742370f06cc513ee307e1;
wire [MAX_SUM_WDTH_L-1:0]        I65354f2069de0c25bbe7cd50fbe892aa;
reg                              Ia17906696bd0e095d7a5297da2e049ea;
wire [MAX_SUM_WDTH_L-1:0]        Ic279867ebf3055980f3d813d5dc8dec6;
reg                              I180d4f3b23b518271d7cb8189fbeadc5;
wire [MAX_SUM_WDTH_L-1:0]        I5c05da8a222ad5effb9815cbf3ec25f3;
reg                              Id79636d195efff260c430978f0bcee9c;
wire [MAX_SUM_WDTH_L-1:0]        Ib8bf21f32c0e8b9cfa42a53807bfe3a3;
reg                              Idbf4ad11ab2a27044193448c8739fec6;
wire [MAX_SUM_WDTH_L-1:0]        I7208256bb198bfce1be71390b01bc028;
reg                              I3051f561a5e1131ebf167cb6ccb5adf4;
wire [MAX_SUM_WDTH_L-1:0]        I49f2a06ceb3a59773c65b19f54ff362b;
reg                              I9322a2a61900943075bbc23c72a3f65d;
wire [MAX_SUM_WDTH_L-1:0]        I86e495dc894d2aace15c1aff89798bf7;
reg                              Iedc463e359dd3003d9f7e50f3e858e93;
wire [MAX_SUM_WDTH_L-1:0]        I0d53bb5344cabe5fa5ce3ecf7122a260;
reg                              Ie7cfdd25541414ff3f8d6e5d7677fbe5;
wire [MAX_SUM_WDTH_L-1:0]        Ib2f5f5fc77ea8b529f2471c54388f2d1;
reg                              I1e93f0470d2818249f1c28ef2a399a0e;
wire [MAX_SUM_WDTH_L-1:0]        Idcada1bfb3c0d1f2a09aab58a2071a57;
reg                              I5d6e576b0fa7e3219aaf9ccc345085b8;
wire [MAX_SUM_WDTH_L-1:0]        I814b62120953991f9da055f118967e05;
reg                              Id962beade26396738ba0e97f67d5e261;
wire [MAX_SUM_WDTH_L-1:0]        I123a212546a8ac394051425db4924812;
reg                              Id0ab747d92288f23cef793567b2363d1;
wire [MAX_SUM_WDTH_L-1:0]        Ie95f1a7e0effcec0aa423dc803056a13;
reg                              Ie536879e6fa9be65376d7f00e0fc40d0;
wire [MAX_SUM_WDTH_L-1:0]        I106deaff50b8480eac31ddbae2ec7c61;
reg                              Ibf312ae4f51fbc44b43848f9df62a45f;
wire [MAX_SUM_WDTH_L-1:0]        I68528be9951f5b8805411711cd11ea59;
reg                              Icfc03646b36b971b9fa57d04a26dbfc4;
wire [MAX_SUM_WDTH_L-1:0]        I0f034a8f077b0ab231727b6298e366d8;
reg                              I4f134c0669b5a6a8c7e03be7eee30c6c;
wire [MAX_SUM_WDTH_L-1:0]        If9c12f8662333fb54a45cfa1bc5da487;
reg                              I6c765e677f42fe600b848698c8a78349;
wire [MAX_SUM_WDTH_L-1:0]        Ie1681d905517daafcc7584725cd6014c;
reg                              I284b23051c85300c2a1e3afe8f25e99e;
wire [MAX_SUM_WDTH_L-1:0]        I2ff3edcdb6158f1e3c9a555aeefc0850;
reg                              I9b560d9baf8a7422b0dd84720e924ced;
wire [MAX_SUM_WDTH_L-1:0]        I43b380be6df7df0d354223d0a0d6d6b6;
reg                              I457ae11ad90c8478751eb4b42764e158;
wire [MAX_SUM_WDTH_L-1:0]        I23eb1dc4d1c992f804dd04a2d823c778;
reg                              I2b7822d5d77aaed61eee87570564df76;
wire [MAX_SUM_WDTH_L-1:0]        I7f90f96c0260560ad5e6dc7448b2670a;
reg                              Ibdad0ab78e4404c852e60a2b04c3a5f6;
wire [MAX_SUM_WDTH_L-1:0]        I07b417cdcc99eaea3413f563e26ddc73;
reg                              Ic4efba3932e598784f5b9ad6ad04772d;
wire [MAX_SUM_WDTH_L-1:0]        I2f3ab9654e515a54e22e73d6c130ccc3;
reg                              Ia03836a4e93d2f36513227d1dfaea0fa;
wire [MAX_SUM_WDTH_L-1:0]        Iebdc41368d57498a04fa73e30b10a966;
reg                              I138fb0c48f2d27e3315e237d9e61d653;
wire [MAX_SUM_WDTH_L-1:0]        I5b4305bef5b4350c1d7ae143667afddd;
reg                              Id0b1c46fa4caa63a4c63a44ba3c5ef8a;
wire [MAX_SUM_WDTH_L-1:0]        I2795d21d343b83a69146314a2407cfa2;
reg                              I3566033cf5c9a06977c9182925750707;
wire [MAX_SUM_WDTH_L-1:0]        Ic6386d7d8813731d612e24b715740275;
reg                              I02812a8a833bb69eb168a1004b6fafdf;
wire [MAX_SUM_WDTH_L-1:0]        I4c366a57920ff090a98a2cb8b9caa00b;
reg                              Ie886c5effc85f1fe0b6411db4a2cde77;
wire [MAX_SUM_WDTH_L-1:0]        I14cf5d43fc9864820a8a25efcc5c6d86;
reg                              Ibab1d13cd6a4f7b0c79c9f845339e53f;
wire [MAX_SUM_WDTH_L-1:0]        I33b99994abbb5ecf8eed4de39033e4f8;
reg                              I7b813d83b13bb7bc13940cf5714c06ba;
wire [MAX_SUM_WDTH_L-1:0]        I7c3291f0250d13ca94802b0b071a95c6;
reg                              I09031235f61238b0e32ff52641aab70e;
wire [MAX_SUM_WDTH_L-1:0]        I2c926fd9d306e9ae13364e07c4b0395b;
reg                              I5402fd208dc7ca81dfd2920a9cfa2715;
wire [MAX_SUM_WDTH_L-1:0]        Ib23edc35fa5bbfe0415fcf0861a22d9b;
reg                              Ia01c82761aeb124cd92fb15ee367ee8b;
wire [MAX_SUM_WDTH_L-1:0]        I3e0e682047f7cc36142e668828cbff1e;
reg                              Ib1a40247057324b0bd810c844bf11f51;
wire [MAX_SUM_WDTH_L-1:0]        I99fb9030e8361e57818c07511479a9b8;
reg                              Ied8bd4b6fd0e4fbcced6d20eb7435f55;
wire [MAX_SUM_WDTH_L-1:0]        Ic87c3d7762a18772972552162e1d1a8c;
reg                              I4ee312036de8c08300c358edcff1e1e9;
wire [MAX_SUM_WDTH_L-1:0]        I7e393e6c1d1bc44daaab120d55f5dd59;
reg                              I477a920e2326828bf026b0a6b6a18e2b;
wire [MAX_SUM_WDTH_L-1:0]        I448f126fd3932d5065abbe7bb2d92c56;
reg                              Ic11a6b77b84c44180eb99220a0c4c9f6;
wire [MAX_SUM_WDTH_L-1:0]        Ifc8c6df8904b97674f2970ebc95b523c;
reg                              If0970d9f7b053fce3ced3521b4885588;
wire [MAX_SUM_WDTH_L-1:0]        Icd0622a90782b9c451950e7ab0399567;
reg                              Ic7ebdc317c978eb275eca41d5b9106a5;
wire [MAX_SUM_WDTH_L-1:0]        I6493b3c087d4685a6b3f98c73dc2ff49;
reg                              Ibe3d3e6bc58efc2e9d9eb1f96cdfe424;
wire [MAX_SUM_WDTH_L-1:0]        I20c2057240417146df144b518b43d052;
reg                              I1dd4671765f8826c2fe20c592c5e32c8;
wire [MAX_SUM_WDTH_L-1:0]        Ied029d0bdea3bf134744c99426fa72dc;
reg                              I6cde57127c5bd2732e71ecb7738fad6d;
wire [MAX_SUM_WDTH_L-1:0]        Icb82c9ff4cb58159a1c3115c6fdd5f8c;
reg                              If6ce2fa9f0b8bc74442ed8262b5089cf;
wire [MAX_SUM_WDTH_L-1:0]        Ia3450e134e4086c35acbdee1e6042396;
reg                              Ib0001d7298ad1f3b1c7603173a70d8b5;
wire [MAX_SUM_WDTH_L-1:0]        I5a0f27df5158309f32f0df31e8ae3ae3;
reg                              I05e739fc87e962848f265e2c73338cac;
wire [MAX_SUM_WDTH_L-1:0]        I17d9e19854cef197fd3267618617efc3;
reg                              Iaaaf373f7e6f55214915b93da9bd71d3;
wire [MAX_SUM_WDTH_L-1:0]        I2993acb61f1abe529f8a60c94a438550;
reg                              I47b0847946b0e00961233ac0101fa2a7;
wire [MAX_SUM_WDTH_L-1:0]        Ic8be2c94235fb40f78da33179ce4873a;
reg                              I2f23d4cdb6f5f827513aa60266936e4f;
wire [MAX_SUM_WDTH_L-1:0]        Ib3367565e4456da15e7c2315dccdb5e4;
reg                              Ia67f9b902a21de0414eb8dda52171991;
wire [MAX_SUM_WDTH_L-1:0]        I15a1671def323cd294591564ae6ef8b1;
reg                              I87b10521099179c18652c86d5887c908;
wire [MAX_SUM_WDTH_L-1:0]        Ic512effb493a06ece58a2af155135004;
reg                              I84057a3b319ab3d6a2ed8f2310f970fc;
wire [MAX_SUM_WDTH_L-1:0]        I2c72248cbe49ec0a0febac2437b8a6dc;
reg                              I67d57e38df8cb35ca686ac2eb44e233e;
wire [MAX_SUM_WDTH_L-1:0]        I964e17c41a134c080e9c43412a514f3f;
reg                              I23955b54e486f0f0d21a2809a9472b86;
wire [MAX_SUM_WDTH_L-1:0]        I94f1724740defe5bb7e40041d0e266a0;
reg                              I1e11f0088959aa40b4ad1a047b59caf4;
wire [MAX_SUM_WDTH_L-1:0]        Ic19486b6ab0373b9c0ad8f7597782d8f;
reg                              I68c35d63dc95baff41b4dc27a86d2342;
wire [MAX_SUM_WDTH_L-1:0]        I31243de90dc2a1656ca9d5e03bdd78da;
reg                              I837183265ee22d080e81fea468ab0887;
wire [MAX_SUM_WDTH_L-1:0]        I242a30bdc8699d8ff550b25dd53d6c59;
reg                              I413b1c1985a6c9c6f202e85ff901e3a8;
wire [MAX_SUM_WDTH_L-1:0]        I9d15f76bb68b214057566cba4b511214;
reg                              Ic32c6734132776c290155a80025fe366;
wire [MAX_SUM_WDTH_L-1:0]        I9cc16a00912e7dfc05fb505a9db23cd8;
reg                              I624958486d181501c7a8ec2642cb503c;
wire [MAX_SUM_WDTH_L-1:0]        Iacf9640cbf486411d6ceb8fe1a2fd5c9;
reg                              I04864c28351edb33b61a103add6fb875;
wire [MAX_SUM_WDTH_L-1:0]        I9015033ab0caf3fa41dae4de43f24a82;
reg                              Ida3dd5e990ce3c237e9628a9a090901e;
wire [MAX_SUM_WDTH_L-1:0]        Ia630e59cbce82a570ae3890a6c0221e5;
reg                              Id182a776b03f48fb139c28194ae7ab6b;
wire [MAX_SUM_WDTH_L-1:0]        I4904ab14b19fa1b6befc218bc7be3842;
reg                              I0c5539373b3868d0664a92157b4b4226;
wire [MAX_SUM_WDTH_L-1:0]        I282d2eb4e74e034694e33273b9cb19d5;
reg                              Ic0191941cb968bbd7644c21767423d2e;
wire [MAX_SUM_WDTH_L-1:0]        I3f33901c407a87e10d86c13c83dd52eb;
reg                              I163cf58b9a308e0439a8dc7c1526e6b5;
wire [MAX_SUM_WDTH_L-1:0]        I43f41bf07836cee48069e9890c1de2a0;
reg                              Ie08ad9bd71329858c1742c8f571a1c36;
wire [MAX_SUM_WDTH_L-1:0]        Id88480a0a350bb5fcf01ed5fff0bbd4c;
reg                              I3c10d579f80bd0106506ad047d75f188;
wire [MAX_SUM_WDTH_L-1:0]        I1d9b9ff357667a362f0442f19986f451;
reg                              Ieca2767ac27170058499d83016447aa7;
wire [MAX_SUM_WDTH_L-1:0]        Ice73589836da9028def6efb24a04dbbd;
reg                              Ib9c194ec16f435a9357cb344cf25bdcc;
wire [MAX_SUM_WDTH_L-1:0]        Idb72c046c5996fbbd80b706666ffbd92;
reg                              Ic920452d5997a8477724fa78c86c0fba;
wire [MAX_SUM_WDTH_L-1:0]        Ie5757e7b1647ab7d43cdbcf98cbb77fc;
reg                              I6eea5fde8e2517554ad6ba25018572dc;
wire [MAX_SUM_WDTH_L-1:0]        I6072331f838d82329a07a4ffa340c7b6;
reg                              I9ad2f6fd2d7f68011fc926ec9abd5c34;
wire [MAX_SUM_WDTH_L-1:0]        Idf6875955525d80dc660ce956f4a84e7;
reg                              Ied33f18cbb778d5ba744d249f91c950b;
wire [MAX_SUM_WDTH_L-1:0]        Ia96955d9c0a8a587e0afab37c8415d8c;
reg                              Ibabf61085ca7af8dfc7927b3656a76f7;
wire [MAX_SUM_WDTH_L-1:0]        Ifec374bce7f5507438f550df22d61a01;
reg                              Iddc5b5b4501f9f13bcaf22081e5a70f4;
wire [MAX_SUM_WDTH_L-1:0]        Ief67e897e57b96e2ec200e82bbc7caeb;
reg                              I67f87fbb746dd937fffc534c596f36c4;
wire [MAX_SUM_WDTH_L-1:0]        Ide604e9bbe35cb55892a4602e18b2527;
reg                              I45bdd0cfe107da0d57cad1333bf95e3b;
wire [MAX_SUM_WDTH_L-1:0]        I262f2390e77ec486ccd3a6ed05816e2d;
reg                              I4d54dd2ee2f32909098d3cc2b6689220;
wire [MAX_SUM_WDTH_L-1:0]        I280e20c20c0b4f26278b3de9b2ff84e4;
reg                              I7bfb4c5d9e22d1bd8811844d9c74dff8;
wire [MAX_SUM_WDTH_L-1:0]        Ib3a0307176d424a4733720416d71069d;
reg                              Ib9d58222da98f29fa302b4896594fe26;
wire [MAX_SUM_WDTH_L-1:0]        I76060709de3ea188748849f043c59ac0;
reg                              Iea3e35ece9fdb3aff3b9ff5369e9a7e0;
wire [MAX_SUM_WDTH_L-1:0]        I8be20605d26d218911e80a883a90d085;
reg                              Ic44eab478be232721e7a43d14beca32f;
wire [MAX_SUM_WDTH_L-1:0]        Ieafa9d74d4a61d28ac4a913db460bf33;
reg                              Ifab075b1437495268b6a3be4cb022e71;
wire [MAX_SUM_WDTH_L-1:0]        I6fd1b4395af175eff85b3bfeef4c329b;
reg                              I2919272e9ae3996a3e1d602ff72ba86d;
wire [MAX_SUM_WDTH_L-1:0]        I39e6d3fb468aa40ea73535e81556ea65;
reg                              Ib6fbe376477afa58bfcc17a8564f78b2;
wire [MAX_SUM_WDTH_L-1:0]        Iae449b74e50e0907feae9e60f2329426;
reg                              I659322a9fd0d5eac514437b02e0491b3;
wire [MAX_SUM_WDTH_L-1:0]        Iebf769a6bdaf214c1006c55c608d4eda;
reg                              Ic68f500938d80460ffdb33a0adc48298;
wire [MAX_SUM_WDTH_L-1:0]        Ia030c08757123aae947f86ab8bfb6d94;
reg                              If5ae6fbf843fdeee17945bc5ce81aec8;
wire [MAX_SUM_WDTH_L-1:0]        I8c35c5b343b552c22000e194c517ca12;
reg                              I94460b6ce7b776bcc5eca149eab80c26;
wire [MAX_SUM_WDTH_L-1:0]        Ibf80bb564263ea85bd886a8617f09bb2;
reg                              I3347717ba9556e69de30ce7533d4f5a4;
wire [MAX_SUM_WDTH_L-1:0]        Ib8dfd9b8badef282ca00a4f793c3c868;
reg                              I2db290170ddae8dc52ce07edaf48b365;
wire [MAX_SUM_WDTH_L-1:0]        I596ad7e132f272cb196b74faa8c75aa4;
reg                              Idd775d9fe6fa8dbdbfb07d4071b9caa5;
wire [MAX_SUM_WDTH_L-1:0]        Idc629414f6d0236ce0714cfaae23f065;
reg                              I6cbc06919b9c695d99621db6f8d768cb;
wire [MAX_SUM_WDTH_L-1:0]        I157fdf8775206858c08682db3039b084;
reg                              I5b8a1e1a6b904b0f6822c224ee0486e3;
wire [MAX_SUM_WDTH_L-1:0]        Iacbb4daf5ce5c7eb1a2afe30d0cb5382;
reg                              I3f5053e519a928640ae49cf4e5b39d1e;
wire [MAX_SUM_WDTH_L-1:0]        I4e08021c0235fafb60200aab97827a8f;
reg                              I7c965c047d862c973d09a81abe03a845;
wire [MAX_SUM_WDTH_L-1:0]        I730634ea15ac94d241f3ad2d6393a227;
reg                              I9b8023f4dced915cd52c91bc9d4ed78f;
wire [MAX_SUM_WDTH_L-1:0]        Iee367c535d9c39f872d2ec043e7e7b33;
reg                              Idc6b6357741c9887a9db1037ccc2d922;
wire [MAX_SUM_WDTH_L-1:0]        I68bb1f26f878862f288c1f57049cf58b;
reg                              Ibe97860165dc5d9a076ebd935385ae51;
wire [MAX_SUM_WDTH_L-1:0]        Ia9b5d9ede006c56a6d83905529c77b7b;
reg                              I777ee54ff20d0544af18ad8a870d6915;
wire [MAX_SUM_WDTH_L-1:0]        I1487170cb1f3370ad45efc801cefc8ab;
reg                              Id18c5a1d4eaa73a94e699e5f9e3c3d35;
wire [MAX_SUM_WDTH_L-1:0]        Id88568dd34fbee42c9cb8cc15ac5c31d;
reg                              I72939e49bf2d9c6a84e404419fc644a1;
wire [MAX_SUM_WDTH_L-1:0]        Ia30539545e66c4cfc16828140149180a;
reg                              I57b7b48f13436b19a8d6a47e014eb41f;
wire [MAX_SUM_WDTH_L-1:0]        Icbfbb37bad6344005dd233b3605a784f;
reg                              Ia3ef2f70c5abaa852586a33c505aee0d;
wire [MAX_SUM_WDTH_L-1:0]        I91a6408a11fab36a8ba3dbd3f895a803;
reg                              I6d423a7d17e05a3c597ec6ef6c5a7cba;
wire [MAX_SUM_WDTH_L-1:0]        I47b878f27c30f79a37e97e022307e9e9;
reg                              I48e3309c61918c3991852b45d9c72ea5;
wire [MAX_SUM_WDTH_L-1:0]        Ie76b0739aec66f8860870e66e87a6445;
reg                              I472352e7027b9df2fa957d9fd68443ff;
wire [MAX_SUM_WDTH_L-1:0]        I50383e3d7c172eedfa00aa50a9faac4c;
reg                              Idbbf2ce4a30787c5f07c3b908a73da75;
wire [MAX_SUM_WDTH_L-1:0]        Ifeaa99e03bda8ded058f98387de3d49d;
reg                              Ibc9a860879ccc58c815b9f6caa23320a;
wire [MAX_SUM_WDTH_L-1:0]        I4255ac1af4367c321567c4e46b06ab25;
reg                              Ia71cf07b645c58cffe33be1a9a960eb2;
wire [MAX_SUM_WDTH_L-1:0]        Ia445bdc7def7d8c1eec31ab892c25c41;
reg                              I0ceb14ac0187d804f9692e0c55b8e941;
wire [MAX_SUM_WDTH_L-1:0]        Ic3b4752136ac08e343933ccc3a4ec47c;
reg                              Ief18a19d451f05f6051e3cc8de16d73c;
wire [MAX_SUM_WDTH_L-1:0]        Ica6707efd6d44ba6bbb87c0593a3d828;
reg                              I30be0b18e4415ca50f2d8149efaaafe6;
wire [MAX_SUM_WDTH_L-1:0]        I739267bcc50c54b8a685cb3c6afc5cc1;
reg                              I7ec15b73b2811b44e1e50c74a9f921e9;
wire [MAX_SUM_WDTH_L-1:0]        I9160d11439c5140c0109b5190eb82e6b;
reg                              I0fd2f706e374a4eb57ee26ab50201e15;
wire [MAX_SUM_WDTH_L-1:0]        I6ff7b86cd7f63f9243646f1be10b2577;
reg                              I44f170d02bae7fe044456e125a98451d;
wire [MAX_SUM_WDTH_L-1:0]        I165653ab165cfafe2b74cd441331f9e1;
reg                              I30c0fcd89e0cc7c5fa348df7b4fa2ccf;
wire [MAX_SUM_WDTH_L-1:0]        I08a8cd6965c23af6650568b654831b20;
reg                              I13a98f98c54b2e412cd88c96f016c41b;
wire [MAX_SUM_WDTH_L-1:0]        I9b6a674dbcbfcf65f1ae0deb8fc3566d;
reg                              I9890f7fc708c7b8cf460849b4a30025b;
wire [MAX_SUM_WDTH_L-1:0]        Ie3a336de822ac7baf8486b1618ef1126;
reg                              I5e69e930a318dcb0594a823b3129d650;
wire [MAX_SUM_WDTH_L-1:0]        I5fc3c26d6c5aa893dfd5caa0f677233a;
reg                              I403303228c0df825f67436f4a7e64061;
wire [MAX_SUM_WDTH_L-1:0]        Ie22b94121b58f17af14c75bfb27f96dd;
reg                              I946246be5b4745508b7d4b578f83aaa2;
wire [MAX_SUM_WDTH_L-1:0]        I0d9f8c99194d9d6e187b4ad02fcce8b4;
reg                              I95f0acd4f955058041c035789c3a4d99;
wire [MAX_SUM_WDTH_L-1:0]        I71e101962e766a4d1484b3235359a4b5;
reg                              I4082b3564c1949a19ed35bd5a88e1ef4;
wire [MAX_SUM_WDTH_L-1:0]        If2539da6722562bbf31786fd0036666a;
reg                              Ia7606050c683ecefc510ba92ac539a9c;
wire [MAX_SUM_WDTH_L-1:0]        I22c8ccd4a9018ad1c129aa058bf579d8;
reg                              I5446c1c323774715371c73bd1be66697;
wire [MAX_SUM_WDTH_L-1:0]        I83330fef69470d2f5def8e6d7d9c50d2;
reg                              I3a8e9e7d2cd6751e8500a5567cef5acc;
wire [MAX_SUM_WDTH_L-1:0]        I0539d598bbe3d50940329a282c801328;
reg                              I621b20d29d3a9a9f41065bc3c3bbd2d8;
wire [MAX_SUM_WDTH_L-1:0]        I202f88fdc946494d55fc8831c2e8a34c;
reg                              I263aad78110a1136eb7012c6983b2a8d;
wire [MAX_SUM_WDTH_L-1:0]        I3ee10f6a7785a236db317515fdd23a2d;
reg                              If4308ed204e33952c9931f8fe257aca4;
wire [MAX_SUM_WDTH_L-1:0]        I453fdf4fbb5af5bd28a20d7643da9eb2;
reg                              Iddcfab4a7022e0f12fd20cb34e9b9d02;
wire [MAX_SUM_WDTH_L-1:0]        Ic4a6c02880a9aead7353332708e3f388;
reg                              I759409e242eaeb144a53e630a8cfd514;
wire [MAX_SUM_WDTH_L-1:0]        I7fb3b66cb48521f8715f66bf5642cdb2;
reg                              I5f96a68d20e3ebc71dad4b43305baa20;
wire [MAX_SUM_WDTH_L-1:0]        I2fd872df07f50688486c0d602cfc5549;
reg                              I5d92fdff96b9cd64f3af2b28b13e9956;
wire [MAX_SUM_WDTH_L-1:0]        Iccefa45795486757515d95e5908b306a;
reg                              Iab2f643f81921ed8464e1bbd9fa8c68e;
wire [MAX_SUM_WDTH_L-1:0]        Ib1357cb20f471f1670ac2448f964f8eb;
reg                              I17d7f36fdade16dbcf621fe302bd7e57;
wire [MAX_SUM_WDTH_L-1:0]        Iab953a8974a1eb619dc0f074c003b5f9;
reg                              I23afd747ecece714e32fbb896b5c022a;
wire [MAX_SUM_WDTH_L-1:0]        I6e37582849c2c98fd15ad92d22c222da;
reg                              I388528eaf83566cc56b23485a9c05962;
wire [MAX_SUM_WDTH_L-1:0]        If004de0cac6e5f7701a1fce48c6936d5;
reg                              Iea424dd9d8916c4951b8746408b8a521;
wire [MAX_SUM_WDTH_L-1:0]        Ic1efa395cc1fd2c5a1d1559fb169a5a0;
reg                              I73bbf90b625d56f663ad10f9d21d8e76;
wire [MAX_SUM_WDTH_L-1:0]        I8e96c69e7d872be23229353808c34953;
reg                              I41796b587316c600bf583edc62649bd8;
wire [MAX_SUM_WDTH_L-1:0]        Ib6aded6c73a8cc3cb964b0ae895b859e;
reg                              I7009c18515dd43d8dd2e5d1ee6779641;
wire [MAX_SUM_WDTH_L-1:0]        I939368b76d98b43826c68c7f468a5632;
reg                              I797c9cb725f88c07be28f017871d17f8;
wire [MAX_SUM_WDTH_L-1:0]        I544f6263f16cd5e0b7cf28c511a8f6e3;
reg                              I06b48093d4c9b0327c3efc6fa4ca7daf;
wire [MAX_SUM_WDTH_L-1:0]        I484545c4d2c869d79eb17f51e11070a3;
reg                              I04c734eb876aa722e84d6b9edd297978;
wire [MAX_SUM_WDTH_L-1:0]        I39289e6385a9bc378a9b8dd440249a7f;
reg                              Ifb89e7ad8ef661959d82b7c22f187243;
wire [MAX_SUM_WDTH_L-1:0]        Ie9cce5746a83479a567bbaeac6dbf497;
reg                              Id1dce2b9eafc35fa71df33ada4aac539;
wire [MAX_SUM_WDTH_L-1:0]        Ic044d7419cc43736d278c2df33b4a3cc;
reg                              Ied19cb51636bfb029ba8a2c390f97105;
wire [MAX_SUM_WDTH_L-1:0]        I6714551e8885ef5e4490673fe1b2dad1;
reg                              Ie46b71f55aef4d00168202431d47dce0;
wire [MAX_SUM_WDTH_L-1:0]        Ie9ab3c88ac62369e3d92d110165a94a8;
reg                              I8c0c1a0a35f4f7a688f516c567242d39;
wire [MAX_SUM_WDTH_L-1:0]        If38feb4f76f761dce6145731ad235d7f;
reg                              I53222c82827cab7c770e057ae91bc10e;
wire [MAX_SUM_WDTH_L-1:0]        I6359856a1843d8c8b65dc478bccb3acd;
reg                              I8015717cd36aabbf2cf4aa3a5c234690;
wire [MAX_SUM_WDTH_L-1:0]        If6f3d91c3c7a43622b9a522492cd83d3;
reg                              Ic0c13c9a929c8c46e8702cef74de8955;
wire [MAX_SUM_WDTH_L-1:0]        Id023a6298e65da1f4da3831f5136afc2;
reg                              I71d7f72d83b7410de31e09ea96adb95c;
wire [MAX_SUM_WDTH_L-1:0]        I6b24690f394792edb0d82b3b9e110851;
reg                              I1db4ea6916125702e7fb09d0f742e60a;
wire [MAX_SUM_WDTH_L-1:0]        I5b55c285f7e3e78447fee68532ab9f7f;
reg                              Idc445d3f5b3b62562b0ac83e5f17e92a;
wire [MAX_SUM_WDTH_L-1:0]        I32701d9e4b96853c53f0ab651a6a4ba2;
reg                              Iee6e52d75c093a24eb4e5e0b45feb256;
wire [MAX_SUM_WDTH_L-1:0]        I82f266e5792cdb6e7ebd264e246161f5;
reg                              Id48fe0672aa98f987162931527e9f9bc;
wire [MAX_SUM_WDTH_L-1:0]        Ibfacfe5b83819afe7fbd4bffa2d6d4e2;
reg                              Idce46f6d03376bea1ba361e8c59f8bd1;
wire [MAX_SUM_WDTH_L-1:0]        Ib8e68a77ad8b9e7cf415bee17645c3f9;
reg                              Ie79ce8adeef2c3c24a3386f054d0cf5b;
wire [MAX_SUM_WDTH_L-1:0]        I644ee0055a55f54ab3544bb532e39c61;
reg                              I0d41bef808860bde56d48792764612d5;
wire [MAX_SUM_WDTH_L-1:0]        Ic5467e42aa377c6ffd8f70673808774f;
reg                              Ib6ae81df8db1dae269437861ee11ec0d;
wire [MAX_SUM_WDTH_L-1:0]        Ic57eb4a034247a4c952d8224ea9f2bac;
reg                              I33ddee677715877c11a1df45cbfb01ac;
wire [MAX_SUM_WDTH_L-1:0]        Ia642db613c0ec1ca4e69afde7a14a839;
reg                              I433dd5092cf1851cd196feade3cfa6d8;
wire [MAX_SUM_WDTH_L-1:0]        I432aa7cb844286c442356954f8814260;
reg                              I71d3a999d88e591e102398409b3adebf;
wire [MAX_SUM_WDTH_L-1:0]        If520c1cd27f9d4bc52d0d029f693b660;
reg                              Iebecd2d19f9174d87deedc1a273e7baa;
wire [MAX_SUM_WDTH_L-1:0]        Ie87075ac979410cc11099a356966b8a2;
reg                              I168afc1863f909dbcb6a9230db9f3e00;
wire [MAX_SUM_WDTH_L-1:0]        I6fab46b1766878b26b53f352fee98223;
reg                              I1c4b29e48d0effac4839037ae5688334;
wire [MAX_SUM_WDTH_L-1:0]        Ieaf14683f40374c4531326d228cb43c3;
reg                              I431fc2e9533012c8571d8158d4777dea;
wire [MAX_SUM_WDTH_L-1:0]        I5149125aaaad943d891df6a3c2be93a0;
reg                              Ief72606c77113ae37845e4aa4a2ae5e7;
wire [MAX_SUM_WDTH_L-1:0]        I770dff588ee1f52f58bea1921cb23383;
reg                              I641539560711ff1824bd90baa0f21f96;
wire [MAX_SUM_WDTH_L-1:0]        I8f0a90e761111a613d2488285534a500;
reg                              I3ac0799861144b599995318bdade2114;
wire [MAX_SUM_WDTH_L-1:0]        I765a8825e42180a6c63f7b33703bb483;
reg                              Ie83fa8157a7cce44c2e25f46ce897dbb;
wire [MAX_SUM_WDTH_L-1:0]        I512cc8f6519aa08aee18225b56d47c9f;
reg                              I8be4711146486fea913843e497065b50;
wire [MAX_SUM_WDTH_L-1:0]        If08370fd0e8af818c6db20f43e74034d;
reg                              I65171c9ee8449407484e5c82d13c6751;
wire [MAX_SUM_WDTH_L-1:0]        I0ff382edfc8051459657ffa3899f5f73;
reg                              I7353ebf3a1cde89d2bb3fa667f7f5485;
wire [MAX_SUM_WDTH_L-1:0]        I9d2864024148337277523ef7fa2e1600;
reg                              I669d34b955d2991ebbb31c149ad1b6f8;
wire [MAX_SUM_WDTH_L-1:0]        I1c85a2d1df6749a194072eb731506bfe;
reg                              Iabb01dc9980b4879a7356712b51df0d6;
wire [MAX_SUM_WDTH_L-1:0]        I3e3ce8b4ead150a6eae2e5c701c7b598;
reg                              I373841aa2bcbad8232d54ac9035a3ef9;
wire [MAX_SUM_WDTH_L-1:0]        I45bc13ae0e0554a79c62cd9c6aa8f2a5;
reg                              Ib6124faff821158c6a2c9a9c454ab68c;
wire [MAX_SUM_WDTH_L-1:0]        I92678f5b52c9c55556ff7f17f0f607b7;
reg                              I6f7a45fe64ffeda9ed120be3a4519aea;
wire [MAX_SUM_WDTH_L-1:0]        Ib4bdc9069d0c08655f5e87f705943eda;
reg                              Id1dafb7e45b860d506e0c2c91b28142e;
wire [MAX_SUM_WDTH_L-1:0]        Idbf9094c94c931f16fba468b9dd59a25;
reg                              I5f1609647f1e71cef4ba2d605c6c8445;
wire [MAX_SUM_WDTH_L-1:0]        I1c3c4ce44610e04c5eef2fcbc2ea5114;
reg                              If17c0096ce34b88007247bf4c429d5c4;
wire [MAX_SUM_WDTH_L-1:0]        Ie84be0ae8311d906eff08f7f5b214943;
reg                              Ifc2963762403a00c4f3662b2863c991e;
wire [MAX_SUM_WDTH_L-1:0]        Ic90b98708faa8c8b75d4bd9a52c292f7;
reg                              I5fdd8e1550feaecd81b82069fe73ed7e;
wire [MAX_SUM_WDTH_L-1:0]        I8eba6f14f42701d22859fbea94bd1871;
reg                              I85654bd3a07b4329aba17d8b27777f4e;
wire [MAX_SUM_WDTH_L-1:0]        I6d83efa9f988328f487e9232bf2633a2;
reg                              Ibf2a253afde05c905d0b2404c5a808a0;
wire [MAX_SUM_WDTH_L-1:0]        Ic23e01562c8a753fd70c343297be288a;
reg                              I3ade5535a79ce83857481ac771cd8618;
wire [MAX_SUM_WDTH_L-1:0]        I5669856f88f5e2c98f64df696db76414;
reg                              I221524a69e18854f029cad30e8f94e8a;
wire [MAX_SUM_WDTH_L-1:0]        Ic3a608b850709286ea0ad2f67425d9ac;
reg                              Ied764ee7730ad129b6f62837ef50774a;
wire [MAX_SUM_WDTH_L-1:0]        I5267fa34449e6eebe891017fc32d0749;
reg                              Ic98f33c6a4613534bcc9b6bc4b4f2d17;
wire [MAX_SUM_WDTH_L-1:0]        I599d01cfe6e54d8e45d64446c446818d;
reg                              I92eb6f60c14ee9eecb01718b01ea980f;
wire [MAX_SUM_WDTH_L-1:0]        I8f94dbafaac589ac9f14b56d4556ff96;
reg                              I97e82e5f6775d1e31537b891597223bd;
wire [MAX_SUM_WDTH_L-1:0]        I754563caea429d3d0e22df5d193b84eb;
reg                              Iba1c0ebd9cefeb0dd7f690bdbbbfec58;
wire [MAX_SUM_WDTH_L-1:0]        If7f373506cac70f8ba1222db135c27e8;
reg                              I235c3a9fd3e8ea1cee762c10bc8e2c53;
wire [MAX_SUM_WDTH_L-1:0]        I69f563e7b7ad483893ac9c4684349769;
reg                              Idd474d80b50992537d6f527faf279800;
wire [MAX_SUM_WDTH_L-1:0]        Ia0a02781c674fe5d769206448d475245;
reg                              I88a89b2d938552458dab9bc34728959b;
wire [MAX_SUM_WDTH_L-1:0]        I1b7a401bc11741e6f011fb9895b5c797;
reg                              Ib105151d91678f81978495ff94b1e651;
wire [MAX_SUM_WDTH_L-1:0]        Ieb528d666fdb708279184bb59eac25d9;
reg                              I4edd64d1f1da865b1eb886e22726a033;
wire [MAX_SUM_WDTH_L-1:0]        Ic3ff7ce12c836bf0693252b9a7a7cfe8;
reg                              Ia7c9c24f8e993526e76c6915e56908c4;
wire [MAX_SUM_WDTH_L-1:0]        I19bba6a58ad3ef959b33701f82761984;
reg                              Ib0dadebad37d9ea9d01350054872863c;
wire [MAX_SUM_WDTH_L-1:0]        I8acc93b34974c1e708b0e1591f7b2d3d;
reg                              I76fd9005abd511c3c5bf6c77de8bf2f3;
wire [MAX_SUM_WDTH_L-1:0]        Ib60d4ac0fcadcdfce5a14fb92f58423f;
reg                              Ic124975d36a292816146a2fe61ab3ab9;
wire [MAX_SUM_WDTH_L-1:0]        I039f05d5be891a37e04556f1eae674d2;
reg                              I70a4926e9e6a05fa9ee51a26988862fe;
wire [MAX_SUM_WDTH_L-1:0]        Id0f75e19b94541ed5c5c352d13390d2d;
reg                              Idc5e98f6958786ccf95d39b922b42ea9;
wire [MAX_SUM_WDTH_L-1:0]        Ife1190f76c2e251704c2960c23330a48;
reg                              I8879df010bbdf6e5fc9370e2fb3289b4;
wire [MAX_SUM_WDTH_L-1:0]        Id3e0c98bff2636e216b4d3a0ffd51054;
reg                              I94a9de743d5bedbea3876de954f479bd;
wire [MAX_SUM_WDTH_L-1:0]        If4d3b31b87c0f723241d35ce7e854eba;
reg                              I17c9d8f658dd6b2916b645d103f4702a;
wire [MAX_SUM_WDTH_L-1:0]        I72369dedfe36cb22269033cc305b730c;
reg                              I384e50fa8daa639124f083dda56fac00;
wire [MAX_SUM_WDTH_L-1:0]        Iec71fe7fcebccf1ae0d10a5d187fcc44;
reg                              Ie165d0729542c81ca89f45d15e0afd3d;
wire [MAX_SUM_WDTH_L-1:0]        Ie11da10808c4ca84f399535df6261307;
reg                              Ie8e29053f122a9247b0dec291c6ef4f3;
wire [MAX_SUM_WDTH_L-1:0]        I280fa9d114e227cd649bf0e55e845651;
reg                              I453dd7d7c0a2f003f0b67e909630d641;
wire [MAX_SUM_WDTH_L-1:0]        I94c4e11670b4233fa072517a8f19c901;
reg                              I5707d30ca29842b6a96cfaeb44ac6668;
wire [MAX_SUM_WDTH_L-1:0]        I4dca2dd40a7127ce44f83b430a34c738;
reg                              I3fbd40faa4c3b78b547b8348c466fd1f;
wire [MAX_SUM_WDTH_L-1:0]        I1a24e98165afa62bd14986911a36fb6e;
reg                              I9a403c511fe2d44472ab319a9477199c;
wire [MAX_SUM_WDTH_L-1:0]        Ife1164cad7cda4aa9a08d94dfe86add6;
reg                              I9db50007841762c9a10f6b7e9d40f858;
wire [MAX_SUM_WDTH_L-1:0]        I8d8d95ff26f33f69a182b32ccde23905;
reg                              I89c5af1a6176cefa1f77ee69996473cb;
wire [MAX_SUM_WDTH_L-1:0]        I2508854bcbab37bd09c9465c377c06aa;
reg                              I5ede62333e0f7ddc5446b653ba9a2382;
wire [MAX_SUM_WDTH_L-1:0]        I140078292f7209eccacd53a8bab18016;
reg                              I69d82ab774d52c219509e993e7cc4deb;
wire [MAX_SUM_WDTH_L-1:0]        I141fb1cbe09f9abe282cffd4de815d25;
reg                              I0eaa22f5eca8f33dd254fe241017a098;
wire [MAX_SUM_WDTH_L-1:0]        If79d1d378f7c6fd29fc3335ec5f5c51d;
reg                              I570c036d0237c53bb069c52d621e539e;
wire [MAX_SUM_WDTH_L-1:0]        I4a41999cea9357a85c73a0af509eeac9;
reg                              I9d7614d286377329eb3999213889b707;
wire [MAX_SUM_WDTH_L-1:0]        I8e517c401d62dbb10dcc96ab536f6afb;
reg                              I3eab1582cc42db0ac7739386cce2a712;
wire [MAX_SUM_WDTH_L-1:0]        I8ad3627f171eadcc960a688ac0afcbc0;
reg                              Ie4827dc0983c1a63053c08de6e36d375;
wire [MAX_SUM_WDTH_L-1:0]        I85c4d3d6c8408c6f38741257ed177ca6;
reg                              I2eed3d32a27d51036e17c4a21382b4c1;
wire [MAX_SUM_WDTH_L-1:0]        Id66c47fd69c175a4393e975a269cf053;
reg                              Ie039ab562e9cf90289047b5425186123;
wire [MAX_SUM_WDTH_L-1:0]        I37dca40506d61bdeab1255ed4892ca20;
reg                              Iefbdf686d9452a62cb99cf023a4d9fe7;
wire [MAX_SUM_WDTH_L-1:0]        I340c98b886123c541a1b8d9fc8a6d48c;
reg                              Idc5dd6caa4ed17a63746d30d381a944e;
wire [MAX_SUM_WDTH_L-1:0]        I2dc64c3b06588542b027f997437bee63;
reg                              I17086dc5193aa55e5c6f56ecd365cc00;
wire [MAX_SUM_WDTH_L-1:0]        Id92a37c091100e9df08e24498ecb4022;
reg                              Ib2fe0f68044c11f879e512a200f8099e;
wire [MAX_SUM_WDTH_L-1:0]        I74a4b9365391fd20c34588002ad40547;
reg                              I768720af835b02a8dab376ef23d17a15;
wire [MAX_SUM_WDTH_L-1:0]        I461195b7ae78743e09ee50486ad6ebe5;
reg                              I1d98943b01a6a2d8c4db18b98dd62f5c;
wire [MAX_SUM_WDTH_L-1:0]        I356d747600182675699a2d2634d4c5ce;
reg                              Id3b089fb6edd5bcfdbca142fddd5ff89;
wire [MAX_SUM_WDTH_L-1:0]        I87d6a5d30c3e4202cf51f33c7a770c51;
reg                              I5196382b75d16892d550f17893de15ec;
wire [MAX_SUM_WDTH_L-1:0]        I960768a84aec9d5b8bc7c1c523024a25;
reg                              I6387919f2426c283e2d70e471cda54a6;
wire [MAX_SUM_WDTH_L-1:0]        I09b5273bb15d48a7fd78559930fa6d1c;
reg                              I3b84dad6d0dd8730312b3e20c6d5a2a8;
wire [MAX_SUM_WDTH_L-1:0]        I5814a85c45fd0f7be21ed325235fe4b7;
reg                              I2a4bbedf880a9a7b4e1bf946f9f96c0e;
wire [MAX_SUM_WDTH_L-1:0]        Ib06b60cf9933dd8952206c5f3ccced8e;
reg                              I49d35ec6369de10afb15be8e0cf135c3;
wire [MAX_SUM_WDTH_L-1:0]        I67347c413b5efd8ff9e0d5bc7ab2a047;
reg                              Ic3ba4531855366e9a060cec1c7694844;
wire [MAX_SUM_WDTH_L-1:0]        I72b1bb104bf2843f161448baf7aab44b;
reg                              I4dbabfd592b74aef93b819163130ef5e;
wire [MAX_SUM_WDTH_L-1:0]        Ib23d889edb5a6d9f27de977d3b1a2616;
reg                              I9ece87047aec25abc02a5eea72f0e647;
wire [MAX_SUM_WDTH_L-1:0]        Ifaff9dd032cf96487be819c59b03000a;
reg                              I3ed6426fbdba8aaf1c948cca7442b3a6;
wire [MAX_SUM_WDTH_L-1:0]        I028ce03be0618b816e0ecdf43d4cd6e6;
reg                              I24075f37c6bbd90c83370de1a2e58af2;
wire [MAX_SUM_WDTH_L-1:0]        I6ae2523095237282533e0b5f1c26b488;
reg                              I3175159add7b814df637c2db8feb43f6;
wire [MAX_SUM_WDTH_L-1:0]        I5aba6218461e8d571be03a3ef041ebaa;
reg                              I0a569f6536789efb7ad2377c11842830;
wire [MAX_SUM_WDTH_L-1:0]        I6ca8a1fa2c72b1c61d11dc7d1ba5f37b;
reg                              Iae6ed7748692f2edf1aa9d73380075f0;
wire [MAX_SUM_WDTH_L-1:0]        I3ec5819176ad4b0895a9118d90ab22b5;
reg                              Ib4ae1cedd09d72c235765a6cd7e91366;
wire [MAX_SUM_WDTH_L-1:0]        I49b64469d298012dbb131d879bff38d6;
reg                              Ie2d946edaddd3c87f328e861f3e72c0a;
wire [MAX_SUM_WDTH_L-1:0]        I95361d5f524ccb9feb42811af5c482e2;
reg                              Id6b508145cd21ba088ab8fda34577c35;
wire [MAX_SUM_WDTH_L-1:0]        I9c4b34b5fb1d59c132bcaeb6258675df;
reg                              Ifa6e3541f5e12bf9677ffc51d0392749;
wire [MAX_SUM_WDTH_L-1:0]        I613d4b1e3b9e812b785c9cf14fefdfe6;
reg                              I21e72a7e5870151c3247d15121e5fb4f;
wire [MAX_SUM_WDTH_L-1:0]        I848ed394bd4f0b199d11c0ff458394a7;
reg                              Iba283e99a57d0a3b78ad2e309c316b65;
wire [MAX_SUM_WDTH_L-1:0]        Ie65a0634454381e24bb3223a333e3ad0;
reg                              Ifba3e46933049cb093d2c1809f3a8a3e;
wire [MAX_SUM_WDTH_L-1:0]        Iad166146f7df5e8068fc6efe4d3e4141;
reg                              I4af3e2bf2ebc913ac902b48da672c5b6;
wire [MAX_SUM_WDTH_L-1:0]        I63e45abd4d27219bddcef06108b72021;
reg                              Ifbadefd3a7ab50719a703400ddd742c6;
wire [MAX_SUM_WDTH_L-1:0]        Id1bacd13718f7c29c26b63c239d04dd8;
reg                              If2042aede3390bd208a281f0380c95a4;
wire [MAX_SUM_WDTH_L-1:0]        Ia3104c69fb4f7abfb5efa3874169a7ad;
reg                              I19b73c5c93a71e90f620572f23f0e6d2;
wire [MAX_SUM_WDTH_L-1:0]        Ie1b7257c99831ec5864f65958ecf14fb;
reg                              I4b99891bed4f5c149cd4a5b4f1dde0f0;
wire [MAX_SUM_WDTH_L-1:0]        I4accbad1b451ed2b622e15ef9ae16d13;
reg                              I3472ee8c06644490252e606b62bf9bd5;
wire [MAX_SUM_WDTH_L-1:0]        I5ce8b2f633011e89356243a1a71edeb6;
reg                              Idb1efe99b5d7fd567a7f82cfd52f7eb8;
wire [MAX_SUM_WDTH_L-1:0]        I3e5139f24e3d082eb31b0e61ea9fa1aa;
reg                              I24f82a3f2c0e8df486fe495dd95cf8bc;
wire [MAX_SUM_WDTH_L-1:0]        I61cc8a0f49e393721a62a776e4793deb;
reg                              I83ecf12f3b38fc14c3b75e47b71ecc09;
wire [MAX_SUM_WDTH_L-1:0]        Ie631e40caade823a196370fc3358f042;
reg                              I74cbc0ec3bb682e0f927890eef8d7a58;
wire [MAX_SUM_WDTH_L-1:0]        I4c971e714427664c59c6371e14781bae;
reg                              I989dda9add29306d7b3c0f376822763a;
wire [MAX_SUM_WDTH_L-1:0]        I36ca732e811d67cd742d24fd4cae887b;
reg                              Ibc929201e2eeb3e61cc8f0acbade497a;
wire [MAX_SUM_WDTH_L-1:0]        I354fdd241d5d07f0d8380fe8924e0a8c;
reg                              Ib0dfbbbca2d3d264065f73b4241caed5;
wire [MAX_SUM_WDTH_L-1:0]        Id38b705f5d2863a020a475ffffc8afd6;
reg                              I339786aa60d4c71d12c65db27ac420fe;
wire [MAX_SUM_WDTH_L-1:0]        Id6e5d67e7bb7c4b999459374ea80459a;
reg                              I3ade020bbdf8f954821f737439513043;
wire [MAX_SUM_WDTH_L-1:0]        I05341013abd4206eb66fcddfd63bfe26;
reg                              Ia50526cd3a3174bebc5a7a0889fda661;
wire [MAX_SUM_WDTH_L-1:0]        I15da71a21f5842cb65b543d9bc3e267b;
reg                              Ie9f37dba0791359bc426a73639ce33ad;
wire [MAX_SUM_WDTH_L-1:0]        Iccf255fb3422c558465e45226068a16d;
reg                              I9518532a8617fc8290eb6a5e981dea94;
wire [MAX_SUM_WDTH_L-1:0]        I1c2674b2e6b269ed539827412c5199a5;
reg                              If66524125bfde5aa48ac70c4e448b38f;
wire [MAX_SUM_WDTH_L-1:0]        I6a3f405bb4a0c4448d9b9d3dd95d036c;
reg                              Ic3ec6375998b05a3e48f6c5fe7b3910b;
wire [MAX_SUM_WDTH_L-1:0]        Ib528bb7a64cce4f694081d151fa6fa86;
reg                              I0ac421af6e311b6005c3e02e93ff94ce;
wire [MAX_SUM_WDTH_L-1:0]        Iaa40bd3abf668a21e0f87c7bda7b3f69;
reg                              Ib9db80f43718305a8a8774d8d80c86c9;
wire [MAX_SUM_WDTH_L-1:0]        I919d36a7f6ad42c4bbc23222beb73106;
reg                              I3b775b06b5d78fcd7373c966a62f44ad;
wire [MAX_SUM_WDTH_L-1:0]        I648d2a279dd1f587b1e45eeb35f2fa90;
reg                              If2372a5956f21f97eeb9c76281b6675e;
wire [MAX_SUM_WDTH_L-1:0]        I194a64bef92ecf6714141eaa5d41c9d4;
reg                              I7b32c2b108e24750e2a24785668af3ea;
wire [MAX_SUM_WDTH_L-1:0]        Id332e7f482524adeac7f7cdafcf5ca46;
reg                              I8ec99197a7d823f5745d382c10161430;
wire [MAX_SUM_WDTH_L-1:0]        I226383d68f89db716cfd8d08b837865a;
reg                              Ib895fec0b3756932b85962c1d129a03e;
wire [MAX_SUM_WDTH_L-1:0]        I2bdf5d319ba9089a4da34b108f5c5ae5;
reg                              I76aab345d13c6678fe37a4a7133cfd7d;
wire [MAX_SUM_WDTH_L-1:0]        Ia91800792941ec7cc60415c3f844e4ed;
reg                              Ib4f368fa3d3ec11d9ffb2ae9a2ae6310;
wire [MAX_SUM_WDTH_L-1:0]        Id7c507d96098ee7a955af8a48ee5d72a;
reg                              Idd0f3cfc5599481c954a2bfe69f044e5;
wire [MAX_SUM_WDTH_L-1:0]        Ie15e4c1bcdb0e18085d4b320ac6a925c;
reg                              Ie624c4dad5036a25ca314b94cf3c4b95;
wire [MAX_SUM_WDTH_L-1:0]        I5485d9edcafc6202f6e5f0969979802f;
reg                              Ibf4b3caa5655cfb6663f9b7e2383bbbf;
wire [MAX_SUM_WDTH_L-1:0]        I7fe364f9f537cbef782e7007848a1c10;
reg                              I049d1c09c15def12ba7bae95fc1c3d55;
wire [MAX_SUM_WDTH_L-1:0]        I52dcf5bace9cadcf8a895aaa6a8c1da8;
reg                              Ide06ba186ddb179b489ba6e3e209e3e8;
wire [MAX_SUM_WDTH_L-1:0]        I13a9eec6175e695ab8bc4516cf57d6ec;
reg                              I1b78785ebe2e7f77a3125a6334c4dc54;
wire [MAX_SUM_WDTH_L-1:0]        Iee73a7c685a4cee03f33d3ef379b1c8a;
reg                              Ie79c93f1703121713fb9401617f349a8;
wire [MAX_SUM_WDTH_L-1:0]        I740dc91716e3906ad078e2c7cc3c925a;
reg                              Icf25f076eec2bf81c899c66f6cfbebc0;
wire [MAX_SUM_WDTH_L-1:0]        I514d2dc697e9b39ba027c418a6df6cb9;
reg                              Ic5c837a0556d1cb66edbf0294d08283a;
wire [MAX_SUM_WDTH_L-1:0]        I782726e317a2aada9e755bcbc4b0d3fa;
reg                              I51ff4bda38746682e3cd4c68118c3216;
wire [MAX_SUM_WDTH_L-1:0]        I11eb26cf0f0b3a334e8f7317bf8d9eb0;
reg                              I1c074a53e6c0f2467bcdd7c952f51670;
wire [MAX_SUM_WDTH_L-1:0]        I26cb63ba20245b2c332b09e25c4409aa;
reg                              I37c49c5a2af240496f5a5706b0d42ea6;
wire [MAX_SUM_WDTH_L-1:0]        Idd7691d31f8d0c09ee988116d574ec59;
reg                              Ia94c439131e1df5c95fc8ad3cfdba473;
wire [MAX_SUM_WDTH_L-1:0]        Iecc02842a2d2b9b9e8187f2d39e62e05;
reg                              I723a6fee3b2496f23c48b3584f8bf9ce;
wire [MAX_SUM_WDTH_L-1:0]        I5551342f1751fc64f32744a46b9649be;
reg                              I648b62fa0bc2185c1756ee531e8e34de;
wire [MAX_SUM_WDTH_L-1:0]        Iff7c29299f005c1cd5a16b64601e727e;
reg                              Ife631f9a3c4c64a3d92aa9586ae75f3c;
wire [MAX_SUM_WDTH_L-1:0]        I17a5446e942bcc1dc2c96930e0a87a70;
reg                              Iaac1d82f0846fce1bd88ebf8e60300ac;
wire [MAX_SUM_WDTH_L-1:0]        I719b67f84e07e90dfd29a8cd5d94cf39;
reg                              I48cd09f035f668536cd288a23010b07b;
wire [MAX_SUM_WDTH_L-1:0]        I2c835dfb3596b8bf057a7cc21122c81f;
reg                              I119b2e5c2fea5338244c4019884af26f;
wire [MAX_SUM_WDTH_L-1:0]        Ib71b3d357c98dcdfae5c777ca3082275;
reg                              I2bd34b2fd12f12bc301fd0d5d69c0fb6;
wire [MAX_SUM_WDTH_L-1:0]        I086bf19f620c8a8f6888e775cb1ed7f4;
reg                              Ib715b1e0061b84ce614a30d961a83e7e;
wire [MAX_SUM_WDTH_L-1:0]        I802c554d5b04af6b949677819a4966ed;
reg                              Ief8c2838abac83370fd7ec25c06d509b;
wire [MAX_SUM_WDTH_L-1:0]        Iceefb06cb3715e1b41e6f7d89420e5ba;
reg                              I561d79eb079915c0b1732cbddb119c2d;
wire [MAX_SUM_WDTH_L-1:0]        I56948bc48c0220893d68004615a6ebaa;
reg                              I8bb75bf828d5ef337fa6a965808e4638;
wire [MAX_SUM_WDTH_L-1:0]        Iec1368f034655d61354ab5b5e94d7d89;
reg                              I11ba339c8250d07b497c88a39a6df1ac;
wire [MAX_SUM_WDTH_L-1:0]        I1e43c0aeeb8a2461d208eba24967af30;
reg                              I173aa69cf52114e223ac1410d90b4bfe;
wire [MAX_SUM_WDTH_L-1:0]        Ia6eb85b127cf9c1a437611556296b967;
reg                              Ia4e89e99acb95f4183474b94798ca35d;
wire [MAX_SUM_WDTH_L-1:0]        Ieba89aa901e61218074af53a2484a74b;
reg                              If4c36727ab1c29bf78f72e8acfc00d7c;
wire [MAX_SUM_WDTH_L-1:0]        I8b3b875c6c07bd97ba598a5139156fa4;
reg                              I6426943b4ab66f17c2b7b399ccc7a6a9;
wire [MAX_SUM_WDTH_L-1:0]        I7b33ddad346077928620344542b9481e;
reg                              Iddcffa815489773b3688fd68dba18bd8;
wire [MAX_SUM_WDTH_L-1:0]        I11d967a5c5d14c88b5587d4cfed1d05f;
reg                              Id00642563679fa9a6696f8e7bbdf6576;
wire [MAX_SUM_WDTH_L-1:0]        I27458d76b3ac6520fb379405c6b2956f;
reg                              Ifda1c55899cd3506853cc82b450b3936;
wire [MAX_SUM_WDTH_L-1:0]        I2525111a2fb5f10d64bbd16e148653b8;
reg                              Ib5d1a7cdbcba0b654c12063d4f1768e1;
wire [MAX_SUM_WDTH_L-1:0]        I7b7cbcd1c6d2a2eeaaff474536a69eed;
reg                              I5e8ed024e2f2548bb375a2ecf1918a5f;
wire [MAX_SUM_WDTH_L-1:0]        Id2a7f0781d18dccc7c4e0b383b7cddfa;
reg                              Id25deba967318f049de8163e67262f4b;
wire [MAX_SUM_WDTH_L-1:0]        If8bc141d98ebe1be7fa81cde5c65868e;
reg                              I925f6b549a25cdc8f85152eb21ea3b58;
wire [MAX_SUM_WDTH_L-1:0]        I8645e1326c66f5efef4b9c923599d1a3;
reg                              I9b49e1acb81ef5b088b808d2e4ce9954;
wire [MAX_SUM_WDTH_L-1:0]        I0426ef66185128dd1ef4dbb68dcda585;
reg                              I6386a4dd26e7c36165dc265b3a2c93cf;
wire [MAX_SUM_WDTH_L-1:0]        Iddd954df5bae9b4240e0512f746669a9;
reg                              Ia20709f08cfff3a51d4af1e81d640400;
wire [MAX_SUM_WDTH_L-1:0]        I29e940970d87e8e09b26ab1b0b8f2286;
reg                              I1ff042bdb52aac5d69791e96e2f9706c;
wire [MAX_SUM_WDTH_L-1:0]        I488f6d9676aa85a55d030bf12e8997a7;
reg                              Iaa2cbf59f6f61198b4fcf5a741cd5bc8;
wire [MAX_SUM_WDTH_L-1:0]        I99d761b75ade1fb2e8afbb1a77752609;
reg                              I01c94743a11042e75638ba6618356203;
wire [MAX_SUM_WDTH_L-1:0]        Iac4e3d20178049f9c59abf374752dccc;
reg                              I0a0340a0e52145f3597accfe4a4e8624;
wire [MAX_SUM_WDTH_L-1:0]        I618d33f26badabfa578908903a613bce;
reg                              I3bb4d24caaa0882a75125e466070f0b1;
wire [MAX_SUM_WDTH_L-1:0]        I822d7973afe090b2764335f1b72dfd0e;
reg                              I44ead0ab5ccc53226fccc03024643771;
wire [MAX_SUM_WDTH_L-1:0]        I12c1035353e553b3b6a13bb174ce6020;
reg                              Iaded125f7fd5c833e7206dd7071069be;
wire [MAX_SUM_WDTH_L-1:0]        Ia6d61947d36fc128c689808c82db80f6;
reg                              I373be7c3f9511a2906584e33e5048abf;
wire [MAX_SUM_WDTH_L-1:0]        Ie9b042f686381739b9ff219041f1e0ce;
reg                              Ie0b5f51835ebdb508a596eeebf0e4847;
wire [MAX_SUM_WDTH_L-1:0]        I0c4268c01aed70ce4fc71531bf4bb862;
reg                              Iddb75e0197b9a76b36a59ac2a7ccdf3a;
wire [MAX_SUM_WDTH_L-1:0]        Ia34e42f8de91fa4861b0c6cac5dcfc29;
reg                              I08c03198b9599b2f4590e3022e398f7c;
wire [MAX_SUM_WDTH_L-1:0]        Ib7c5850b4f7cc77be2048d114a2128d9;
reg                              Ia4f3cff223e24815ee1d86bf41756f06;
wire [MAX_SUM_WDTH_L-1:0]        I32bb50faa2b246b2d3b462a79be597c5;
reg                              I56592e1452c4b559af19465b30230ec0;
wire [MAX_SUM_WDTH_L-1:0]        Idc6d40a49f05c5422758cee50f787eb1;
reg                              I213ce488e5345fa405a9c5df297d6f74;
wire [MAX_SUM_WDTH_L-1:0]        Ide1d7dc22a4b271ef764df14ac22366a;
reg                              Iefac1e428116a797c2c0803410ac5601;
wire [MAX_SUM_WDTH_L-1:0]        I7ace6778ac86b3e05939a3fcc716136f;
reg                              I8b419d5827e5b1af9649d602401c189a;
wire [MAX_SUM_WDTH_L-1:0]        I044e01e8d2df46e03f00a0af2beb0bf5;
reg                              Ie989550c9101de382056dd60d5da0e01;
wire [MAX_SUM_WDTH_L-1:0]        I45a7ddcda2662e36b7617dfe64514346;
reg                              I259010e323e1e8dcd9dd719091131f6c;
wire [MAX_SUM_WDTH_L-1:0]        Idada779a1ac7b844867571d77054b657;
reg                              I389ac86954fd70464c9550e3fed4ed33;
wire [MAX_SUM_WDTH_L-1:0]        Ieeba01b18a244ab8c0ac263c138fabcc;
reg                              I77371f0e55b4684d1af196ed52d3d997;
wire [MAX_SUM_WDTH_L-1:0]        Ie4c9797a955778694dd8615219cb51e7;
reg                              I5a21996f5724a2a49fcf8e928c01b062;
wire [MAX_SUM_WDTH_L-1:0]        I28a5ed4c239e64c76bb6e566b50cfd23;
reg                              Id46108963921efa50aff64d4dd7d1701;
wire [MAX_SUM_WDTH_L-1:0]        I79a705ee1e414fe4a5fb14e9b3ce9597;
reg                              I8da50e5093acefb6f809aed64564a53e;
wire [MAX_SUM_WDTH_L-1:0]        I04f90a907f10a7fa1ae3591b48094d5c;
reg                              I03b0694777d0160a83cbc82ac1397736;
wire [MAX_SUM_WDTH_L-1:0]        I31d25b1b49e65216e90b39aa27acd6be;
reg                              I85c2bffb93569d9fe1b1bcb10b98bcac;
wire [MAX_SUM_WDTH_L-1:0]        I1f6540c5f037d861dee2c0091cba01ec;
reg                              Id00274c88b93867a80606343add1cdab;
wire [MAX_SUM_WDTH_L-1:0]        I9632bb500b7faaaaeb649d74c21cbe8c;
reg                              I61e829cbf7d6c0ef8ddc11677981e2cf;
wire [MAX_SUM_WDTH_L-1:0]        Idd0217a35c3adc8abc7bb581a5df7a2d;
reg                              I9e8ae2aed048068b01b3bd46f30baae8;
wire [MAX_SUM_WDTH_L-1:0]        Ic05b46168884322644db4e331d37d759;
reg                              I7dab71adbe62687846fc027d2789451d;
wire [MAX_SUM_WDTH_L-1:0]        I53c88dc237bb2cd02d50fd7f0a168a48;
reg                              If1295608bd218ed60922a0b95bf1d098;
wire [MAX_SUM_WDTH_L-1:0]        I7450d4ab3ef0227e93a02bfd620d047b;
reg                              Idf04e08c120ed116af14a62659675b44;
wire [MAX_SUM_WDTH_L-1:0]        I2b16e5b4e279bb29c3c675b72083e5fe;
reg                              Ieb7614ad1b1bfed3e2b0089a72fe214a;
wire [MAX_SUM_WDTH_L-1:0]        I70c92e8ada46476d15ef4b3c620d2601;
reg                              I589062eca318b25dfe5735da455b6fe1;
wire [MAX_SUM_WDTH_L-1:0]        Ib193b07804d6d5f111b06bda487bfa5f;
reg                              If3db87afb3ea184c9e4020c5e45cb161;
wire [MAX_SUM_WDTH_L-1:0]        I885433b0ab16c6d87abe45af13c9e529;
reg                              Ia14bc1fcd5bbdcb60b8e68298f7d716a;
wire [MAX_SUM_WDTH_L-1:0]        I198c055930cb89d0390c336eda8fed4f;
reg                              I268b60cb371b3d46dc3f8b0009f541b1;
wire [MAX_SUM_WDTH_L-1:0]        I688a2c72e69b217d2673e8da75146a83;
reg                              If2cd93b57cd1c2b91ee7a73a97dd19f2;
wire [MAX_SUM_WDTH_L-1:0]        I3b6fde4ed14cd68af1468ae1d4cc1a22;
reg                              Id81305359a07db527e49fda05cd2784f;
wire [MAX_SUM_WDTH_L-1:0]        I5d3df1e7563630311f56143ee6d97a8e;
reg                              Id8292eca087c1a17dc8b5a572a76f21f;
wire [MAX_SUM_WDTH_L-1:0]        I90a7ea789d3bf7f9126c786474a56da0;
reg                              Iddb19725b093506e5e521d8d68dcb8e1;
wire [MAX_SUM_WDTH_L-1:0]        I5029424c9d9fe923eeb858b1e62cd758;
reg                              I0b573d3a86a3111451da661e46384876;
wire [MAX_SUM_WDTH_L-1:0]        I1e805c70d50c2765b4a03ad2982dc421;
reg                              I0ff479e61d1a0cede88ebffb073c60be;
wire [MAX_SUM_WDTH_L-1:0]        Iba58175a7fd5c5da650222193caff0b3;
reg                              Icd6f8f5df6b4ca4c81855e974db76526;
wire [MAX_SUM_WDTH_L-1:0]        I7401a0501ba69c5559fbf00c77e58dc5;
reg                              I7ce064a756dad56d37684d5d7d168047;
wire [MAX_SUM_WDTH_L-1:0]        Idd9f7ea657ea9cdcb45a7e4b573b9d50;
reg                              Ied2ea62cfb21602645babc36e27b8218;
wire [MAX_SUM_WDTH_L-1:0]        I53f275395dd6be17961a5edc3e8da7f2;
reg                              I79b85da6e5ce0b02ebd1619115c98e24;
wire [MAX_SUM_WDTH_L-1:0]        Icab010d78cd66b02e089c74f04bf4e75;
reg                              I8e1ddd7e4185c28caa71d30bc28138f3;
wire [MAX_SUM_WDTH_L-1:0]        I376a48b7e0195a5aacc76a0ad8bd14b2;
reg                              Iab0bff1633e2f3ea0bfbc291f3ab5d29;
wire [MAX_SUM_WDTH_L-1:0]        I241622b0367dde514f96ece55c8c3964;
reg                              I5f0751fceaa008feba5c6867ced453dc;
wire [MAX_SUM_WDTH_L-1:0]        If94a1abfb972f63629d07e64dc23863c;
reg                              I9f6751c15237c20b0cf2175575195ea7;
wire [MAX_SUM_WDTH_L-1:0]        I07b9b1f4fa01b16cc69356057d3b6154;
reg                              I6ea50be10bc990a1206cdc9e28e0c4c2;
wire [MAX_SUM_WDTH_L-1:0]        I2288a6ad3b748b716249f4adc42d52c4;
reg                              I43c2fab87f70ea883321ab82de85f133;
wire [MAX_SUM_WDTH_L-1:0]        I022df337bcc05ac5648b8ae2e42f3a76;
reg                              I1af02ed6cf00d4cb0704b5e44c83bfa3;
wire [MAX_SUM_WDTH_L-1:0]        I60d9a7f95fb8623753002ecaf9a4efcc;
reg                              Ib71611afdd0381cc1884f5ddbbae1acc;
wire [MAX_SUM_WDTH_L-1:0]        I23a74ea5e7174d95e6d16a5e85ac236b;
reg                              I38fc49afce0298846ae8ed63ae715e81;
wire [MAX_SUM_WDTH_L-1:0]        Ie697d28d757df82b3901564bda43251c;
reg                              Iddc3e44d83e8253e5129b6cbf5082df7;
wire [MAX_SUM_WDTH_L-1:0]        I8572aedc94f7243ce5eacb332c81eae2;
reg                              I975a87bdda30c5b6be8d2f0e4b107450;
wire [MAX_SUM_WDTH_L-1:0]        I6734123aaf6320da75638b212812732f;
reg                              I582bd96afa764ded148202f738b7a1df;
wire [MAX_SUM_WDTH_L-1:0]        I7f6dc6f0f403c58f9aaaa70c2383a666;
reg                              I6fb88d97bc9ed37a06b729020a1df140;
wire [MAX_SUM_WDTH_L-1:0]        I66391978843c39b6acbdb4847a01050a;
reg                              I1500943c4a550e78fc169437b0a663b7;
wire [MAX_SUM_WDTH_L-1:0]        I4f756e4125c8af5c412944b273e01cb0;
reg                              I0b83f4ef8ba9badb27e81b32765ec5b6;
wire [MAX_SUM_WDTH_L-1:0]        Id2c9f7ac95de07148c54803f69347f56;
reg                              I2c420acf428e44cdd9ca9998e276f258;
wire [MAX_SUM_WDTH_L-1:0]        I5061e13a179d27e1ba5f89ce8ee0fd4a;
reg                              Ic7b6dae3017b55dd3cd27423d5f1b0ec;
wire [MAX_SUM_WDTH_L-1:0]        I0f7c32fc1548fb49b8041f55c157498a;
reg                              I4a91a7c9b2a0f3552b8f2ef4e2398be2;
wire [MAX_SUM_WDTH_L-1:0]        I89ffab735ee30423c82e079ed98216c5;
reg                              I99ff29c7ba68b5d0819f1e1bead51287;
wire [MAX_SUM_WDTH_L-1:0]        I9494921d8487ee0b314f75cf0380fd2f;
reg                              If06b00be0356a2be5074d958ddcdb2f9;
wire [MAX_SUM_WDTH_L-1:0]        If2b3e7d1541cbd8ffc2b4cfc3ad13a57;
reg                              I604283449f13c7b225ea03f99f2e296a;
wire [MAX_SUM_WDTH_L-1:0]        Idf3d79da44f2d686f5bd43c3c1427430;
reg                              I2b600e5f5c146ee97c4044c08e1f5ad5;
wire [MAX_SUM_WDTH_L-1:0]        If8125ad3c9e7f0a2b84106064d320996;
reg                              I9fe16403fc21bb1159a5e0305fd1ef69;
wire [MAX_SUM_WDTH_L-1:0]        Ic9018b88fa91fb638bbab0613795ae13;
reg                              Iabdb9374e5caee281c25b003624b2c4e;
wire [MAX_SUM_WDTH_L-1:0]        Iad4ea0196eb32f9a152c9e6fe5059e46;
reg                              Ibd12036702fe60b57354b3aac921559d;
wire [MAX_SUM_WDTH_L-1:0]        Ia8ff29ed728e7f2ae4213f00328b495d;
reg                              Ib1639811de6eb1c38257800c201fb704;
wire [MAX_SUM_WDTH_L-1:0]        I70717726200ec02929f679ef05496455;
reg                              If926d98f659e8fe4bbf36ad2c5c852c5;
wire [MAX_SUM_WDTH_L-1:0]        Iaf1e4c7dae6ad89567836877c08f57d2;
reg                              I211f8d7f97ebb8eb3e50313513abfb1b;
wire [MAX_SUM_WDTH_L-1:0]        Icd09aa81e9b43528af73e23b2f0f80cb;
reg                              I304ac9f96945546cdf1b6f1fa7136731;
wire [MAX_SUM_WDTH_L-1:0]        I6ebb2b94f0f80425f8401ae823d92a1d;
reg                              I7a9800418bd5c195fc47a72370680b56;
wire [MAX_SUM_WDTH_L-1:0]        I4a2c3204a6a9936d4a215b46c0ffd045;
reg                              I5f6a61c9f0c67510e148e596f553a4d6;
wire [MAX_SUM_WDTH_L-1:0]        Ib02c0694762c4815448b2c8d3df767c2;
reg                              I8e313ceb21359bcc44114ab217b1c394;
wire [MAX_SUM_WDTH_L-1:0]        I98cee6efbbe565d3a4de16703189782f;
reg                              I4c9518755c33d725221ad79ee6badba9;
wire [MAX_SUM_WDTH_L-1:0]        Ibf981c01a9d44cbea3c6d8ead92bc2ab;
reg                              I3c3cffec9f47c9979cb9503f222f370c;
wire [MAX_SUM_WDTH_L-1:0]        I864c33e8ea204d20a9baef4584f22d4e;
reg                              I68d6769541fdc3df321e192f645c667f;
wire [MAX_SUM_WDTH_L-1:0]        I6ad3228e0e2e1f19648d73e83ba5a229;
reg                              Ided55428cbb77f454c2607ac783d7548;
wire [MAX_SUM_WDTH_L-1:0]        Ie099210a99a4899c53baf39559592690;
reg                              Ifd3d4f3e2a388b3c70e7704d6351e0ba;
wire [MAX_SUM_WDTH_L-1:0]        Ieeec71d9df4613555fade2ced7b3baf1;
reg                              I17d32f292758416fe02527dfd938fa0d;
wire [MAX_SUM_WDTH_L-1:0]        I4931884e3544af182bcda9061091a42d;
reg                              I9ce3942aba354c1fd7d6b9a39c994d7b;
wire [MAX_SUM_WDTH_L-1:0]        Ib3fb10da528d450251764a9b9ede0dba;
reg                              I2c6c6041c9c69c84f4d64af6458955f5;
wire [MAX_SUM_WDTH_L-1:0]        Icdc9e676957b2223d60c413331fa982f;
reg                              I830a4fffe1244e071eb82c28ddc4a308;
wire [MAX_SUM_WDTH_L-1:0]        I381f6051282c062ccf53866830344cd4;
reg                              Ifad8e46fc3844bbfaf434a14f6b5869d;
wire [MAX_SUM_WDTH_L-1:0]        Icfc21935c007fbbceb2a67ebe1a68a0b;
reg                              I10a6c6a8fdb0003de1f360c148777d0f;
wire [MAX_SUM_WDTH_L-1:0]        I120d597a80158374726e064fb0f099fb;
reg                              I4cde586fc28f8d03fc9934d56f7ff7b8;
wire [MAX_SUM_WDTH_L-1:0]        I2520aa556aadf851f58f0b1820498730;
reg                              Ib83a067fb08e118dcf794902beef9405;
wire [MAX_SUM_WDTH_L-1:0]        I6203f49a08107f7185ebadeecf2c16b0;
reg                              I358cf9609272a4562423a85f9b2f56bf;
wire [MAX_SUM_WDTH_L-1:0]        Ia706fb593b63cebbee0321c154cb859b;
reg                              Ic1e9d9113150ad57954c0e369259dc62;
wire [MAX_SUM_WDTH_L-1:0]        Ia4b5f2b07556629673fc6576bc49a5dc;
reg                              If7fe3f5ccbb5b279e41fd183c8ff3974;
wire [MAX_SUM_WDTH_L-1:0]        Ic532c6b85b156f821e0742f47239a65c;

wire                             I40a85f3ef46def30cd7707afd2c7fa44;
reg   [MAX_SUM_WDTH_L-1:0]       I18d11d94a39d5d7687736d266d3e1902;
reg                              Ib64114b4af6a37b3d52bd38cb83459ee;
wire                             Ib8963a4ab143aba7fadc61d89f937f4e;
reg   [MAX_SUM_WDTH_L-1:0]       I6b9ffa985ece553b83f7227e7a85141b;
reg                              I06ed412c4554e98837146a5c7a6c4789;
wire                             I9565de7442acee8455d1c4f8ab43ab07;
reg   [MAX_SUM_WDTH_L-1:0]       I49fdba80df1c667dd264e5105a530332;
reg                              Iefa11849e46b6ccd923e622fdb878315;
wire                             I26b11eb80b9a1752998f7ab1379e4124;
reg   [MAX_SUM_WDTH_L-1:0]       Ibf4fc04c9e0aa536a8e4b8a6192d8498;
reg                              Ia4245ce0efa56b1234283f4969246280;
wire                             Ibb068f313ff784191769e8da44f023e1;
reg   [MAX_SUM_WDTH_L-1:0]       I899abb7dcba235ff2afb410a87e16973;
reg                              I671b766473f67c92b75716e2bd9a9596;
wire                             I2348d423bff186f1841ecaaf44f4f2c6;
reg   [MAX_SUM_WDTH_L-1:0]       Iab322f0da75316ca9937802a327dd537;
reg                              I24b5cce7252356b606027b301ac6bf48;
wire                             I3b28138cac28625778c34d4bb1a4aa55;
reg   [MAX_SUM_WDTH_L-1:0]       Iba0a4530bce787d70253a92c123f589e;
reg                              I2f0d19d012f0bd45308356fce1a50049;
wire                             I8928563d2510725797f96917767f9bae;
reg   [MAX_SUM_WDTH_L-1:0]       I4475d6a1e59d35444a6a2d9647c6761a;
reg                              I939c483ddfc18ee8dca73a1c98e6ec4d;
wire                             I989726d5ee5f23a016e85b0945573f05;
reg   [MAX_SUM_WDTH_L-1:0]       I217e2e1eb3404ba9ff06d284a18256b6;
reg                              Ife63de208f77b322e1c885e78790f997;
wire                             If88711683bd32856ce45937b841581e3;
reg   [MAX_SUM_WDTH_L-1:0]       I2003418e663144ee49f1ed044f6a0062;
reg                              Ia065f925c78015a3736219a5c7129439;
wire                             I015cf78df7e3417d5296eb0ad3019674;
reg   [MAX_SUM_WDTH_L-1:0]       I4496255218b6d0f5374328803aeeb412;
reg                              Ie02e0e9e2627b178d6c54ea743b3993b;
wire                             I31908b38609b532f9f142a97e0442e55;
reg   [MAX_SUM_WDTH_L-1:0]       Iecbb3f290db6dad3393b592ca946fa13;
reg                              Ib1e432e0b2d7979227d2cc591ed8e383;
wire                             Ib98eadb333ebca2f58c40b8f93d87250;
reg   [MAX_SUM_WDTH_L-1:0]       I9f88e23f2a17035b31840356a5d0bfde;
reg                              Ib05aef46725afee38240d81738c673f1;
wire                             I4a0f0579aa9b7af7b516780074ca6560;
reg   [MAX_SUM_WDTH_L-1:0]       I3fd4a13843fc09ca68b827a8b09e6c49;
reg                              Ie7bea07eac0dc36dbce430e6dd088b5e;
wire                             Iaebca9b574d490aeab28fbbfb1e8fd9a;
reg   [MAX_SUM_WDTH_L-1:0]       I1530e79da3803bb87787397f19822dbb;
reg                              I3f42e9b5ae0fc5c9315670cad33374ce;
wire                             I3ad613d80a126f03fb9125fe6da1bc8d;
reg   [MAX_SUM_WDTH_L-1:0]       I613821692bb99a8a6739d3c3ab7211ac;
reg                              Ie6f54d5d349ba8e19295a9ce17ba3f35;
wire                             Ic116b21b5744ec42a9f41eff3ddd1707;
reg   [MAX_SUM_WDTH_L-1:0]       I5ac600834d567934bd2f0b14a3c38ab9;
reg                              Iab7ce2d8e89a5862f98bd812751d1d17;
wire                             Id9f7e6885737ee2d3128081915a685b0;
reg   [MAX_SUM_WDTH_L-1:0]       I84fe1a1ecad408b16557957b01cc94b9;
reg                              I8a4157cd8206e66109f979bd9bde53b6;
wire                             Iad36872fbd9ac694d47cc0491f3d021e;
reg   [MAX_SUM_WDTH_L-1:0]       I7d03cdddc264c89446cd80405c34d69a;
reg                              I5f0937deee06e2177807a6d0fbc2e2b0;
wire                             I0794dcad0f96cf58fda60c561a1144fe;
reg   [MAX_SUM_WDTH_L-1:0]       I5cf7e3cb90e84c3ac6a66fb6dde220af;
reg                              I598fa274e3ada377f2e7a43d7dfd9231;
wire                             I8b4cdd738b1ed431764d4a51be668460;
reg   [MAX_SUM_WDTH_L-1:0]       I602c2e5bfa93cb3c87af70dd69b0375d;
reg                              I4a3da449219c7068a0bfd3a192d2ead1;
wire                             I79e67c70ee26ab7623355ec5042dcb28;
reg   [MAX_SUM_WDTH_L-1:0]       Id50fe525d660f0bb0ac3bbe6e68758f1;
reg                              Ia7a0522cea2126afdae3fb9f123d51fb;
wire                             Ie0a573c73ca9198012dc8ff4f8373973;
reg   [MAX_SUM_WDTH_L-1:0]       I6a68067b177340dbea2c53f7d8bd5f14;
reg                              I5d901ed468b60a31e199d12612a0b396;
wire                             I6a4cd5680e34df5ccfea4a7eb72113ec;
reg   [MAX_SUM_WDTH_L-1:0]       I9efdcdeee8883d30159881f8831a2c03;
reg                              Iceced38b8b522d1679ed4e1cad38c282;
wire                             I9885460698fe454e65fea4a6022e5df0;
reg   [MAX_SUM_WDTH_L-1:0]       I46290d63552b8cac8d22358cb38c5887;
reg                              I7d3d6075ca3828a533b52dc3cac3a652;
wire                             Iee7e507956faf7cd903ac2dd636b7819;
reg   [MAX_SUM_WDTH_L-1:0]       I6435c7b1b3bfc5dae42cb1b3b03aefc5;
reg                              I0869d337e6cce62a05b29c5baa4ed436;
wire                             Icece56258c1ffa7a0257d68ef9ff5ee7;
reg   [MAX_SUM_WDTH_L-1:0]       I63b2f1c2148e595a40bb41968e4b9a65;
reg                              I36ae963a57878d2c5b647910e003dea0;
wire                             I6c15ea618986f2043f402959ac23fb1b;
reg   [MAX_SUM_WDTH_L-1:0]       Iafb6296c59c2dd241c880c6d57352617;
reg                              I5851ca9a7e932378c2bdf2c118b498dd;
wire                             Ic45cade04982e60abe32a359999a778d;
reg   [MAX_SUM_WDTH_L-1:0]       I0b982beca6221db7b3ec2afb3833a60e;
reg                              Ia5597b68eb3f1c1d371cda63fa1fe034;
wire                             I670dbb51097dde1f56eeb7e25ac50369;
reg   [MAX_SUM_WDTH_L-1:0]       Iece8968796771c1ef094808823da8962;
reg                              Icc939d3c403d238cf5c9c196cac91886;
wire                             Ia3fb4901b185e64ccb788dcc1d7cfb1b;
reg   [MAX_SUM_WDTH_L-1:0]       I05c7cb4a076239b8976a76d418ad6149;
reg                              I0bd90c7dbb94917bb46a3e008484f582;
wire                             I15a23e6922630f6d409706b1c4100d22;
reg   [MAX_SUM_WDTH_L-1:0]       I9076162e7b10bffbc9473e35b407e986;
reg                              I6ec7620a49b53a8377767e363e88d471;
wire                             I08eb91ffc153d5007de61e2938407d18;
reg   [MAX_SUM_WDTH_L-1:0]       If702042844ed38f5e7103382ef4263eb;
reg                              Ie512ccdcaff0cc5c29277e28f1ba5fa8;
wire                             I642d63513e039da95a66c1cd4336f84f;
reg   [MAX_SUM_WDTH_L-1:0]       Ide63b2762649761944db237c8efe69ae;
reg                              Ia115f92bd6dcb4167f0771941a18ad59;
wire                             I1e35f6f8ac9e61787a3b263e5e4ac62c;
reg   [MAX_SUM_WDTH_L-1:0]       I1cec628c6d6e22895a0f0c0258851171;
reg                              I7c8174a3579ed90c0ec89941ac53e287;
wire                             I5af04bd644d9c14f56884acd1f6674a7;
reg   [MAX_SUM_WDTH_L-1:0]       I46b0b74552e89df91c0027f0f093e1f5;
reg                              I7d6b68dbc5ac773ce97df3a6726c6836;
wire                             Ia9bc04087c3926bdf993858e683dc3f6;
reg   [MAX_SUM_WDTH_L-1:0]       I68dbff67a1910346ddc0281b445f4439;
reg                              I5045f1311d1e891577f3f8a09078fe79;
wire                             Ia8c23f2c6c80bc389fd66aee524975cf;
reg   [MAX_SUM_WDTH_L-1:0]       Ia42f547c0b02c2de66f2ff383ca1741b;
reg                              I105c3326421f25d3b9931e2178c794d4;
wire                             I74ff51ab0824be97bf311b50b4ce5401;
reg   [MAX_SUM_WDTH_L-1:0]       If456045711d535cea07d9dd5ef9b04c6;
reg                              I838c5c183e758ef4f28ad86d16befd87;
wire                             I22cf21c1e88c0b8ff5d5b43835b1f61f;
reg   [MAX_SUM_WDTH_L-1:0]       I9585ff28ce0f3bca71d582b1cb8937d7;
reg                              I33c782b29a89c2ec375038b88919b564;
wire                             I2fc87e59765765e16bae0761ab5741ec;
reg   [MAX_SUM_WDTH_L-1:0]       Iac3dfb28a343cbb391fdf58684e091ef;
reg                              Ia21ec0ad85852d1eea449283d1d45a7c;
wire                             I6c6297e7aca3c7d8a9f8c3542f8b070c;
reg   [MAX_SUM_WDTH_L-1:0]       I82650d4bf0a9b51e245665259f40fe60;
reg                              Iae32e0aebc2719c3e476a5300f1bfdea;
wire                             Ifbc2ba75815cb3aece1d327a5c15dba4;
reg   [MAX_SUM_WDTH_L-1:0]       Ib21e67aa9696222891a0b33c414b1bbd;
reg                              I6914a92b8da6d6db6f2e8806c7efc5aa;
wire                             Ib1bba2d65c2224f05a444c6170aba187;
reg   [MAX_SUM_WDTH_L-1:0]       I1e168bf1a0dd18ff31d3560be00095f1;
reg                              I60cad827424e4799360141222a80ac57;
wire                             Id75ce45a6df04b3d173b288b52d82138;
reg   [MAX_SUM_WDTH_L-1:0]       I97e6d2bc8c1ad455f7c61de81e8d4826;
reg                              Ie3389948b5dd781ac9087e62cf93dd2d;
wire                             Icd148cb7a25bc30aafd0271e00356527;
reg   [MAX_SUM_WDTH_L-1:0]       Ie1170db51d408ccc7360ce53c94a9644;
reg                              I566475d003c9fc40aebaba87655a0668;
wire                             I80e8b0fdd6bfadac9c8a788bd9be4b97;
reg   [MAX_SUM_WDTH_L-1:0]       If58c2c1e1dffe04295f3313595ffe319;
reg                              Idb2467b1104f5b924d419208f2573df4;
wire                             I471dd2bc897a40a9463f4984952d4fa6;
reg   [MAX_SUM_WDTH_L-1:0]       I9a9fb4da9fdf5bd42cef32c7d8fa65d9;
reg                              Ie0a8d219223bc68ea3040cbbd349caac;
wire                             Ic61bade7088606659ef8568dc134f686;
reg   [MAX_SUM_WDTH_L-1:0]       I785e4a1f2556289db0bd024e429bbd3e;
reg                              Ide01b9dcf3a3019d689d79f4d7ce0f32;
wire                             I298e98803772a458fbeed1de632c0555;
reg   [MAX_SUM_WDTH_L-1:0]       Ib6ca0cbcbaadb956d19a482fc099b175;
reg                              If33bbe9993ff895a7bd07bb8ee4ca970;
wire                             I605674982abba50698d4d3c2220b0db8;
reg   [MAX_SUM_WDTH_L-1:0]       Id52b94ae6662bb2137d8b9d53280bcdd;
reg                              If9a84cb15af69dab2d9e4ed921f4deab;
wire                             I201d44bd3cdf2b34fd2564188190b27b;
reg   [MAX_SUM_WDTH_L-1:0]       Ic3975e4171d618ba53e1569e4fc93440;
reg                              Ieba9f76cfb4c1a8069e2bfae0320ab0d;
wire                             Ia764576ce7e8ec4fc7120bcb8c038422;
reg   [MAX_SUM_WDTH_L-1:0]       Ib4e0f05afd881adf14a5eab850c75a3b;
reg                              Ic85dfb2e44272dea346bdb4352a88c44;
wire                             I66d5eccef31484a090c91507a3d38a85;
reg   [MAX_SUM_WDTH_L-1:0]       Ifb875d675aa28de930d889ae4d37b48e;
reg                              I9f0f8b22b39af997db900c486fc37a18;
wire                             I93cee05370c836746d1ddeb0f74456bb;
reg   [MAX_SUM_WDTH_L-1:0]       If98948e5f60b2c3ba1d7338e24dc0df6;
reg                              Iebc1dd048a5c7e83175ba1030a4bb587;
wire                             Iaa19be06695f47ff7d10667289dbde36;
reg   [MAX_SUM_WDTH_L-1:0]       I732bb69d248d700bcfdb287932839da8;
reg                              Ie8340c2226ffbab8f79e95ef17594210;
wire                             I21adefc729265cc5ae67ce279a0a78a2;
reg   [MAX_SUM_WDTH_L-1:0]       I403a8ece76036b3ce6277435609548a5;
reg                              Ic7dcd6d9c98422e20947712d0f4adc62;
wire                             Ibc0592b70bd60e475066554f0c7c4171;
reg   [MAX_SUM_WDTH_L-1:0]       I5a6cf1bdbcb2a342e548fb44c171aaf4;
reg                              I7df25ee69290c62782cd05715b0a6ecb;
wire                             I14f80574ea80b02ce13079854991febd;
reg   [MAX_SUM_WDTH_L-1:0]       I83a16a5be8d92896234bb9f2a36a22c9;
reg                              If904894b9cd6236c35bd9de268fab07d;
wire                             I09aae1dd6d02bd2a65dc7fa06fd848ca;
reg   [MAX_SUM_WDTH_L-1:0]       I6cad1cb66561eb6f0e3bfe5070b290c2;
reg                              I5b890a24c074e7f2ebfee20ce4e15951;
wire                             Idd698fb3a64825b43803642fc91bf674;
reg   [MAX_SUM_WDTH_L-1:0]       Ia50c447d5838d7979b2e19796be6221b;
reg                              I22f4468c482ed815d200d72ac2da570a;
wire                             I73c9bd7e52f6049b733b3a594ad6fae7;
reg   [MAX_SUM_WDTH_L-1:0]       Ief62ab0263b74086ae23a208da23e9c7;
reg                              I091ae78d995382a96c68c47a60844a9b;
wire                             I0fa2b3408156b2b0f656db4947670fe3;
reg   [MAX_SUM_WDTH_L-1:0]       I564999dcc2f67c8f82fb5cd16af0ee12;
reg                              Icbddf0d9df1bad66ea2f7352834bc759;
wire                             Ifd85deef561f76562208a8798b540b99;
reg   [MAX_SUM_WDTH_L-1:0]       Ifb0e4775ffb73bb2533844db969ab900;
reg                              I9a0db2b202a01aad173d2c8109cc596d;
wire                             I9d6eec32202aeaf66e7815492ac483b2;
reg   [MAX_SUM_WDTH_L-1:0]       Ib109fcaa55c3094cadb0c1f5f40ca752;
reg                              I724071f9e582e988d8f2d4c98ab9c070;
wire                             Id771356ebafcbb0e2bb8b03e49148b99;
reg   [MAX_SUM_WDTH_L-1:0]       I56aeb1bd0b0e9857d9cfd2c6b347fe91;
reg                              I31e8ca0bb1f64410501bb3c55bbb60fd;
wire                             I7f4f192560919410f2526392d10776a1;
reg   [MAX_SUM_WDTH_L-1:0]       I02651642fc35059fe9b4141c2fa1f34a;
reg                              Ib7b1834c1a9867cb8f42c9ab177dc11c;
wire                             I4e2247be1d2dd1af7467039a05447631;
reg   [MAX_SUM_WDTH_L-1:0]       I1f1e04979c8a5badc8a103809f76dadb;
reg                              Iaf22f59aaf7fa5f0e87a8d7504427627;
wire                             I5146e2d888c120b7afc430cc8d1dd34c;
reg   [MAX_SUM_WDTH_L-1:0]       I19fe22e1104703ddc9bbc94a5368bbc2;
reg                              Iea702a29812bf0e4b61cf21351648fe4;
wire                             Ib34be78c56c66ff7d85745612cd59f60;
reg   [MAX_SUM_WDTH_L-1:0]       I4386a95203c4fe83c6db7e25a288fc4c;
reg                              I05fa85d0596e05c1df86434a2083c4e1;
wire                             Ic6f48b24e0247c43666af5f25f03c1dc;
reg   [MAX_SUM_WDTH_L-1:0]       I2ddabc0b4bc45698fdd877c93bcbe280;
reg                              Ic61a806c6bc223d2c23cf24dbf3e85db;
wire                             If9f312c27d80be62969c60eb9b67586c;
reg   [MAX_SUM_WDTH_L-1:0]       I5adddbf99d0d39c5d70ec6a0978f3ef5;
reg                              I8284c12f98671842255420333096213f;
wire                             Ic7e3298aeb02d5829de1904288687002;
reg   [MAX_SUM_WDTH_L-1:0]       Ia24d776498719aa6cfbdb5df69d648e3;
reg                              Ide2e42206ceb5cc9ddd1646dea75776f;
wire                             Ib45f271c90e7bb32cba9dbaad5334c67;
reg   [MAX_SUM_WDTH_L-1:0]       I038ff8eadf1c551dc42d09fbadaea5b9;
reg                              I47512947d0532033dfa2b015aa107642;
wire                             I727821089976c74cd540ec58ecce2da2;
reg   [MAX_SUM_WDTH_L-1:0]       I102dc8709a274d21c09abae1d2ac1272;
reg                              Ia5ec36569a57a6256966da94a52875d1;
wire                             I4ed27d0c804891ee239ae8259d200712;
reg   [MAX_SUM_WDTH_L-1:0]       I136256458e71d84e850b61a950f279e7;
reg                              I07ea72a5755bd2b0da6e89389df44f69;
wire                             I421ad50f600133f1e7f6a52625181d36;
reg   [MAX_SUM_WDTH_L-1:0]       Icda6fe755f2d840f8e404d84b231e827;
reg                              I89b6e7810b2a5d45238819a6a171dac6;
wire                             I172379505892287217e08c060285018b;
reg   [MAX_SUM_WDTH_L-1:0]       I1f6cd53f31f27d86d78d5079e84c9716;
reg                              I2e6141be9be5edab8e67a1e7f640903f;
wire                             I8ac36cb7b4e56689efd4a3de1fafa0cc;
reg   [MAX_SUM_WDTH_L-1:0]       Ia1f69042d447cb17772b29f634344b53;
reg                              Ib438d8ef5fdd32b2811e0e755acdfefb;
wire                             I002e83f2fb7e5b07710a802aa505b2bc;
reg   [MAX_SUM_WDTH_L-1:0]       I84648f139f0fd470a62f0638aeee9e97;
reg                              I21cc09d0a95b4598c5614b7af3c6fe03;
wire                             I26fe780ca6becdc9f86a7be04c6257d2;
reg   [MAX_SUM_WDTH_L-1:0]       I6ebc0ad14d76d3a80a4929ba8b5e7848;
reg                              Ia7a6617c92f999d7c19d3c338cc60e8f;
wire                             I3a8d18e570ec3aefcdc29d7bc783dfde;
reg   [MAX_SUM_WDTH_L-1:0]       I26cba2d4920ff7fc40b1723c29ed8391;
reg                              I5ea3e9e13e199daf8df53389a405cd0a;
wire                             I4ddf83c90adcc1bec65f265e898568fd;
reg   [MAX_SUM_WDTH_L-1:0]       I27980b3a1936a92a1751588f91a5f542;
reg                              I5a202e3ec847e13fa21134123db7a027;
wire                             I0c06a37e120e59f19578c68801a4b6ec;
reg   [MAX_SUM_WDTH_L-1:0]       I5464cf638e0ca778d4e113b216084180;
reg                              Ie697e69bd62cf7bef4a4934843967cec;
wire                             Ic290ad8aeb51c16106f9311b06134a2d;
reg   [MAX_SUM_WDTH_L-1:0]       I1804dfc05236c728f563342eb011f4f8;
reg                              I6979425ff99d598782f2a45b1d463f8d;
wire                             Ic4c7c898ca601e4d44076ec5bb475979;
reg   [MAX_SUM_WDTH_L-1:0]       Id219264de5f6b67cff866b2bafc660b5;
reg                              Ie735fb63c3d40f44ede25d0a213847a8;
wire                             I380cd867541300f76fc359d72f49bdbc;
reg   [MAX_SUM_WDTH_L-1:0]       I03e4f803d4b82aa774662e02b188b0a6;
reg                              I2f132b8b367a5eb3d7029b1c27991dbe;
wire                             I350f20848080cffa45a31e2f1e553a3a;
reg   [MAX_SUM_WDTH_L-1:0]       I32e079707d9ce4b31aea8fd2c998c27c;
reg                              I55291a60dc5b1255d71ab749eaba0404;
wire                             I912b9be8432d4eb792d79566a8280703;
reg   [MAX_SUM_WDTH_L-1:0]       I488f60405ded7af04c941bdbf55290f8;
reg                              I804b17fba020affb1ed32666d73607ae;
wire                             Ifaed59e29ee3ee9166192bbbf04bc682;
reg   [MAX_SUM_WDTH_L-1:0]       I26d314b69785bdb0ca8cd52c258c3b35;
reg                              I478f85d129f1f538304e6cc74b9d2234;
wire                             I7eaa9f70586b12e371db5964758ee7c2;
reg   [MAX_SUM_WDTH_L-1:0]       Ia490437ab050e63e611dfb4d9366017c;
reg                              I71ef5d9d9f272131a3c7bf864c0b4863;
wire                             I9a8946bbda4bfe72fab3c2f59533b3ae;
reg   [MAX_SUM_WDTH_L-1:0]       Ia6cc50c8b7f83dd80d7058eea40338e9;
reg                              I65ed551a24cd36ae20d1ffeac42fb99b;
wire                             I29fd8dea7c3c39722614210cb7f65851;
reg   [MAX_SUM_WDTH_L-1:0]       I3652208cee3ca6dcdef63b7df53e4329;
reg                              I4c99cb1e56179799079d9a484edf2a02;
wire                             I54bed2059ffd24ac2fa91b038c0256ae;
reg   [MAX_SUM_WDTH_L-1:0]       Ia9a4760f6a2bf8f8f660e2b0c31dd823;
reg                              Ibd985ec8f6f4eed7f14ae2692367cc00;
wire                             Ic3608e6a6c45ee04ccd8198c88c69003;
reg   [MAX_SUM_WDTH_L-1:0]       I5ec267a535ad08c629940d70c61894a5;
reg                              Ic7eb65782a34589e2b015442172d7568;
wire                             I37da881d3575c055944719409ddb66f1;
reg   [MAX_SUM_WDTH_L-1:0]       I17fadd913ac1008fcbefff48ad366d8f;
reg                              I3bb60f8d4ccc5e40e97af6f6718c90c9;
wire                             I2b6999fd13f9e57ea33c0b4602594c66;
reg   [MAX_SUM_WDTH_L-1:0]       I275728fecbd15ba77f57860bb329da16;
reg                              Ib109c4220b1113561ec1319a0ac74498;
wire                             Idee62819bc831a9ba7c73dea46f3da9a;
reg   [MAX_SUM_WDTH_L-1:0]       I8d0bc446761559f2188e78200eb0a895;
reg                              I91ec97b5793a453f81b1780157e12d47;
wire                             I48c95e9ee4d7dd54b6bf21a9a5b20635;
reg   [MAX_SUM_WDTH_L-1:0]       If9fc4683c2f0545e1f077541fd25da66;
reg                              Icae10f8dc7273f91884f011b6a88cf91;
wire                             I26b2a20b53a3ef8531d6798c4b272422;
reg   [MAX_SUM_WDTH_L-1:0]       I1c8e7559160d5a1fe1fa0002cc414d1c;
reg                              I8b7efa4f096bf761a8df08d1a3f1b77f;
wire                             Ib814d21cc76c4f3135a4aa813dcb748d;
reg   [MAX_SUM_WDTH_L-1:0]       I059014ede8b9092d817c0aaa1c7ed388;
reg                              Ib0dfb26e39fd974f64d54a0f9c0cd552;
wire                             I44dcb4df87d1cf32ee2c9bea836223ea;
reg   [MAX_SUM_WDTH_L-1:0]       I6294fc2c9181871210e0cfbb9834c3c7;
reg                              Ida3a51bb8109fd4c3e494b736889efaf;
wire                             I96ea91e1bf398f6b2973e815a6a10aaa;
reg   [MAX_SUM_WDTH_L-1:0]       Id24dd0ede5504678fbd809ffbacd0dcb;
reg                              I6a47d611882f8af53484f22ce5b74fe6;
wire                             I75458b8dd7bf267526c36af5cbfcaad1;
reg   [MAX_SUM_WDTH_L-1:0]       I496994e784eb114337ac9e78ec0c4d3f;
reg                              I52af26697dd18d51e902642e19045d9a;
wire                             I230ed2d0ad383ba3a6b5b69ce09ab4b6;
reg   [MAX_SUM_WDTH_L-1:0]       I44c28351f261765c28a066a581c27c13;
reg                              I38b0b02379864bed0b097754dac42dec;
wire                             I6c09d773366bca735c15703f7c2c5a11;
reg   [MAX_SUM_WDTH_L-1:0]       I84419e016619a3a33224eeaba85e68b3;
reg                              Ic3f80e7837ab46f58cfd4b6c775d4e72;
wire                             I146e4737d01377560ffeb78fce84973d;
reg   [MAX_SUM_WDTH_L-1:0]       I67d114d975d5d65f575bbb8c819fa22b;
reg                              I87b9dff79eb8389488e97e427d59d767;
wire                             Iaa4c0cb6fd4dcc74d6ffd2bde42b7947;
reg   [MAX_SUM_WDTH_L-1:0]       I6a452adc2501774b55e5fe73c642ea26;
reg                              I44926d094aefc5aa52713fb52704f84f;
wire                             I49d021b0957d65a6c2608de826c2676e;
reg   [MAX_SUM_WDTH_L-1:0]       I33792929f4428ddf0629231288e459ec;
reg                              I57127b05215e4faa4e32d5ca38611eb2;
wire                             I72393e4bfc85c2b9ee24a4395b3568eb;
reg   [MAX_SUM_WDTH_L-1:0]       Id0013f18ab77416e08d994c360b13473;
reg                              I79aadc384d50af92ae1af6760ffe3b3b;
wire                             Ic9f855b66d25668256912f2e434b4854;
reg   [MAX_SUM_WDTH_L-1:0]       I5683f67c7d462c01c55b8be9b6d1fca6;
reg                              I28effe4aa10b24a221d5e1c84f2c21ff;
wire                             I27fe4e83261eb6a1789a8f7d77a0caf1;
reg   [MAX_SUM_WDTH_L-1:0]       I4a5e3cf3066a4c2f7f5f8dbe824ff88f;
reg                              Ia0d7cfa22522e5b4f7b545aacff7fa59;
wire                             I45c158cf7145668cb8524f7fa06f9302;
reg   [MAX_SUM_WDTH_L-1:0]       I93879adfa4333a80be696d846e34d799;
reg                              Ifdac0b0a75dfcc09291fd95e842e68f1;
wire                             I16d2a9270452f0d8b6eda06ea939fc6a;
reg   [MAX_SUM_WDTH_L-1:0]       I199e944b303446e2cdafb6f34d0d12c7;
reg                              I1bbd0d48cc6bd8a4d4d520d38798f74c;
wire                             I1ab974ad9718ea8350d76bbc1510d2d1;
reg   [MAX_SUM_WDTH_L-1:0]       I91d282de42df72b1c439fede384d6336;
reg                              I06ede5ab6bc97827c4f866dca1aa17bc;
wire                             I31467f39d6b5c20d4e155d19afa34e95;
reg   [MAX_SUM_WDTH_L-1:0]       I8a06d2c278af9d552fa36a61128b8a9b;
reg                              I4b7f22e0b9e1589fbc1d558b37cceb37;
wire                             Ia8762fb956b52535ad6921e9191288d0;
reg   [MAX_SUM_WDTH_L-1:0]       I5a36e45af7599ec00703dfc81f9d1176;
reg                              I6e63e4047456268e73ad16a5cde93681;
wire                             Ia018c4c165c5af9a329a63aa365ac038;
reg   [MAX_SUM_WDTH_L-1:0]       Iae09429ca8733186fdb3c50f36895746;
reg                              Iec7997b0018f4fb3572579a5bf1e4728;
wire                             Id85085de57a0152aad8cf5e27a195052;
reg   [MAX_SUM_WDTH_L-1:0]       Ie5f74b33d06ddb8b32b57c8c82392001;
reg                              I11cb6032d99f05b3f908418a70fd3d6e;
wire                             I461b443279e5bf47de450846e3da7d8e;
reg   [MAX_SUM_WDTH_L-1:0]       I7d3cdb71cdab3a85122130207d872476;
reg                              Idba56a073e34e530c36025914f7646d9;
wire                             I71d07a22b66aed8c24fe4dd203869fa1;
reg   [MAX_SUM_WDTH_L-1:0]       I68ae9f2a14b161c940f6685073eca97e;
reg                              I3a7582a1c86f2b49979372132ce98c87;
wire                             I173b85306dc75e596cfe67f7c518f36b;
reg   [MAX_SUM_WDTH_L-1:0]       I778f907b5eacdfac02b0bc4547af4ea3;
reg                              Ifaed912ee00082f8458ae37bd47179a5;
wire                             Id57948138d3091aa350db0d906b06b34;
reg   [MAX_SUM_WDTH_L-1:0]       Ibcea5bf1e21fa764ac9f2d2702c8f79a;
reg                              Ibecc30f33083404bf48eb0005e14bb83;
wire                             If6b37dd338e28ffd7fb888bc56f716d1;
reg   [MAX_SUM_WDTH_L-1:0]       I93a3e1a8e414d4775f19c0c9f16d07a8;
reg                              I87009d289b53c6e366b73e275e414caf;
wire                             Idd412a66c4a434eaaf337b6b4ab6b0a5;
reg   [MAX_SUM_WDTH_L-1:0]       I8772034840834e51187950d320f9eb40;
reg                              I5d5b08cc3fd13b96621143655a806c7d;
wire                             I5829341b8f12f906ffc53c9d716e6556;
reg   [MAX_SUM_WDTH_L-1:0]       I3d0aa00b61d4684ad46f49329197c901;
reg                              I94ce074b29f44c5e4a63ff6e00d2b9c4;
wire                             I449b6fdea575e92fa4603f141ff359e8;
reg   [MAX_SUM_WDTH_L-1:0]       I146866a6d46604c47d87afa3c88308c6;
reg                              I2fd3e923d1adff22ef7718dae5632b29;
wire                             Ic6581fe8d97a45b71a1ca8d9ec97f97b;
reg   [MAX_SUM_WDTH_L-1:0]       I84cf7aa78617faed2f1762bb1961cc0e;
reg                              Ibe2d184a52eb5d33cac0ca4a5dab55f6;
wire                             I4af6879c6d4d2b96562b1c2ada8f92b0;
reg   [MAX_SUM_WDTH_L-1:0]       Ib1f43a0b9c86d236b2ed71c35c296b9c;
reg                              I0907dde542619e162f45f3dac8c0c16f;
wire                             I7a176a15ab2c5396639be387bc43896c;
reg   [MAX_SUM_WDTH_L-1:0]       I88aaa7538f9007ce204319ec639d1c7e;
reg                              I9bdfa0d38ed6d215e7ef7ecb12185b60;
wire                             I38c29f53b042f039a908cca7d09cc2bf;
reg   [MAX_SUM_WDTH_L-1:0]       Ie3a171564602e9936d7960e83bb0fb3a;
reg                              Ie0e096809efa587a070562473e9a2fff;
wire                             I1e5c60072bcfdc56b1928040edf9ecb2;
reg   [MAX_SUM_WDTH_L-1:0]       I732b452fd9521b3a13ff1f965c443325;
reg                              I8c2c0b7861868365bc3935ef8d0fe309;
wire                             I03998667df412d12539d57112b6b6f76;
reg   [MAX_SUM_WDTH_L-1:0]       I16cd75fd747b600e90763d8ce9c08210;
reg                              Idde6e2f615f8ec0aa66b7397e5581651;
wire                             I2ae5c6ae2de0db31a656018e19d086b9;
reg   [MAX_SUM_WDTH_L-1:0]       Ic6a7d6bfb12f40ae8823db716cfe017a;
reg                              I3098e45c14ec08213883f7879c30150c;
wire                             I1e27f59e10400144106861daca51e721;
reg   [MAX_SUM_WDTH_L-1:0]       Iea38a3c260d0caae4ae042264a0f4787;
reg                              Ide3c2fa1d5da990a0566c65a12d1d7da;
wire                             Iba8577f8233fe013584171e588868e69;
reg   [MAX_SUM_WDTH_L-1:0]       Id6240152bd22a9655b18bdfd91812e03;
reg                              I6ece8c59f986da73f00e104ff5966189;
wire                             I1d0a95c7cced8ede694d02936af63047;
reg   [MAX_SUM_WDTH_L-1:0]       I07eeb34c9dfb9baadb9f263b6f095ecc;
reg                              I5c002c1ec0c63a2c04ca2711fde50254;
wire                             I8b072ed41d990e6afa6fb5d22990f4df;
reg   [MAX_SUM_WDTH_L-1:0]       Iedb57db3cbaca9f9a469d91ed81466a8;
reg                              Icb5a521ae9f45d8c9101fdde8925e64f;
wire                             Iab0f19858a1a01fe09fa3c99d92a79fb;
reg   [MAX_SUM_WDTH_L-1:0]       I2972b771a4e99ddfa2178349a805b16f;
reg                              I7b72bfdf546647380e6b1f9a810fd1d1;
wire                             Id88441b410f55c15465eff4cfa216691;
reg   [MAX_SUM_WDTH_L-1:0]       I6a61cdadaf987763080e6ce4d1605ee6;
reg                              I84581a99221f2aab1e7cbbcc80296ad4;
wire                             I894540936535dd20ff1ea5c47546e5fe;
reg   [MAX_SUM_WDTH_L-1:0]       I12e430f1ccaa6099ba9ff803c85d9532;
reg                              I27d48bcfb04bf11d76b496d459ee1b48;
wire                             Ibb40a1e09cc59e00ce8ba1460e0712d4;
reg   [MAX_SUM_WDTH_L-1:0]       I2cc3c84149c81572357c01219248aa3b;
reg                              Ib89fb8b901f12120ab0bdff5207c74f0;
wire                             I5349c1efb5233e8cc6c472ecae80ccc3;
reg   [MAX_SUM_WDTH_L-1:0]       I6d4b18dbba5c2b058f93a8d46bed38ec;
reg                              Ic2324007897bedbb70a77faa1fd301ef;
wire                             Id90c5bcfdae1c4abdfa194477917dfbb;
reg   [MAX_SUM_WDTH_L-1:0]       I32ca5d01c39fe736d6ed57d70fcbd555;
reg                              Ic75af8091015d4615d0c059ceb16371b;
wire                             I1dafa9e7b2a353dee90a0b0f9685a826;
reg   [MAX_SUM_WDTH_L-1:0]       I8807f2f633d64cb064fbc149ebd30412;
reg                              I5b98fb653fa4d3d4ce2ebccd24085f95;
wire                             Ia75e6368415ff53bdbfe81ac2bdfb290;
reg   [MAX_SUM_WDTH_L-1:0]       I822d3b3516499e58ee7777b99259a206;
reg                              Ic9320f9ad332f511422f5b805de9488a;
wire                             I91217ca822fb03fdad03b8d005edadc9;
reg   [MAX_SUM_WDTH_L-1:0]       Ie706bf8dd49322fc1d5d83e40fb20f04;
reg                              I71574a4f01fc2e2fdd051a90b9115524;
wire                             Iccc6e66d1f26c4a5874ba02980dad6a7;
reg   [MAX_SUM_WDTH_L-1:0]       I9975f2ca851119d7ec85cfdefda150f0;
reg                              Ia59c01c2e6f19ee93a091dbd1a1da83c;
wire                             I15e9479f1c9aae3c1f12f0f301ee275b;
reg   [MAX_SUM_WDTH_L-1:0]       I2e0639bf4e48a7b1486beebcc9ad7c0c;
reg                              I5e8e70c7ad583c0c4f09cacb60602c00;
wire                             I14692ccb24148a020dda28c6f61e3611;
reg   [MAX_SUM_WDTH_L-1:0]       I6131789039de7dc431c3b9b59ecb7654;
reg                              Ia180d785ba74d63500c25e3a04d21c03;
wire                             Id237c89ded30e926343fb68d786a76d0;
reg   [MAX_SUM_WDTH_L-1:0]       Ia20482fd064712397fe2f9f77f4d854b;
reg                              I4dbcb057b2076d4efd4e05e818d976c9;
wire                             Ib56bd244f7a9876fab3d51a21ef163c7;
reg   [MAX_SUM_WDTH_L-1:0]       If052875ec5a78a68428a1ff09df623df;
reg                              I24e240c3d018053712e0fb7f861acad7;
wire                             Ic1db9806badd4e959a0f0a769e15b6c0;
reg   [MAX_SUM_WDTH_L-1:0]       I2e27abc9297a3fa647f50859af7cb094;
reg                              I78d4209646fe0f2b8027988024b947ae;
wire                             I3649823bb60a4740b6a7f94dd26e45a1;
reg   [MAX_SUM_WDTH_L-1:0]       I5d5e3b64ed1ca16d65d8eadb8100fa06;
reg                              I62fa50cc71ade42b52be1de668da6b7b;
wire                             I8d7596d25b93595ffa1ef7d273c98c14;
reg   [MAX_SUM_WDTH_L-1:0]       Ie91a08b49b9bf23270dd3fa331e64968;
reg                              I5145e1005293c49c849599347a4a2b46;
wire                             If607fe1cc3901fc74590a81a26ccb4a8;
reg   [MAX_SUM_WDTH_L-1:0]       Ib599712a1e8fadbdf7e3712bca6c0b74;
reg                              Id77a6df77f3d714b6b1f60bad2462f2b;
wire                             Ibe2cd0729747659786b76f044f3caa6e;
reg   [MAX_SUM_WDTH_L-1:0]       I1791c009b0838ef10233015f80a5c4af;
reg                              I6cbfcd474a5a76538db10b8c3235986b;
wire                             I38e96074261512c31ebd15c6de4b440b;
reg   [MAX_SUM_WDTH_L-1:0]       I3dead2d8d18ea8503a578469625f3aa3;
reg                              I17c80f6af6d201a1214d251778a9e534;
wire                             Ie72e9c0aa298ff1809a47908ff86b6c4;
reg   [MAX_SUM_WDTH_L-1:0]       I2fc47140b9df2544d7ae9c82cd38ebd6;
reg                              I468342d7ba88b0a9313f38d0ec2a81e5;
wire                             Id6e349e3f114f328958052a680a95411;
reg   [MAX_SUM_WDTH_L-1:0]       Ice09150d69c67cd2d08d6e63b8a9bbc7;
reg                              I189be0be892f48991d69acf5a0d42533;
wire                             I6dff6c5c76c92ba9626512b35a573ac8;
reg   [MAX_SUM_WDTH_L-1:0]       Id67765c4a6b11f6ee0a4524ebb2d1ca7;
reg                              Ib5bdc1c490d7d2fd11359fc6c79372cb;
wire                             I5145ca1a0b7eb68adb93316264ed0084;
reg   [MAX_SUM_WDTH_L-1:0]       Ia17bbf4b7f063de0bf0701276b7b0c20;
reg                              I85e112a43fa9046e94da6bdb7b3a13d7;
wire                             Icff67cd5e9472e77380eb812deb625b6;
reg   [MAX_SUM_WDTH_L-1:0]       I9f9075a7745d475331f0b25bad830421;
reg                              I03ad487e845cce369a813b0c7f32e59d;
wire                             I88adcddd217c9b2363fe254b0be469e2;
reg   [MAX_SUM_WDTH_L-1:0]       I4d832ef88af4d4244516b0bdfd2b461c;
reg                              I85aeb073e949fc999464ce61479790db;
wire                             If149258ed84a848bc38011bef172b6ea;
reg   [MAX_SUM_WDTH_L-1:0]       Ib2038174dd555b1d058778fa904aee65;
reg                              I7534524f9d9c64bdf0bb88ba351b3ca5;
wire                             Ie70f8bcc335351e60eecd70b90d4432c;
reg   [MAX_SUM_WDTH_L-1:0]       I959dff5d57b4c2adb85c3602d5874c90;
reg                              Ic4a902801adb86fdb2481f5b868daa8b;
wire                             I5277100478097db96b41fe0988046442;
reg   [MAX_SUM_WDTH_L-1:0]       I30dd112c5a6793cf37bfaaf8dfdebcaf;
reg                              I1141271b2c1fa529b7f4e4ce9ac10c95;
wire                             I0aced2534542d8d2c488c7082ca214ca;
reg   [MAX_SUM_WDTH_L-1:0]       I4d4a0930420b4d7da8b6e91b2b25bc51;
reg                              Ie62709fd754ca31b0e5d830901bd6433;
wire                             Ifad6157e5199a5b5dbd2465f4cae5b3a;
reg   [MAX_SUM_WDTH_L-1:0]       I7ae1d318fd0df386e0c8bcf0f0a94e4b;
reg                              I6c6a99a66fe46ca1532fa898123a6131;
wire                             I2bf55a177a00da61ccd463a450de2bb0;
reg   [MAX_SUM_WDTH_L-1:0]       I06cc62e12d5a261d672b5428dbc9767b;
reg                              I963a6698cd1f83ce4e7ecaff7f53ce25;
wire                             I521e3e69d81a6034183d2ba861ec7726;
reg   [MAX_SUM_WDTH_L-1:0]       I9798b16b4658501d739d46182d7ab169;
reg                              I451d9f14e13b272ea041178627ef7f56;
wire                             Ife32264cdbf7445987f5f39d6361d1e4;
reg   [MAX_SUM_WDTH_L-1:0]       I90bc85b7a6e56250bf13407ddd32bf11;
reg                              I3e7f571589d773eaf3435c03bd13c9ca;
wire                             Ied102cd26c4fc50aa354b16a35d3490b;
reg   [MAX_SUM_WDTH_L-1:0]       I88990d32bd34da606660f1c078b36ce0;
reg                              Ie823a06acbb6935875c5cb9088389b27;
wire                             I5900a9bf6a83b1965f0dd9749d90e317;
reg   [MAX_SUM_WDTH_L-1:0]       Ib32ce57f2840a45fce8e66f71b37719d;
reg                              Ia4c876fe77f09258fb130d03b8cdc67b;
wire                             I1b4d2bc08a78865fb281a44e84088fa5;
reg   [MAX_SUM_WDTH_L-1:0]       Ib0179c2048d6c9d1865d171b48c521ff;
reg                              Ie6bf8e5060074ce2dfcf7ddcbb158bff;
wire                             I70724327149d97d4d4f3f71a1500427e;
reg   [MAX_SUM_WDTH_L-1:0]       Icc8ffcc0641f0f9405590338e6b5e517;
reg                              I706ad22942f1cfbfae4fde958450189b;
wire                             If91997f00102c66a7630ffb2d041d949;
reg   [MAX_SUM_WDTH_L-1:0]       I5d6cb688ef094e1f119d8536f0f56766;
reg                              Ic64d1cde239aef0df4f227a64762f9f2;
wire                             I25da82603d45fc12f685407e8dc2f6f1;
reg   [MAX_SUM_WDTH_L-1:0]       Ia5aa7c66d2818982a661e4d048876d1c;
reg                              I719f60bd29522fded995c8230b4f3a34;
wire                             Id2fdc5b6c996c567743aaf021a5e6371;
reg   [MAX_SUM_WDTH_L-1:0]       I449e514b6afb3e8e337691fc64f7431c;
reg                              I1bd8505e6f316488bb1cdd74932c0314;
wire                             I8d57ad30940b8351a829b8ca99921a10;
reg   [MAX_SUM_WDTH_L-1:0]       Ibbd5f0906646560a903abcf6848ee80e;
reg                              I63e645f447ddd1fc9409879872479bef;
wire                             I2ccb382adcd7799634c86273c8a39199;
reg   [MAX_SUM_WDTH_L-1:0]       Iee607ab8132caf0f678324d20394f533;
reg                              Ia8298013e67424c2d5fbe03634170080;
wire                             Ie521ecd231d7bfedc8de182c5050f6de;
reg   [MAX_SUM_WDTH_L-1:0]       Icc90fd3c992755ac7e4aec1370600e06;
reg                              Ib404a1296714f45ddca6351a918ee875;
wire                             I855892c34f1706745dda4ffc3e5e5a98;
reg   [MAX_SUM_WDTH_L-1:0]       I81e0ea92e07ed7d29b4ab769443b55d3;
reg                              Ic08905e9ffee26c630277db86cd5be95;
wire                             Ib945fab3df6e5a7494b7fe463384ff4b;
reg   [MAX_SUM_WDTH_L-1:0]       Ie7554e9d2bb6287b440973a9effefb50;
reg                              I674e937c017f29d18946139b00db02d8;
wire                             Id4fa22c6f8634ae38892953bd6ab55b5;
reg   [MAX_SUM_WDTH_L-1:0]       I3fd483389e4ddb927e7be7636441f0f1;
reg                              Ib3f5f61eaba0c2dfdf6c75e46e4233f0;
wire                             I3d8295457058e1d34bb136753b69aaae;
reg   [MAX_SUM_WDTH_L-1:0]       I3d7a6bd63d9f66b068c08cf9046474f7;
reg                              Iff1039ba558287ef96daa7dfd15d6294;
wire                             Ib8df0659486e8ecfb5c52bc2db3a8436;
reg   [MAX_SUM_WDTH_L-1:0]       Ifdb5bd8e8237676fd8d2816bfa53f0c0;
reg                              I017268444024bc19b209dbb4322de15c;
wire                             Ice8927db6ef88a90daf77ea5be2a34bb;
reg   [MAX_SUM_WDTH_L-1:0]       If2865b698bf9c511fcf6724856074335;
reg                              I22e4741c472c64c846742391d81f682c;
wire                             Ifde5beb333f350ce581a137dae22b99b;
reg   [MAX_SUM_WDTH_L-1:0]       I077ad1ef2fe0a7e791fdb45026788641;
reg                              Ie3c87a536250268b1012b6166173108b;
wire                             I9fe47549e560319ae8decf04a9db5240;
reg   [MAX_SUM_WDTH_L-1:0]       I4c67ed6284da547b599a4602a3cc51dd;
reg                              I54204328537dbc383a3a03352e9d6fb6;
wire                             Idcda31b4dea85b3acd88cad806aef569;
reg   [MAX_SUM_WDTH_L-1:0]       I3d0babc64a3400a1ee57fff14920d1e3;
reg                              Ic5d81213c2d23b0549006ed162d9e6dd;
wire                             I54da9f6048b299dd7e94962912b86407;
reg   [MAX_SUM_WDTH_L-1:0]       Ica1731833fd3d6a881b3a17a5916f7e7;
reg                              I0ac628860f9fb9e6daae572ff007f34a;
wire                             Ib1da5f847077624a37594c2db1b444fc;
reg   [MAX_SUM_WDTH_L-1:0]       Id5705e57bc5c050342e82a302b73902e;
reg                              I2487101836608b77528a49d037c40fb6;
wire                             I80c640a2bc35e9012dfdda839dc5ed1a;
reg   [MAX_SUM_WDTH_L-1:0]       I4606e0ec878c615753206459716b5d25;
reg                              I99d49fb5c921d2d837ac7b02716d9ada;
wire                             Ic81ffedc7f65fc4d390acd0a30d5e427;
reg   [MAX_SUM_WDTH_L-1:0]       I5ac4f231a175a60f63db8d4d71cfabaf;
reg                              If4d0af4a78a49e861adbdb1a3f6e7ae9;
wire                             Ied3448df1f31122d619b1a4cb316f200;
reg   [MAX_SUM_WDTH_L-1:0]       I26a3cd9ec3a564df04ad20559039598f;
reg                              Iccefd72e7e22a425ced6974251245da8;
wire                             I017d4243cafbd5d4d615393de3a29aa8;
reg   [MAX_SUM_WDTH_L-1:0]       I26801bb91e66797982b66ce815da85a8;
reg                              I3fcc5c32415df9710be01f0f35ac68e5;
wire                             Icb2adb3572c2ac780b4fb413c6ebb375;
reg   [MAX_SUM_WDTH_L-1:0]       I3b617a013c15e8b623ad517e08df3a00;
reg                              I0bf8339802110abb8bc94e481647f25f;
wire                             I711042dda213300a90c51b09057b64b4;
reg   [MAX_SUM_WDTH_L-1:0]       I65f5f9a3f7f68f4b2fd7695ce6bf4629;
reg                              I6ae57b8d68417d1ea8ef70d43a943e0b;
wire                             I59b7772e832e814877d4f9e7726f5143;
reg   [MAX_SUM_WDTH_L-1:0]       I7d405b59e360b17d7f2eb1805b796fa9;
reg                              I07dd0ed55fbdeaace398ab7644a5189f;
wire                             Ida6ee8eeec2fa7a6bc1eeb8b5c3fbffd;
reg   [MAX_SUM_WDTH_L-1:0]       I033ad5c570f42830b265d7bf6a102757;
reg                              I69cfa3967387c5e8e48994b6466673a0;
wire                             Ic7fb6a8351310bd93953232556a692ab;
reg   [MAX_SUM_WDTH_L-1:0]       Ia00376ef5aca6a428280f2dbf25ab1cb;
reg                              I2ce599e7a40a71d9fe09f80269accc31;
wire                             Ib2ff62fd117b50bc0c190b8111b85f4b;
reg   [MAX_SUM_WDTH_L-1:0]       I252b17144e39018fda208bd18b555c09;
reg                              Id424746e76cc70f9292ed41659973621;
wire                             I4d46847f77bb17019eaba7ead1549a87;
reg   [MAX_SUM_WDTH_L-1:0]       Idb756c313694457c14b02431f3f076c7;
reg                              I45528f9be6a8f9a0f646d83223307e79;
wire                             I1d6145f5c5d5049a1ba3f3ef8a09924e;
reg   [MAX_SUM_WDTH_L-1:0]       I0c1545b312d755b14ee27b399a1d3079;
reg                              Iabcd2910bddf2e544c707c553b2ef370;
wire                             Ie5e08b5111cd2baacecc68000f84a9ef;
reg   [MAX_SUM_WDTH_L-1:0]       I903842d13327b74a952be0aa6c7ab0e8;
reg                              If01521dbf7dd9aa5196a9130ba47b149;
wire                             I3d61c9137cc0cdc892bc50c659fa8c47;
reg   [MAX_SUM_WDTH_L-1:0]       Ic461c1b7bd09b59297193d388c525ece;
reg                              I9284cc53534eaf3d6e5b4e9d9d93bea5;
wire                             I15411a1495f104308964c62a1ac7fe6a;
reg   [MAX_SUM_WDTH_L-1:0]       Ia14490057ef27f5df5f1b23ca6440a65;
reg                              Id5fdf11f0bf10ec37b11ced0a3268ad7;
wire                             I99f350aa0b468f89e8ac4b3da627a81a;
reg   [MAX_SUM_WDTH_L-1:0]       I2d3c1e36bd952fdbe4fac5f3af07e666;
reg                              I36cc6827c8e4c7831078c8f9972ee78a;
wire                             Ie23efd54df7880569e2d45a8572c02ba;
reg   [MAX_SUM_WDTH_L-1:0]       I7fcea0a5f9987b2414ab443bd07c05ad;
reg                              Ied6cdc5d7aa6335b2c32d8ab6ee6d889;
wire                             I29de3d73d38639aacb693c8080f4a168;
reg   [MAX_SUM_WDTH_L-1:0]       If0f5bf08d96033f6281121230c1e47c9;
reg                              I70709dd8c55168e62143f56d0bda1239;
wire                             I09fe5010524903c8b34892f6c308d670;
reg   [MAX_SUM_WDTH_L-1:0]       I19412627d5c573ceaa981cd7f1027e83;
reg                              I73ce9bd4312ce9a6cdc0c6b6aec72a55;
wire                             Id1af840781c6093921ea2feef85b6bb7;
reg   [MAX_SUM_WDTH_L-1:0]       I7c72a1709b233f745fb0323d04bfeb1a;
reg                              I9d0fc48c488109406aa9cfef80ac3b48;
wire                             Iab8c6e113a90faf59bb550681b0dc7f7;
reg   [MAX_SUM_WDTH_L-1:0]       I2639cefc25ac6f4982e4eeccf8fa810e;
reg                              Ie09336ee55ee45ac0297849f7b814f4d;
wire                             I2110f3928229bc70d8ec9ec7f1c92520;
reg   [MAX_SUM_WDTH_L-1:0]       I76340f05f74b295583bd9353884979be;
reg                              If919b9778437e1c4366017968d1ea582;
wire                             I0befd079483b2da8d410fa137f71d801;
reg   [MAX_SUM_WDTH_L-1:0]       I00974459262f29ec2b5472472e49faf6;
reg                              I71cdff133cb7a645e623c4bf06588fc3;
wire                             Icd1a2b8c1a50f9a1bab48ebfbb87ca73;
reg   [MAX_SUM_WDTH_L-1:0]       I075efbd3c4d87df8d733f0b3db008b1f;
reg                              Ie7fd0410103d16e27611f9ac30c657da;
wire                             I4422278d28ff2a983cc3a4ad8f2d655f;
reg   [MAX_SUM_WDTH_L-1:0]       If8bd6a5d380075f1ee7f7a4542531dbe;
reg                              Iab93975104312336985d4736015098b4;
wire                             I3fc4400a93546df2e2aad374a4d8c7e4;
reg   [MAX_SUM_WDTH_L-1:0]       Ib81b730d107434503c988ab9f00e1605;
reg                              I564a4d4a94f9951d85287b2ac35479fe;
wire                             I6c6a02b572e98d30ea5a0406be5cfd11;
reg   [MAX_SUM_WDTH_L-1:0]       Ib05cffa1bb31054450391bf9e17f8ef9;
reg                              I09c5b4146a3c48ae706d3041ddfe074d;
wire                             I91c29953d4b53657da39b53d8c909fd8;
reg   [MAX_SUM_WDTH_L-1:0]       I627097c06e3be5a4385171f3ec7ae5c9;
reg                              If205c7d745e5372ea61afa389f1af2c2;
wire                             I10441dc2915fcece28b38aa6b4156f5c;
reg   [MAX_SUM_WDTH_L-1:0]       I76e2c6001e1ae97670539bd471fc74e8;
reg                              Ief37a022c34d4e670413f5b7db306876;
wire                             Id26aa7283f70b13f1eb0b97ab1222da7;
reg   [MAX_SUM_WDTH_L-1:0]       I8b4433056d26f4aa60f18418b0114930;
reg                              I5ac36d471eec2b3ac068a2d20283f674;
wire                             I98b4bf6c27d9420941d252a98806344c;
reg   [MAX_SUM_WDTH_L-1:0]       I99601176686afd8fb85a85ec43849e6f;
reg                              I68acc6967dd156d6373abd6cc620f247;
wire                             I7814b43f7573d005d6b9350b311f93df;
reg   [MAX_SUM_WDTH_L-1:0]       Iad8276d5be3d9c6fc085465f05ac2aed;
reg                              Ic830033c7861645951982dc630e3385b;
wire                             Ia378bb83b0f76d4bf7de347a8bfd20cb;
reg   [MAX_SUM_WDTH_L-1:0]       I5e5dfce3ceb4fbbfce344bd471901736;
reg                              I7f9305c8bfe731300ad0a9d1ece97db4;
wire                             Ie814322ac906e4bc9baa42fef66e9b8e;
reg   [MAX_SUM_WDTH_L-1:0]       I22ace766690e445ff36176eac2473368;
reg                              I0bb61f163279dc993a94e647611f6e06;
wire                             Ic3f5c7e9a546509687973efde6a8a8f7;
reg   [MAX_SUM_WDTH_L-1:0]       I896c57162e4384f021d822789b4c01a3;
reg                              Ib5effb1b2c147179bc8c8febce7657c7;
wire                             I5a7668981b781cea8cd3de0aa6687bc1;
reg   [MAX_SUM_WDTH_L-1:0]       I3d0367a799090b3c9048235436a39063;
reg                              I81dd944eccdd3dd6fd84727d21efd0ac;
wire                             I4951067363d095f73676e08c2be255fa;
reg   [MAX_SUM_WDTH_L-1:0]       Ic0f25799f0dc7cc33de95e47ebcc083a;
reg                              I986e7c899df08e35fa2347e282e8c90e;
wire                             Ia02db0467aa519e8920344525ed30dfb;
reg   [MAX_SUM_WDTH_L-1:0]       I7186b368e297d0db1f746c6241eae65d;
reg                              Idb764022b3ae49281c7b82f6e309cca9;
wire                             I303114e80311c7f6552446bbcb0fe6a9;
reg   [MAX_SUM_WDTH_L-1:0]       I21d63f6fe5c72798aa4636527c02613d;
reg                              I311eb64d22cff4b1424f3ccdd33dec45;
wire                             I7a5c09537045dcd633095a86a6c530ed;
reg   [MAX_SUM_WDTH_L-1:0]       I15e0219f2da6f52177e76580198d0e6c;
reg                              I128183dffb32a1461db0c2b851559f68;
wire                             I6aac30f1ecc270161a81bccffab85efa;
reg   [MAX_SUM_WDTH_L-1:0]       I4cac308bee8801c4f9716673e39da4ab;
reg                              I817fbe1f44196264e2531197ca8da9ea;
wire                             I79b86b24bfa472a80487e7ea64f9dd82;
reg   [MAX_SUM_WDTH_L-1:0]       I6f4f7b4e45a495fe139955e0605ff208;
reg                              I3e74c445193a1c9ec9dcb31f4aef2117;
wire                             I208d1c07cebe2f45b25b562dd9109f7e;
reg   [MAX_SUM_WDTH_L-1:0]       I79ae5f2981b7dd91141b0a22f012f4b1;
reg                              I70f3cac8f36ef943672bbe7a9d6be5ed;
wire                             I86a3b6dc06c6c99cb1fa88023d920423;
reg   [MAX_SUM_WDTH_L-1:0]       Id4b4d757e50bc2721e8725ae10d88c9e;
reg                              I26b4d738c45246201073f4b4a786078a;
wire                             I9c0e0297c0e5042f1ed791d9d97a6f37;
reg   [MAX_SUM_WDTH_L-1:0]       I4513152c34d5d00ddcc4f099481f659d;
reg                              I6c4f341b9eeda21a97806084196421d3;
wire                             I3af891fd5da91085a79886d82e6bdf48;
reg   [MAX_SUM_WDTH_L-1:0]       I7bd4e77993fdd5a0833f1cdc7a382b56;
reg                              Ibdf325321ebd9a7baa25435537c159bb;
wire                             Ia1c63f27861c8e594f01ffb31a29ba0a;
reg   [MAX_SUM_WDTH_L-1:0]       I13b0d404e7a96cd53147b574b242ef41;
reg                              I626a4c66bf0cca36dfa2bcd8c24bff35;
wire                             I62b87c6aa6ba054ab5e80842ea738020;
reg   [MAX_SUM_WDTH_L-1:0]       I4acc3bfa99b152c6ef6d11608f639b70;
reg                              Icd6ab7be501038196ab2674cdf764453;
wire                             I429241122829d9e51a3db90b33a44ac3;
reg   [MAX_SUM_WDTH_L-1:0]       Ia1ec7ba972ec6f0049c4cf00b9d42125;
reg                              I31c6d68ecdb4d0a6790a12343f59731b;
wire                             I162416616ce392c679d22b115c192356;
reg   [MAX_SUM_WDTH_L-1:0]       I4fb5494e6f04e29d76bb8d3bc8bf6cd9;
reg                              I8eb06ffb6aca72c66cea97d9caa26f1c;
wire                             I62edec03adbb7bbda313abc2220a6a5f;
reg   [MAX_SUM_WDTH_L-1:0]       Iaffb0ef4e18bb7b582275b43684fcf3d;
reg                              I35ecf6ebd98d91d12361beef01dadfbe;
wire                             Ic3e192f5abb5526a54ea249e736702b7;
reg   [MAX_SUM_WDTH_L-1:0]       Ia5e3649f8e32a81606ee34353c54350a;
reg                              If73961b42bf31d49c78c3fbe86f8d2cb;
wire                             I1ae99cfc5ded208c2dbadbabf36fd629;
reg   [MAX_SUM_WDTH_L-1:0]       Ic675cf7eac5ece436feb5a8acd642f6b;
reg                              I560157aede2c2c3b6dce019e2fb4314c;
wire                             I1ef8bfbeda31b3dbbff053cd36de4859;
reg   [MAX_SUM_WDTH_L-1:0]       I71357943bbe307c9ae9099d4bcbff882;
reg                              I075a8e7435a4fbe97304b4d379bcfee4;
wire                             I6d76fd8af44893ab0f82a282aca12377;
reg   [MAX_SUM_WDTH_L-1:0]       Ib2684f54caebb1a1c079a2a4f2cf0dab;
reg                              I09a1ad6a0fba78d4984fee238fd95bd7;
wire                             I86247340bd399afebac1ffe403a3331e;
reg   [MAX_SUM_WDTH_L-1:0]       If19836577f9a254b365f0dcfe0ae55ce;
reg                              I5c03de756d46517f2158e4ffb019edd3;
wire                             Id932053ac235b3035e2f3d5986b7d398;
reg   [MAX_SUM_WDTH_L-1:0]       I2f47a00b58779b836c08b472d305b031;
reg                              Ia897f60b5c256180be523c5ff8ba6b77;
wire                             I4b43b5eb71dffb4bcb9ee541a537b427;
reg   [MAX_SUM_WDTH_L-1:0]       I8b2593fd0e35c37f68097187a41596e2;
reg                              I81a7d30b51b1d7f9d9bc9a97d2f3caac;
wire                             Ib481c772e0ef5d172f6b079dc8df1ae1;
reg   [MAX_SUM_WDTH_L-1:0]       Ibbcdc1c30d3333cbec65d264890cf3e5;
reg                              If46a830ca08eeb2b8b3d8b2f996491e8;
wire                             I2e046a6e848cf2da29e103872a10c26d;
reg   [MAX_SUM_WDTH_L-1:0]       Iec6e9640b0494777c013c97613855ce7;
reg                              I13e6271176ef80d03f8878441893c467;
wire                             I2a64ca51e05db642281525ccc7cf9a06;
reg   [MAX_SUM_WDTH_L-1:0]       Ic10f396b52dda0dcfbf2a847cfed617c;
reg                              Idb5b4ae9bb42a053d9db8b8c71a0b9cc;
wire                             I4275f1683058cfab72e02f2631d2ee96;
reg   [MAX_SUM_WDTH_L-1:0]       I94ebfb633f3272b8f40303ce768f0ade;
reg                              I96c6deed53888cfe0b1fcbe6832a1d61;
wire                             I592fab4d3d2c1bb3956b89eabc06dc56;
reg   [MAX_SUM_WDTH_L-1:0]       Ie975a6fd78adbad8b8a56bd6a3802e4f;
reg                              Ibb40e3b624d2f19eeccfe071e540021a;
wire                             I6520a98d1357fc57d687f9ea9a60508b;
reg   [MAX_SUM_WDTH_L-1:0]       Ib852991e38422ba6de5e18a879ddc3f9;
reg                              I93bd27a068e6fd416060bd5d919b3451;
wire                             I8a022ff37fcd6f34531af4dc7f31a223;
reg   [MAX_SUM_WDTH_L-1:0]       Ife665c9aa6794cccffd04923f4359047;
reg                              Iaf516c91fe1544bd0a6f671635eda05d;
wire                             Ia95cd411b17d1c5aaf9e5b583e9398a6;
reg   [MAX_SUM_WDTH_L-1:0]       I076cbc669ff4fb135ffc85910c888241;
reg                              I6029a024d76e9357223c6fea077501c3;
wire                             I526597e8561c75326b96e85743420a1e;
reg   [MAX_SUM_WDTH_L-1:0]       I50245c953aab8c513b17b894afb36a6c;
reg                              I8dd3c6c27d8fea2b67906c78715c5854;
wire                             If2c489abf57879ea491d9a95ce7e1cc1;
reg   [MAX_SUM_WDTH_L-1:0]       I33ac557ef59d79e8b1b359e499a00119;
reg                              I244ab0a87c282939527938b5d43c90e8;
wire                             I1dfa9cd65fb0f7c62439bc0d9539e45d;
reg   [MAX_SUM_WDTH_L-1:0]       I173fd30c1a5367b61e3fda352365f557;
reg                              I8b9861dd9f6dbeaedffc07a3e088cf49;
wire                             I5799e21b9e2fdc554f8ec65b98120544;
reg   [MAX_SUM_WDTH_L-1:0]       Id6f5041043fa4fd352e74016c4e7de48;
reg                              I71c3dc98a45a807f146ec052c8a9fb82;
wire                             Id109dde61c0ee952c9053905ee54ccd8;
reg   [MAX_SUM_WDTH_L-1:0]       I6d863254c7f0b52f803b2af4b184f99d;
reg                              Iaa6c753b09c2244d22a8680d73670deb;
wire                             Iafef3ac31f22ba4f5ef06b13165e97eb;
reg   [MAX_SUM_WDTH_L-1:0]       I1eeb9c94908cc9ddeb8e3904a145ec6e;
reg                              Id8e40a0bd35259f34ffc971eaa7f2fc5;
wire                             Ifc59d693d6dc2fa6848f37a134fbb316;
reg   [MAX_SUM_WDTH_L-1:0]       I6211e241282624fc50fb4ca1842ff9db;
reg                              I59df806ee758f4db794635ec24232ae9;
wire                             Ie83012a17bd2730837939cf0454395c3;
reg   [MAX_SUM_WDTH_L-1:0]       Iba09e22ece1eb1639d2bb940d3273fe0;
reg                              I7bd8b1c89a39e4dccbde5c5e040c162f;
wire                             I1f37257664651a57575f7ae53ab4e180;
reg   [MAX_SUM_WDTH_L-1:0]       I2fe99e4fb8c660d83508bff50ab4929b;
reg                              Id3d37273d55ba1de64f97f6d11e704d7;
wire                             Ibdf8f7dadf142fe8a166328bb5461308;
reg   [MAX_SUM_WDTH_L-1:0]       Ia73db0428763da3c0feffc94a8a8f4f1;
reg                              I4ff07696ccaf99e49d575694d3a2670e;
wire                             I0ce12cc00bd66d743ab82e89887190dc;
reg   [MAX_SUM_WDTH_L-1:0]       I6542fbca90e189048b15deaa3af5d836;
reg                              Ib89e0144bfc6be3be9a06a08e4f297ca;
wire                             I70145dd478e7f0c74c0299cdc0ab8ad5;
reg   [MAX_SUM_WDTH_L-1:0]       Ieacf022fc976bf397946d6481468d6a4;
reg                              Ife372091864d6ae9b770b69db66ff3ca;
wire                             I03d54826d217e4209d0e0f82beda4100;
reg   [MAX_SUM_WDTH_L-1:0]       I1cef7e6e0555e076b68bbc57de8f289f;
reg                              Ie81b8b84cc2795e2e92168bfa496ece4;
wire                             I0aad448f6b0692670432efdd1b92d115;
reg   [MAX_SUM_WDTH_L-1:0]       Iadaaac832a1422494d4206edee770d63;
reg                              Ia6eb1062be96666c061e5fc1f830e1d3;
wire                             Ia5a7e36b324b3a34be321ef63db22f50;
reg   [MAX_SUM_WDTH_L-1:0]       I905b0ec8983ba423798bbe8282728af8;
reg                              Ia0947c561ef360d78d0dae68baee6161;
wire                             I01399ecad74618d26fea1ef278a3125f;
reg   [MAX_SUM_WDTH_L-1:0]       Ic646b82fb6e3d0afb3a58c4e0d68f06c;
reg                              I3cd67e0abb8ff03aa1068dcb61aa3468;
wire                             Ia56986ae4171b36a362b170920663c44;
reg   [MAX_SUM_WDTH_L-1:0]       Ie57f41c62e23092974664f967a27566d;
reg                              Ic64779388389bf13a0e5240613caefc7;
wire                             I7785a1b6345c7a2086b3d2a032970fa8;
reg   [MAX_SUM_WDTH_L-1:0]       I34524ca1dddbeadcc060954238175e7f;
reg                              I767cd611a030d15fc5eebc6e1b9ea2dc;
wire                             I778c7251ca1b16e1ea1a4720ec7ba2de;
reg   [MAX_SUM_WDTH_L-1:0]       Iaf2a93993f99814321951a6bffd8bdd4;
reg                              I03e14765645af77dd39ed51320bf7a95;
wire                             I1fcb2b0e5beab6a80ce06aeca85610b6;
reg   [MAX_SUM_WDTH_L-1:0]       I97e4f7a9a8a42be813c6e4128936df3f;
reg                              I29e966dc25c12cd095c25c5e6fd6d872;
wire                             I3f8184c2f7e604f0581e5c02f5b9563b;
reg   [MAX_SUM_WDTH_L-1:0]       I682a67100f862bac0155a870cae0528c;
reg                              Ie8b68c8c51e2e03a3797a2ec3f8a56ae;
wire                             I25be48f72f47043fb6e8b7f774db1912;
reg   [MAX_SUM_WDTH_L-1:0]       Id5296b03b99bbf52d3ec04dddf3e84b1;
reg                              Ibbcfb7c284a2c99332d9261a4de199f1;
wire                             If75d53ea58491447eb2344e993b4881e;
reg   [MAX_SUM_WDTH_L-1:0]       Ibb089d47014f9002f2ea6b431156d9af;
reg                              I3e33a1f3e03bdb35d7c03f17f4ba4ebd;
wire                             I4951621739ec145bcf3004b0f72e26db;
reg   [MAX_SUM_WDTH_L-1:0]       I83496522139d35aa028dc9cb8a78d442;
reg                              I0f81337862e31b6a4a6db462533d17f3;
wire                             I959793f388e50197e4e31dae019d64f2;
reg   [MAX_SUM_WDTH_L-1:0]       Ifd4ca5a83fa0c09b043ad54d25971410;
reg                              I5029faffc78b92bc6e76d08fc4cd822f;
wire                             I8bccd3ff9583b2e33bf26d779f1c6233;
reg   [MAX_SUM_WDTH_L-1:0]       I6efbc715be55b616551a7d4650a446dd;
reg                              I11262f431003b344ab224ab5488995c2;
wire                             I177f26189ade299e79c1406cc8171ae0;
reg   [MAX_SUM_WDTH_L-1:0]       I572bf74835f5acdf5a17de2063c293fc;
reg                              I3f0fc144d868b4446b6d261b3ac80a67;
wire                             I93f3cd21e4819405b800ade59c9ccdd4;
reg   [MAX_SUM_WDTH_L-1:0]       I5f8194ef67d22bcd38f415fe8d9a6ce7;
reg                              I463736cac698d2366442abf5fba61580;
wire                             Ie655403fd0fb16aaa04783a2ff742064;
reg   [MAX_SUM_WDTH_L-1:0]       I3d3f2dff1f64ce14071e5f315bb8a57f;
reg                              I6cc14595c5c11f3ef8daa2a0b0634f73;
wire                             I1c3163e355c43d0a134c88fa671c41f3;
reg   [MAX_SUM_WDTH_L-1:0]       I8e3880fe0374bc068ed14eeff9f6d009;
reg                              Ia2345aaec32840b490d4b58c6ab3f115;
wire                             Ie378961bdb2de01ac733e765bba5eaa4;
reg   [MAX_SUM_WDTH_L-1:0]       I51d8f49653c7468b2923390dc5932a2a;
reg                              Ifdca49a87cf807777f2e460bd3d3a4fb;
wire                             Ife404037f29f17b3edcc4d1334298781;
reg   [MAX_SUM_WDTH_L-1:0]       Ibeb380f8f935c8e061fe00734675662a;
reg                              I4fab81c713b53f66f545f4f614713462;
wire                             I4109fd0e3086c344f926c4a83b378296;
reg   [MAX_SUM_WDTH_L-1:0]       I641f4280286c9343b7ce001a8b43fa21;
reg                              I1dd4557e3f4df4fa18a9198f9f36a98c;
wire                             I5d9e11667955d8128b76d9144463e59c;
reg   [MAX_SUM_WDTH_L-1:0]       I796970d7c73d8fbd7d25793d0dbf9872;
reg                              Id2ac1ca1ab4cb5eaba4ebb9dcb31d857;
wire                             I70c06d2f51ef27666c8c39e0a13ff5cb;
reg   [MAX_SUM_WDTH_L-1:0]       Ied0b1d10ae09c523d1cd1cd3e5b184c6;
reg                              Id40872fc0d4f1e9ce25d366069af2f1a;
wire                             Iacd270f7fbb94c91757a4f8780616e1e;
reg   [MAX_SUM_WDTH_L-1:0]       I7d0d39d94d929741158c39f69e8169e4;
reg                              If3b1c8b7c2296e5664f105adc761fd48;
wire                             Ia95e1a8c5bce4673824d56d6fab81f4b;
reg   [MAX_SUM_WDTH_L-1:0]       I2349636f6ea8796c7b798aa555641a9e;
reg                              Idd694db68c0f91155fd81a106d596d8c;
wire                             I49137af52922e3872901905fd7c70601;
reg   [MAX_SUM_WDTH_L-1:0]       Ia3739201eb91605fc115bf320d4c24f0;
reg                              I89473d1b100eb64c951e986819a4bc59;
wire                             I548d9239de9b536e1b581327961b53df;
reg   [MAX_SUM_WDTH_L-1:0]       Ic74cc511acc98510da011e126edaf3a3;
reg                              I4351f5987566977330a1e69b78d4e6aa;
wire                             Ifad4cf6d79d76caa33927ba4a6b94b45;
reg   [MAX_SUM_WDTH_L-1:0]       I89b1312c0696711956ddcf787e37f3c9;
reg                              Ic067d44971ef80f6c63c6e187a583e3e;
wire                             Ie78dd544469009d2b182d2b76694df6a;
reg   [MAX_SUM_WDTH_L-1:0]       Ib2ef1187c1743da2cd83eb9231a7ddf1;
reg                              I9d46fd2fca52ea2ecb6242801a4378a3;
wire                             I69122b791a8f717c501f2842240a51f6;
reg   [MAX_SUM_WDTH_L-1:0]       I21710bdb6874ab83e2b2a2cffb026ab8;
reg                              I916104565afa11bfd9b3ef53551ade1d;
wire                             Ib89ed0cfe4ba481ae28b835d4248babf;
reg   [MAX_SUM_WDTH_L-1:0]       I2ec8afd22c84596550412a5d2c7129af;
reg                              I48812dfaa796a851f23d230227be8969;
wire                             I6ec25bbba8c41ebdf4efa95fc1d8e1b0;
reg   [MAX_SUM_WDTH_L-1:0]       I57056cc2fd4bd1ea6e980cf90c22e871;
reg                              Ia2d3db44f16c9bf381145ce71ba2efd2;
wire                             I92953d645060c118de19fafee18e34a1;
reg   [MAX_SUM_WDTH_L-1:0]       I233becd31032d63e65371119edb2cf79;
reg                              I849110a991c42aefaead8d9500a18912;
wire                             Id89c23eca2ed6103c87dc296082605ab;
reg   [MAX_SUM_WDTH_L-1:0]       I0142623400f5994f581a4797fd9d327c;
reg                              Ic4988fc07458064e44f882807bd13c4b;
wire                             I070e631601f2529f8f18ad0be6a70316;
reg   [MAX_SUM_WDTH_L-1:0]       Id3e298c9f2709d8dc01c18626ea846e8;
reg                              I0fdd344f1ce42003661bb06c2c0d2fb5;
wire                             Ie1e3e5fbe2e2ae4cb3218616bcaa0ae1;
reg   [MAX_SUM_WDTH_L-1:0]       I1044e090bdf84a1bd30438137d6ed056;
reg                              Ib2ab217127041c49acfc86ef2eba3350;
wire                             I6b2795593e93e47b2733c1e0003a7806;
reg   [MAX_SUM_WDTH_L-1:0]       Iff0f43c1fb40bdb3271a3a38d89f4d6d;
reg                              I5d6dfd14a38b207a97ba02a357965d5e;
wire                             I467646a701c26d253f43251aceac9527;
reg   [MAX_SUM_WDTH_L-1:0]       Ibc71a0c3641097c144513810bc9a0a7c;
reg                              I963472efe41928bdcd4c87ae5d6d9781;
wire                             I280a8abed1540ebaf599c094a0a75797;
reg   [MAX_SUM_WDTH_L-1:0]       I6ef3b025eb065f833efe6daaab699efb;
reg                              Id8cde19539c6cdf7186230e34b96dc15;
wire                             If75560cad0cb26bd315f3711d1e9711d;
reg   [MAX_SUM_WDTH_L-1:0]       If76152e9435e7300b19095a9b070e0f4;
reg                              Ia31ee8ac9735d3bd38298fd5d9812aa1;
wire                             Id0d79e0b7361bae1b007c8a7d606f6fb;
reg   [MAX_SUM_WDTH_L-1:0]       I5fa63303ab85db9c8cd268528eb604ca;
reg                              I79bced0e80e2554a4e748644c5985896;
wire                             Iac7bb2fe5935b53852a63923c53f13a1;
reg   [MAX_SUM_WDTH_L-1:0]       I69d6adcd3d35a24b393e97ed6a99c061;
reg                              Id0216555323efdec39d0448568f59f23;
wire                             I4554a553586d9966e7d4e8d99a5c799d;
reg   [MAX_SUM_WDTH_L-1:0]       I8980eca0e5973840121576b6eaaab736;
reg                              I35c6735d2fa06f57341b6010f5bb825d;
wire                             I84a85d995e807610f153e72ea3df3ae0;
reg   [MAX_SUM_WDTH_L-1:0]       Iadbb5c4f7b7c02e151d5118a7ede1f0b;
reg                              Id2e8b17327e8c85999d3d6b3dd31a164;
wire                             Ic68f898ba0d0073df41bbfae0944c9de;
reg   [MAX_SUM_WDTH_L-1:0]       Ifff90bff22a3bcc33261004136d2e655;
reg                              Iccd9ca809045617acea3364a6c86fde9;
wire                             Iab98e00ea4dca63c81eb8f78a133b1bd;
reg   [MAX_SUM_WDTH_L-1:0]       I8d13628f322640414a4b556ee48d3bdd;
reg                              I8ce27f01f84ea9babfca8074bb57417a;
wire                             I67aca5b07f66a9f3e8a5550020802c63;
reg   [MAX_SUM_WDTH_L-1:0]       If7d187cc56b1014b1582c5f5b94759f1;
reg                              If6bad1b3865cb4cec97a730043863b3d;
wire                             Id4b0e0110bcd34cf8f0a9a92108b88c2;
reg   [MAX_SUM_WDTH_L-1:0]       Ia01d5a33078abf4b2d6c625af01c25f6;
reg                              I0c88089ad1c5fc9928c091c1c677ca66;
wire                             I29ee6514004941d4280cf4a93e7baf5d;
reg   [MAX_SUM_WDTH_L-1:0]       I4c74240688b5635b5323ce3a8ac666fb;
reg                              Ida2ed38c156200b9511c3b4515f42e5e;
wire                             I3bb0ea6e5c41271be14ed45d4b8ece5b;
reg   [MAX_SUM_WDTH_L-1:0]       I943e9afa0dc80fb50b5869cf34726823;
reg                              Id322e4a2b0197e5b0f67a220134ca540;
wire                             I0a1dc75c36d5fb043c80dde4e8c5e577;
reg   [MAX_SUM_WDTH_L-1:0]       I44d8779f30245bc7f1475e6feb762cec;
reg                              I935862d2f7c82e05768f55434167ba47;
wire                             I89e39167f230c52eaf64e8c5ce8fc38d;
reg   [MAX_SUM_WDTH_L-1:0]       I479e7456c445ad604ebc134872a0fbfa;
reg                              I1c6dd243cd7d2b8d00eb59e2ae30331c;
wire                             Id6e88b1c05e5f4e7188f4b646f428b55;
reg   [MAX_SUM_WDTH_L-1:0]       I484f372e3a2e74e0791b06aa666b781e;
reg                              I8ab7b4e7f78fa63ec77224c7e5a31198;
wire                             Id9b024743e4060a62c6dde2646b5c998;
reg   [MAX_SUM_WDTH_L-1:0]       I64b07241996c48963595f28e35a75be5;
reg                              If20d6cdf73bb1a925317f35de01b6f62;
wire                             I2bc4cf6682dca441749b95f63592dd8e;
reg   [MAX_SUM_WDTH_L-1:0]       Idf678798bf4e1cd316a49a2b413cb29f;
reg                              I8c2bc7a3c5c7e798a9dbd0199d37bfd5;
wire                             I05d8735777c75ecc9f1e5d2f972f5c21;
reg   [MAX_SUM_WDTH_L-1:0]       I35fd5e5e93f992ef5ff6b11f9d69609c;
reg                              If814b033c7e3229ba1475b305fe98307;
wire                             Iaa201a0537ab3cbcb5bc065871e0153b;
reg   [MAX_SUM_WDTH_L-1:0]       Ie72397edc1c597c0a8213b67a030a482;
reg                              I6e69f6d33a933441458f5a46decc4e8d;
wire                             Ib76deffcb8cd38d5643df9447f3b060b;
reg   [MAX_SUM_WDTH_L-1:0]       Iae50178e99a07cee0eea6f7cfdcedf1f;
reg                              Ie2bb4ef41cf43cbea46b7a6d492bf03b;
wire                             I6483a59c7f2bc77b445b202f0448eb2a;
reg   [MAX_SUM_WDTH_L-1:0]       Idd7082c7a65d7f8e0ea88142312a631e;
reg                              I757b0e2104a4d9913cf6b3a13ad7d6d6;
wire                             Ic1ffdfe961dc8458b1d4cb36642a386a;
reg   [MAX_SUM_WDTH_L-1:0]       I4b580dc4cfac9e9315d03b60e2a915d9;
reg                              I46c7f4a6ef4b3ac3eb74b4ba2552fcdd;
wire                             I0fb493a1f8f2810ddf67a6cbcb2c782c;
reg   [MAX_SUM_WDTH_L-1:0]       I77cdc9841414221c3f6c3cf35397059f;
reg                              I247479fee56f209f758feeb4770e50de;
wire                             I2c555af9585a50d2cd6a27c223c8722c;
reg   [MAX_SUM_WDTH_L-1:0]       Ie59619c3e78e616e1febd2db2fa940ae;
reg                              I2ada4b104b94c163f3d9201808d21121;
wire                             I5f93af2953a9f1aea5cf55a037f7af6e;
reg   [MAX_SUM_WDTH_L-1:0]       I5bc8079a5896f59bc6137b59c4b7e750;
reg                              Ic7f0721d5160d4ce266b21c53aad0b4e;
wire                             I25b3e2b9f55ea811784ba8ad8c5f516d;
reg   [MAX_SUM_WDTH_L-1:0]       I239bf978d991f702ad23bc6b4b8be1dc;
reg                              I9af70dd16bd606c4b9588ce32ce9844d;
wire                             I93fb55e460d75b8d36c19833849bc1d2;
reg   [MAX_SUM_WDTH_L-1:0]       I450351fbb31246b49cfb2d622b9e90b4;
reg                              I30c5fca5bab3bc9cf5c024c3302bbdbd;
wire                             Ic51082943371a401c48202b4e655e84c;
reg   [MAX_SUM_WDTH_L-1:0]       Ia7c17a0979f3bbb9e9e821bf69a239b7;
reg                              I09db79951c2115c2db0a3036bcb2b63f;
wire                             Ib53122ae54dc4ac5b090ba8aa3ab9959;
reg   [MAX_SUM_WDTH_L-1:0]       Ic22975c34b92a39bc8940076e80d3c0b;
reg                              Id76636b29db2c1a69d585b68731fc3b0;
wire                             I459abcd025ce92565cbbfaada735a325;
reg   [MAX_SUM_WDTH_L-1:0]       Ia7be8cf38ecee4568a939cb2ef727619;
reg                              I2ce42f5733f4d0cf15d1a7944fe0344f;
wire                             If8abbbaf2986196395e63aa49b1022bb;
reg   [MAX_SUM_WDTH_L-1:0]       I3e475cb1733d494f5f7c4b26a07d5852;
reg                              I87e7191f5ec3f0847afbca81660a7608;
wire                             I830ffb778558295001c003f114b66198;
reg   [MAX_SUM_WDTH_L-1:0]       Ib2c0df16678f6aac19f7af4ad4e53ef8;
reg                              I0f8f4304c88efcc90c021be7764be01b;
wire                             I56e732494aa029b716ac04289d951e27;
reg   [MAX_SUM_WDTH_L-1:0]       I8bd2ef39eeb7089409db02e3806956ac;
reg                              Ie8b6b834bdde210d6f7a3e60fc78275d;
wire                             Id077045b00947ff1b4de86777d84a48f;
reg   [MAX_SUM_WDTH_L-1:0]       Ie3669e34cd19462f524932b3d232b546;
reg                              I591b99ab1b55e2eb4c10996efab5e0d0;
wire                             I7ce7ba4f90dea6eb91d61cb456134df3;
reg   [MAX_SUM_WDTH_L-1:0]       I1ecea23a4e56948365dcb04c5bf6d6d6;
reg                              I27402f7d7892626f9b5ea1fc39987c23;
wire                             Iaee8dd8470306340982baafd8c9e28b5;
reg   [MAX_SUM_WDTH_L-1:0]       Iac222e9e39e300d7161ed05153cd9ca0;
reg                              Ie6e9475310530f511d38602f2c58a28f;
wire                             I35088305c303ace3b0bd194f5efa557f;
reg   [MAX_SUM_WDTH_L-1:0]       I292683f8453be58f65370a286c1a4505;
reg                              I30eeb2d396c381acb08253d886025fe1;
wire                             If28f074339d099d0c8f0e582c11f57e8;
reg   [MAX_SUM_WDTH_L-1:0]       I1dff7459553fccefc94a6020cc248a49;
reg                              I9a9a3b834bb25862cbe40375e20c2163;
wire                             I55b6efd25a905ab958ff62e0334d0116;
reg   [MAX_SUM_WDTH_L-1:0]       I9acec7aa4b420b7c820028b669a8bfb4;
reg                              I1152ba49a018ec527bb8091c0cebd737;
wire                             I859a2864cbe2fffc01b411e7b0a2c3d0;
reg   [MAX_SUM_WDTH_L-1:0]       I714b7d8b39c4135183b605dd97ff15d6;
reg                              I1cf3b72b3aa02961788688172c1ad2b2;
wire                             I3ede6ae83cec11aecdb308142c26f6d6;
reg   [MAX_SUM_WDTH_L-1:0]       Ie5856c36d9a310f890ecc5220590fc3e;
reg                              I09293a7f47ffb53331aad25a876d2562;
wire                             Icb7fa4f4271f536afd96934a45bbf0ff;
reg   [MAX_SUM_WDTH_L-1:0]       I062b1d8d3b6fe6d8e158ede1f0af9eed;
reg                              Ic00d9c70df8f473695a4aa76827ef690;
wire                             I4dfd9e0bf539f3077f2d5a8bd3b5e469;
reg   [MAX_SUM_WDTH_L-1:0]       I0fbd5b5eef6da9adaf918390f6bdbc27;
reg                              I36132477ed96c4731e46d24e9ca1e9e8;
wire                             I795091257b4f78363310623b731b347e;
reg   [MAX_SUM_WDTH_L-1:0]       I73fb14b30841cf67e96ba329fdfa3e35;
reg                              I2cb80c174e5ddbbaca6eabbfa7c669c7;
wire                             I6ff1f76a6ad568b5fa0cb300a67ceea9;
reg   [MAX_SUM_WDTH_L-1:0]       I6d6cfca51988c5ac32471fe8f4399bbc;
reg                              I359e17e055d03931cac7b41c77be575b;
wire                             I5864383518b7c9a70f69b0fd1a64d4aa;
reg   [MAX_SUM_WDTH_L-1:0]       Id7940e4951c96c3de9f45119043fbffd;
reg                              If466ac9d4d278b49b4aa91650b30ec2e;
wire                             I30959187f5ac883ab77af90ccfce5704;
reg   [MAX_SUM_WDTH_L-1:0]       Iea71361c5f846419eaa18ae4b9463ee8;
reg                              I17d171b83e60410ce78a7e4fa9d17001;
wire                             I0d2bcd2e24e64ad5703a580ddc415f3a;
reg   [MAX_SUM_WDTH_L-1:0]       Ib67ac5fdd6e068ee799965b51aa893ba;
reg                              Id79a4b98545d81fef573054b93ae80d4;
wire                             I4d1ef379c32f93cdd18e2415ba83a5ea;
reg   [MAX_SUM_WDTH_L-1:0]       I0bd84509dde112f3657bd5a12a8df72c;
reg                              I4e8f5e83e32143008d70a8edf17e2ff5;
wire                             I921c8abbe15effa3769c5c3f81427274;
reg   [MAX_SUM_WDTH_L-1:0]       I2caf86026460a024f752fa71b44f743f;
reg                              I57cf1069290a2a5f30b75eb592752b88;
wire                             I40cce0292c07026fb144dc28ba228485;
reg   [MAX_SUM_WDTH_L-1:0]       Id81d9c9ffa81c2653dea2e872ab2f71c;
reg                              I7447d4584dccf4dac9f0d359748ae327;
wire                             Ia1401fc86b9d014a28f1c5bfa7aefc2d;
reg   [MAX_SUM_WDTH_L-1:0]       I0b4d1a08307d452870c3e762bd038568;
reg                              Ic4571481454a10eb7f8c0b58f9d35178;
wire                             Id3899a9a35b467c103ed0dfef20dd4a1;
reg   [MAX_SUM_WDTH_L-1:0]       Id75cc40233cc8648e21a750d882d5ed4;
reg                              I00810b2849a3d3097e028efac18c0a06;
wire                             Icff78887751d68045a0bc21e69047c79;
reg   [MAX_SUM_WDTH_L-1:0]       I3ea9815ba887e373a0a477654f136856;
reg                              I19be1cf97631f5bd782d8358fb55954b;
wire                             I9a2e36db1aa972536df63a24462eba98;
reg   [MAX_SUM_WDTH_L-1:0]       I8b26e270c3ca5563da39e7092ef830dc;
reg                              Id7fe36cc9d5c1d7cc54ee1040e6578de;
wire                             Id74033401d8494d013fcfd1f69537592;
reg   [MAX_SUM_WDTH_L-1:0]       Ib03f94d7e5ff830d5063cd514e7f7998;
reg                              If6984aadfa0583c3281a04ba48f3d765;
wire                             Ib64741c15a5f128b008851c36d55c0ca;
reg   [MAX_SUM_WDTH_L-1:0]       I00b05bb0b225b27562d6629725ac2126;
reg                              Ia7750161c32ac0507e1ff6a8fe896148;
wire                             Ie75e57f87e9c8cc7d29519f0419f1b22;
reg   [MAX_SUM_WDTH_L-1:0]       I1f273682cac5644f1fcc30ffa20f8cd8;
reg                              I97d6084735a682ba654fc70a9e07f27d;
wire                             I95bc08d218c4a924f810b69c7e2b923f;
reg   [MAX_SUM_WDTH_L-1:0]       I483725645504999df82a4d0660873c1d;
reg                              I3e9d85c0ca08314fe2da0fa6977942b7;
wire                             I6dd9a12bbad2fd4aded0354fbb09c6cb;
reg   [MAX_SUM_WDTH_L-1:0]       I689dc18b56442b8db01bd7ca4c44d615;
reg                              Id28d0dd03217797390811bdd3564191b;
wire                             Ie78ca77c4a9cfac31f52cc1f49e5c6d1;
reg   [MAX_SUM_WDTH_L-1:0]       I805d665f394ff24f230bebfa6d252122;
reg                              I0eb20560e7e211b67cfa8ca9e056c1da;
wire                             I771cf2bb35d06a6009955936e2530f07;
reg   [MAX_SUM_WDTH_L-1:0]       Icfba3f165f1cdf2e6070239100e9ac3d;
reg                              Id089d9523253f91c670099157325af05;
wire                             I2d9d14b5c585e74db793171f304e5d61;
reg   [MAX_SUM_WDTH_L-1:0]       I93c51f71db0e3df7f6e2978fd93fbb54;
reg                              I4db3f0e5ff2cc72e499ab5f1b9fd1d14;
wire                             I1e7165374d01b2b7abb1e1883daa4463;
reg   [MAX_SUM_WDTH_L-1:0]       Ib7410e44d23eea21613074695b64bd2b;
reg                              I082972cc68873126a258e9db29e524f9;
wire                             I783fdf0d5058b09d9d0d5c87d9926c50;
reg   [MAX_SUM_WDTH_L-1:0]       I93cc273684a376d76a2e3468b3dc8bd7;
reg                              I3ba1cbc9ff352842d6d687b2218b6c0f;
wire                             I1c66ca0e94ab96e8420e97641a5a707b;
reg   [MAX_SUM_WDTH_L-1:0]       Id133dc3fa65840136b1157fe97a1e962;
reg                              Id8fbc7f9a403b07efd27c20d6d78e661;
wire                             If5f2d3751eb3af97e20c680475976bb6;
reg   [MAX_SUM_WDTH_L-1:0]       Ib792104b6cf946d632f7591f2cd5e104;
reg                              I0628944b437e239b25736381fa59901d;
wire                             I96f91ace9649929071ca3e6e87eda861;
reg   [MAX_SUM_WDTH_L-1:0]       Ia44bcc8308360d3e6fa351bc108df3fa;
reg                              Icf6bf0aab709fb68c18e26f9fe7503b7;
wire                             I27968f9d2e9dc75bfa55b1e5ad6f8c8e;
reg   [MAX_SUM_WDTH_L-1:0]       Ib29a26c41a3ba089efd30c3256106a7c;
reg                              I15947ee18296366e3e13cc9727ad2ebb;
wire                             Id53e488ea1a69e9d1e50dc276c14bb43;
reg   [MAX_SUM_WDTH_L-1:0]       I8999f385aaf15b67e4c12e56c7dba7cc;
reg                              I23b16e4f6f2fab529ae42009d38cee85;
wire                             I8440ba68619a5a3aad3510ad6ecaaea6;
reg   [MAX_SUM_WDTH_L-1:0]       I202980f6263e3b312c38061224992740;
reg                              I51e128a639866ca032029880ae59e874;
wire                             I9e00e6e111b313b2efd5c9d32eae6a8e;
reg   [MAX_SUM_WDTH_L-1:0]       I1fd9ed3763ff0ce0a671360f83bc3613;
reg                              Ib14c75f869e8f09519517f3fcbdfaa7b;
wire                             I1836b01cfa5570153a8e4387baee29d6;
reg   [MAX_SUM_WDTH_L-1:0]       I4b58194aa6a5b5c825f14bb926a0ae9f;
reg                              I9ceea65912b0a100eaa0afb42e84e5bd;
wire                             Icad06a6e006badf38d87cd3c4fd0981a;
reg   [MAX_SUM_WDTH_L-1:0]       I706daad77f6a6eddf5576c238fa4714d;
reg                              Id93be78cd06b38e1d7ec35ee66f878c3;
wire                             I8c061e6f5fb7e2be23d69254f0d0f59c;
reg   [MAX_SUM_WDTH_L-1:0]       Ibceceead1cdcf8805e9a9f93b3b783ca;
reg                              Ia61e18c0042f8ec7abb670e7f0648b45;
wire                             I5411a76d49de45984ac852d98159ef5d;
reg   [MAX_SUM_WDTH_L-1:0]       Ia5956c899daaaa0b2b0c16f524feaf98;
reg                              I117b1ef192f2b24c6764c2d96864cc5f;
wire                             I826369ad5207f64f64ff58abdb9f321e;
reg   [MAX_SUM_WDTH_L-1:0]       I7f353333180ccbf6a271c9745430b199;
reg                              If5224b5f45318dac2a64dcc72c6afad1;
wire                             I4c266cd72fd1cd92f21511071a51c361;
reg   [MAX_SUM_WDTH_L-1:0]       I958f0106e3ffe429d0450f4b6e9ada3d;
reg                              I41710bb2545ba34f65e6d9a24086185b;
wire                             I76aac239cb31a0bdcebd7a3e3829f274;
reg   [MAX_SUM_WDTH_L-1:0]       Idf02454b4aacb6ff03288bb19a4771b1;
reg                              I15a9f9397a5d23e6885ac887723a8a19;
wire                             Ief0092617ed13bebb791c57c0da0b12e;
reg   [MAX_SUM_WDTH_L-1:0]       I42f39cecfe5c3d77b3fffb624cdb2c0b;
reg                              I46f40fec14e2e6d5060c97f0a0d86696;
wire                             If1a6e0ead8f7aec9046bf22a1f59cf68;
reg   [MAX_SUM_WDTH_L-1:0]       Id7b0871cafd2630ba4dfc3e058613908;
reg                              I06e512c9097f76687d65c87f99c74764;
wire                             I26ee3d378528d4a8469eee34a7b5652e;
reg   [MAX_SUM_WDTH_L-1:0]       I18c1c4d71799c5da8172f6cc63d2d37f;
reg                              I17759c97920685cd28c898441838531b;
wire                             Ic8f3b5e177f927b64f1213625abc76c2;
reg   [MAX_SUM_WDTH_L-1:0]       I7d53f3ce487b0a2446d5205868c29175;
reg                              Ie7da1180f2c4eb8153421db4c6317a50;
wire                             Ia813a2600edc508e2eb59a9856e8fc4f;
reg   [MAX_SUM_WDTH_L-1:0]       I37fb9120bfe27a0e7449583dda735479;
reg                              Ie6fe42c4fa7e64067960cab4edee83d5;
wire                             Id04ad2fc64d6c346ae479abcbf3df41a;
reg   [MAX_SUM_WDTH_L-1:0]       Ie7e15e6743a750cbf1b272da694b47dd;
reg                              Ic064e5425fd7a36be5860a40bc765994;
wire                             I2827f1757a4ffc394869610f710291c4;
reg   [MAX_SUM_WDTH_L-1:0]       I66a1e62b25bce18e36d78c382b40b1df;
reg                              Ifc8326ba561071589aec67a7de4276fb;
wire                             Ic8c6fbb1e7408869e5d11d0aea83203b;
reg   [MAX_SUM_WDTH_L-1:0]       I9b81ec12daf51cb61f7dc0b9ad01cc1d;
reg                              Ibc55f69c8c895e9fad768b4b1a4a7a20;
wire                             Ibe0134da146c0c96af213013c5215943;
reg   [MAX_SUM_WDTH_L-1:0]       I9d76cb6c99a69086774f7fd471dadf53;
reg                              I50b89d077d160ee7d56376ae0abd9c6a;
wire                             I46a2e76ccab8ae201f78845054028074;
reg   [MAX_SUM_WDTH_L-1:0]       I4c59798356c8e05f8b2cdb4e202fc4bb;
reg                              I59a2c5b8dc1924b8503c24efa60c0c4a;
wire                             I1ee771cad3766a589cd62746062401c4;
reg   [MAX_SUM_WDTH_L-1:0]       I395b43b11730131a5f4331b2ce82717d;
reg                              I57a7c62f6cdf0fa0bd65df83a4904e36;
wire                             Ic37d0375083a9415f7c0e9650ef0ecb7;
reg   [MAX_SUM_WDTH_L-1:0]       Ib3f07793c2e2cf7b6ac988be01a55829;
reg                              I733e71d48b2ae728b9d7b6a86261a156;
wire                             I73167dd9e24b49f6af3f7493cc2f9c0f;
reg   [MAX_SUM_WDTH_L-1:0]       I05ad19dc723fe482f93cb524c8c86cf6;
reg                              I20386e26c247b478dd7f2c89e73a1016;
wire                             I156970479a68c248bffd30be0097ff8f;
reg   [MAX_SUM_WDTH_L-1:0]       I1db8d47c1852578aa6325919279419b1;
reg                              Iaa6dcd47c9356b0b3b93d83f87c7fa05;
wire                             I851f4bdd95d1297f7ff05f01830c93fe;
reg   [MAX_SUM_WDTH_L-1:0]       I98ec1bdbb599febfcdc06dbf807ab781;
reg                              I8913043709d09e66411b5e70b0e3c969;
wire                             If6f8ef7f0cc4860dfb264b645ab0898f;
reg   [MAX_SUM_WDTH_L-1:0]       I86f73b27c90bbd800b521fb8953d5506;
reg                              Ifdcd9ff3c567f73e0366261dd09dee05;
wire                             I5b983a4c1b35218893ed1bb0aaae26c8;
reg   [MAX_SUM_WDTH_L-1:0]       Id117870de7302febd51da982ab8b524e;
reg                              I95af25eeba42e7fb3dc0dff9b702f61e;
wire                             Ifd281eb29091bcaf3a2929983366e637;
reg   [MAX_SUM_WDTH_L-1:0]       I6cff1d82f4c1bf7789e39b964dd9e6fe;
reg                              Idf7fd041b837ee19551784f305c4efa1;
wire                             I5ef5030a4e29e5e3c981d2616cae1ccd;
reg   [MAX_SUM_WDTH_L-1:0]       I5d9786c9b4566669e7981654c3c10da7;
reg                              Ida9601d0e04fcfa1e448b681c4aa6bdc;
wire                             I3051150debf8f223b936ea5f169623f8;
reg   [MAX_SUM_WDTH_L-1:0]       I83dd9071e7e35d7165d556a67d2d1658;
reg                              Ibf6735fa3cd381ba501ab67979729a08;
wire                             I9b76f1b49c0faf3f89256a1fe04c4597;
reg   [MAX_SUM_WDTH_L-1:0]       Id62c5db9d4a4e5eb91ca4b6876d36a9d;
reg                              Ic78e2d18e11538916e6726418f181e48;
wire                             I62626dac5bf648ffad6e6e3cd836ab9c;
reg   [MAX_SUM_WDTH_L-1:0]       Ibeb5414f37bbb8176c1a9ac51957dba0;
reg                              I4b62c23b8d6b70c44af359b951424df1;
wire                             Ic527dbbf40cb847b5e5400f177a635da;
reg   [MAX_SUM_WDTH_L-1:0]       If40561e9d6ab97e7dc2c6eca6d0725d8;
reg                              If6467cc6d4b393b76586f5b65ace1435;
wire                             I44683db6537a0ae1bfdca8b6448c3772;
reg   [MAX_SUM_WDTH_L-1:0]       I630618151200231dda94b3fb59a24829;
reg                              I1e79f24aac8988678a3ac91e9dfa493c;
wire                             I5a03f223dea2bc87a454b29c3fe6058b;
reg   [MAX_SUM_WDTH_L-1:0]       I45948c2ccae2bd2c2fcfe9c75787e2b4;
reg                              Ie3e87c23a6fbd77afb7a98ba764d937c;
wire                             I8a7824d737ac024ffd25428f6599c070;
reg   [MAX_SUM_WDTH_L-1:0]       I73048e349b470dbb16b2b3e69aebcb3f;
reg                              I6406707a5545040df609c67f677e983d;
wire                             Ia7e5724b4f05b0b6bdedaf264e797855;
reg   [MAX_SUM_WDTH_L-1:0]       Ic3a706eeb522f64147d4946983a9fcb4;
reg                              I6aacacd072438b5172d5bd0be77c9ff8;
wire                             Ic8d1cb210627d8d6e717625ad3dd0fbe;
reg   [MAX_SUM_WDTH_L-1:0]       Id8934e8818877e81d701105823366043;
reg                              Ifea8a5d86f6681180539911cf637e785;
wire                             I313adb9858a6a31cce5af3d108459bb8;
reg   [MAX_SUM_WDTH_L-1:0]       Id5fd5653bfa014fa0e956ef4b1d83291;
reg                              I8101cabc2e8401f77a50d561a53b385f;
wire                             I36dd39ffe6e62b2518e12bb8e544ac20;
reg   [MAX_SUM_WDTH_L-1:0]       I41821f6b5a613fde6539e41a6a0c7b65;
reg                              I9574b260963de729540209c0138de41c;
wire                             I94337aa2c4ca0ec7a962962780f21f11;
reg   [MAX_SUM_WDTH_L-1:0]       Ie8d437ed136f7f5971638d1f62ffdf15;
reg                              I791728546a36e98c0d5c4eb1063082b3;
wire                             Ib2443922534953e49e1af5343c028fc6;
reg   [MAX_SUM_WDTH_L-1:0]       Iaf46eedc430b55905d73486ac0752c8f;
reg                              I338183bc2bdb39e2a3820a768d78ebdc;
wire                             I08d6c121fbd306f3908a88ce10779ac5;
reg   [MAX_SUM_WDTH_L-1:0]       I32671ef3896bd0b586f13c092dd04b9e;
reg                              I4197bb0d6d0465aeb6fd7f0a8189a368;
wire                             I1b947b03d2db27afe8faf78f580c90aa;
reg   [MAX_SUM_WDTH_L-1:0]       Ie8bfdf207d647c9f161bdf265a8472b4;
reg                              I8f0d7e1f97b611f6c4a231338aaba68e;
wire                             I05b4915602c4c635f9e91ff69432ebf2;
reg   [MAX_SUM_WDTH_L-1:0]       Id44fe933294cafff88d133a0ddc1a832;
reg                              Ie50a86c3b69d3884c72948133083e099;
wire                             Ifdd87b92e70f345ca64fa4e96d732210;
reg   [MAX_SUM_WDTH_L-1:0]       I20c1f8e56a14db0665160ecbb277fb1a;
reg                              I2cf91b227a82701d912cf9e9e1040ddc;
wire                             I67335037a5b54e1b5bb316cd3519e790;
reg   [MAX_SUM_WDTH_L-1:0]       I7627f96e870f6a3e8abd7ac494bc178c;
reg                              I0f50e2edf3586292da17ce7214d37038;
wire                             Ic0feb7035ff8f8962a79aa20f4129bbe;
reg   [MAX_SUM_WDTH_L-1:0]       Ia2d3997dce108f85ed64e88780e99efa;
reg                              Id7666dd5135e45a1e42f13ffbb8558ed;
wire                             If11c3d720e491cfc18684f3a23f6b93b;
reg   [MAX_SUM_WDTH_L-1:0]       I6a25dc88186816258f1237123ee4968f;
reg                              I3dbcf0199e35f410c38ab3d9e2cac2ef;
wire                             I5d4a36427e26532bca590796e4107dcc;
reg   [MAX_SUM_WDTH_L-1:0]       Ia9d61848b5384a8cc63321201174f3d3;
reg                              I06c6db30fc7e63facd144d0166702e6a;
wire                             Ib0eb8c6ddbbcd4825e8fc5b1c55495b3;
reg   [MAX_SUM_WDTH_L-1:0]       I53ed79856aae53b180f28b47822e89b6;
reg                              Id20d5070afe5748b50833f0593777c49;
wire                             I0d5ab203120026f15a1d563bb65fa1ab;
reg   [MAX_SUM_WDTH_L-1:0]       I76503bcb779e039edc9acfc03a2d1ee6;
reg                              I3d041f7cf6c679d8d9677445eac96640;
wire                             I35ca485dc9ef601029877a4ee46ed942;
reg   [MAX_SUM_WDTH_L-1:0]       I18ae85d6725cf0ab3b69bedeef651425;
reg                              I51d27603f0a87b78857b8e064182d925;
wire                             I8c1c4b4851ed06bce6af5b392c75c6b8;
reg   [MAX_SUM_WDTH_L-1:0]       Iaa3bbfc6704e70a55b8e1083c326820f;
reg                              I9b6d48e71d050b9b0b5c5e7407288103;
wire                             I00fc4e266ce9e790501c78809bfae38e;
reg   [MAX_SUM_WDTH_L-1:0]       I8c1c3ee4b57d56ab362672dfeb4e0ae9;
reg                              Id05706fe9e0fc4776e0446aacd4c118d;
wire                             I35fa53ff8ca5fab19b6de45beda84ff2;
reg   [MAX_SUM_WDTH_L-1:0]       Ic8e0765b1cf95f2578a7ec656d027f6e;
reg                              I2ec61e0e1b707857ca39f532bf970e03;
wire                             If3c4067202f592fabf77cd76db5575dd;
reg   [MAX_SUM_WDTH_L-1:0]       I39eaefaae486119c8741c5e9b7f85bd3;
reg                              Ibd1b4a1010823cc9e4a78a0fcefd7d01;
wire                             I64276a920c9ccf7576c15618812fd152;
reg   [MAX_SUM_WDTH_L-1:0]       I6ac8d8000e434fcca222525ac00f9849;
reg                              I6da2861072f65e35d46d224b982eda7a;
wire                             I478a999d16ad8a5266769d1b8caa79db;
reg   [MAX_SUM_WDTH_L-1:0]       I114cfd3fe8f5db92b879e0dce592af3b;
reg                              I860c7e185d38d907c4ed20a64d238dd6;
wire                             I29f2854aec43820204ceb8f3eceed6c9;
reg   [MAX_SUM_WDTH_L-1:0]       I8db1c7f6b5c7c04f71e7fcc18f7b9941;
reg                              I76e06fe466c43e4aef0ef860f0274fa8;
wire                             Idf664119a34b4692c0cfaa4c742480f4;
reg   [MAX_SUM_WDTH_L-1:0]       I89e516738a408ccbd495e4f5aeeb38a6;
reg                              I3c00d8a5dd8c99ee527ad4180e469ab7;
wire                             Iae32c64d9bf268ccacaec2d40efe70f4;
reg   [MAX_SUM_WDTH_L-1:0]       I0c02b9318bc4f50969f8d486e587a627;
reg                              Iba2018bad14888e510fc7f4a4e040ed5;
wire                             If30e09a7c080fd91758eacb33912b8d6;
reg   [MAX_SUM_WDTH_L-1:0]       I79224b17e2d1f87175f3118287351e0e;
reg                              I2e3d469ef08219887c92189ad3759da9;
wire                             If000ebe4f2ddbec4afb6c0e41abb2f9c;
reg   [MAX_SUM_WDTH_L-1:0]       I41ee2f859df1db26618ab9c2c0a57be5;
reg                              I74628364cf049f0e6de34bd1f9853985;
wire                             I714abef2427918d8967e5fff40fd48d7;
reg   [MAX_SUM_WDTH_L-1:0]       I15a667ea371ed0fd464f42fb9ef61766;
reg                              Ifec818042c24c8eb96832c782f09ab04;
wire                             I6229267ae259aa8193a90596f8c1d432;
reg   [MAX_SUM_WDTH_L-1:0]       I25c2d3dd7fedd28f0be0e3d8dccddff8;
reg                              I0aa52a892c8969087bf3f158aae7078a;
wire                             Iaa26fea88e8b3f2ce1d402b48c7a9eff;
reg   [MAX_SUM_WDTH_L-1:0]       If22b31d70158d864ca6b0201ffc2b7c3;
reg                              I31b799a3279d7d66b53f4be544498602;
wire                             Idc0f6e44fa41f76f3ddff9628d25c005;
reg   [MAX_SUM_WDTH_L-1:0]       I7950b8505327240095538f60d81834d1;
reg                              Ie8e004bf6e301a4ed9d9dcca91b2dc85;
wire                             I7c14c6e871660c6c830de981c07f6b2d;
reg   [MAX_SUM_WDTH_L-1:0]       Ib75297152c09323c7a6f674c93edc01f;
reg                              I9995a84609ef3fe477c73f136515ffe9;
wire                             Idc5ee83aa6a50531e6de2d9abaa26843;
reg   [MAX_SUM_WDTH_L-1:0]       Ie813deeac800a6b251209a1c8e2adb12;
reg                              I54e519ab156fdf2054472d4684de064a;
wire                             Ie0ff06499371f17cb8c56c9f0c7ee666;
reg   [MAX_SUM_WDTH_L-1:0]       Iada283b3152a5316b6c7077292ac0a29;
reg                              I527950bde49a5c46e818225e41bec4f9;
wire                             I59976ed14d4be22603d2d164399389f9;
reg   [MAX_SUM_WDTH_L-1:0]       Ic14e12a907c5d6b7ad2615905a64886d;
reg                              Ieb876e18857117935ca3aecb6a525b1f;
wire                             I9e94cdbd4a445883fb45fb3ed1b05d7b;
reg   [MAX_SUM_WDTH_L-1:0]       Ife78b0889c9c7129a3000cca66ae4aa2;
reg                              If22f8fa601e72589b3a5779f23ca7454;
wire                             I581b4fe258cb92d51ffc1482da718625;
reg   [MAX_SUM_WDTH_L-1:0]       Id926d49513e089a52b17978a9ab84372;
reg                              If222f8f81e40570854a512fe828f9ea9;
wire                             I19f794db275b2266dd9a91b3b0174329;
reg   [MAX_SUM_WDTH_L-1:0]       I4dfbf2a2c01ce39fea9b756f9b106fc2;
reg                              I6bea78584853c37d7c4993a45668542a;
wire                             I7d4b8ac371172cf90b31890df5693875;
reg   [MAX_SUM_WDTH_L-1:0]       Iad7cce628396ce9ffac3ba9dde7ac494;
reg                              Id7cd91008312189123519e44cfb2e141;
wire                             I1f02219120214ac3e5f5279031facc56;
reg   [MAX_SUM_WDTH_L-1:0]       Ib71f9f92515c200bd16591c656d69ee7;
reg                              Id3c95ac844fe01a85e6251683bb3f9cb;
wire                             I569a8645fa9f5476d122bccc7f40fd75;
reg   [MAX_SUM_WDTH_L-1:0]       I8e39b301e04135b8ab88d54e7c1e22f7;
reg                              I49b96dfb05812ec7b0632bc722d417df;
wire                             Ie620ab2c461442bf7c7ddd962dd65839;
reg   [MAX_SUM_WDTH_L-1:0]       Idadba73fb37b81563818e82af3d89a58;
reg                              I89b8ac7adba1c7fe4f04e408857c92bc;
wire                             I3dc4a3e2c52f2f74aaf1e640543fcecb;
reg   [MAX_SUM_WDTH_L-1:0]       Ic19accaf42ef2b61fb52ab3621622ef2;
reg                              Ic1a67160ca63763ce6b850bed5371d32;
wire                             I749c798e403cefc3782b3a63de02e227;
reg   [MAX_SUM_WDTH_L-1:0]       I94f508ac67f07b73b3ff1d5aa5955eea;
reg                              Iaa1ed0cec8df6dec4fb0ef9c57c98d19;
wire                             I3ce1a50aa7de5d1dae422eed03c450b2;
reg   [MAX_SUM_WDTH_L-1:0]       Ieb8588293562c9c25897044b9e5ed6a4;
reg                              I76465e13c5a9ac236635e663e543487c;
wire                             Id9474b1f0f1ab396654b7048eea873c2;
reg   [MAX_SUM_WDTH_L-1:0]       I671d71d9ca760cc759b96bbacd361f90;
reg                              Iff18998e317563a12db412950315b397;
wire                             Ib7d69d239aac1a9de86e2f2f1337c5f6;
reg   [MAX_SUM_WDTH_L-1:0]       I3f793de7fcfd045af3970e4ec219128b;
reg                              I279642da9295f410b7482eaedfbcde75;
wire                             I40a799391b45437a24bf9c7cbc2ec409;
reg   [MAX_SUM_WDTH_L-1:0]       Id49f950b3679093b10f8b64ae89c5558;
reg                              Iecceba6850d58cd1500bb5129abc8035;
wire                             Id81eae2229fec7726aa687d711d1b998;
reg   [MAX_SUM_WDTH_L-1:0]       Ib70c7567e552969a2757c1f48a2468ef;
reg                              I6ede97dfb1484ba6fe621c7034e22c0b;
wire                             I7bab2b945804593835eb8b63143a3345;
reg   [MAX_SUM_WDTH_L-1:0]       I6dbd0c3ac9f2b3887d87e316b8b40b55;
reg                              I57bf6d033eb5643e96bcdefcfeb76a46;
wire                             I4e7f07fa261e44488cb5b0903d2e8c5d;
reg   [MAX_SUM_WDTH_L-1:0]       I8c309d7fe6aaa8c996e39b8f3dfafef6;
reg                              I5ba33277f07eadbc27835afa96bdc535;
wire                             I5d69471b78cf5aba461a12cfe6d7d11e;
reg   [MAX_SUM_WDTH_L-1:0]       Iefdfd7b1924f8b6049b02576f9948027;
reg                              I256096a960771679c9a7a391448aa711;
wire                             Iba0af171e17c12093f5dbde019fff4da;
reg   [MAX_SUM_WDTH_L-1:0]       I2c14ee79492962576e12ff1698ac0fe1;
reg                              I220f38bf301ec4abcd1e07727fc5bae8;
wire                             I580c7b678e4f2c08a4d521c335392c07;
reg   [MAX_SUM_WDTH_L-1:0]       I56e90395afb09c7d775111d19856da1d;
reg                              Id6cabb7608d470ad7dec1951618efa8c;
wire                             I8016fc36bc9614afef570a084942081e;
reg   [MAX_SUM_WDTH_L-1:0]       I90f0c524f6b98c28d18db952ac40c83e;
reg                              I30ac677d67ab06a6f5759da2717ef6e2;
wire                             I744066a189658aad33b32468934ca485;
reg   [MAX_SUM_WDTH_L-1:0]       Id50649fc4e9de24fdd9f06499a733b87;
reg                              If0881734b6b8bb6e3e22823408203887;
wire                             Ic2a5d82d3e19ff84f46d2d71b3d544eb;
reg   [MAX_SUM_WDTH_L-1:0]       Ifc988e99b4c4c1ba2d5cf3a76695900d;
reg                              I29502a6df7b40a59cb84f6c1a0d30fbe;
wire                             I935a700d902a104974a961beca5ac99a;
reg   [MAX_SUM_WDTH_L-1:0]       I53c579c64f0d911fe3fbc43dc3e981de;
reg                              Ied5d76051c9302e2594e5f1c34dbe8a9;
wire                             I902f91dfb3bada8a106f46923239c93a;
reg   [MAX_SUM_WDTH_L-1:0]       Id729d27d6424495fdb4deb2ffc038f01;
reg                              If6c801f61074108c3342f1c3d0b4a39d;
wire                             I4d4f46a02cffbf72298704e8a0504fe2;
reg   [MAX_SUM_WDTH_L-1:0]       I8816c4edb8c7f5fd6e7a3c81013116ce;
reg                              I3f15fe479ccd6715b63db728ffa8b49f;
wire                             Ie8fd35237928694738b464d52847c2b6;
reg   [MAX_SUM_WDTH_L-1:0]       I88ba486c5bca54f6c120a654b81e0a90;
reg                              Id7e322ddf8565bb59e6377bfc7b3ab36;
wire                             Ib73fc8722db87e7be4b14ce361b79719;
reg   [MAX_SUM_WDTH_L-1:0]       Ie1ba6d92c19ebbc5c994d9da3881f6c9;
reg                              I5a325c188a650a75ab298719c0287618;
wire                             Ifde9664e13fe94aca97da5824ef0c08e;
reg   [MAX_SUM_WDTH_L-1:0]       I023278cb7d70d4608259e10c89e97117;
reg                              I763f7f930d12bef17e0aa5ed0d6abf96;
wire                             I3d25580e525216c23557ffa5ed998bab;
reg   [MAX_SUM_WDTH_L-1:0]       Ib8c744194310bd59e983e392b828e9b4;
reg                              I0e34522d1f95f50998246232512bb60c;
wire                             Ia3d21a8d9a8c24b112965d6eb966de8c;
reg   [MAX_SUM_WDTH_L-1:0]       Iaa2aba39e0454008fbeff8f9aa87a481;
reg                              I45b69f889fd15cce35f6812afe0f4894;
wire                             I7d7923beddaf4b873ae819914599f02f;
reg   [MAX_SUM_WDTH_L-1:0]       I61a43aad15d7a9943f74617f434af306;
reg                              If4db281fdcf771156956dfa30e36b29c;
wire                             Idc6a066b872fa91ce73e9aa21d668e83;
reg   [MAX_SUM_WDTH_L-1:0]       Ibd8114af3027bd3364395e7b94484272;
reg                              Ib312a09daf5e5c38dcd59128256a3ebc;
wire                             I5ea37c7893e55ef146fb831d8c09e87f;
reg   [MAX_SUM_WDTH_L-1:0]       I49167fd9caea095581855b45b1f85d49;
reg                              Iaf3e2d448016a50829b4b0ea6f144b27;
wire                             Ic38315ea78c667a1f77a5fe34ac62412;
reg   [MAX_SUM_WDTH_L-1:0]       Ic502f151ee9ee01786e216d90a29403b;
reg                              Iddbd5820346c3ea47bea79b2ee1ab7e5;
wire                             I2b954aae3ff5e2a0ce92a55107a86a46;
reg   [MAX_SUM_WDTH_L-1:0]       I25f89c7f7f11c7e2811913d6254dbc8c;
reg                              I1b024f329d24692f8d143aeeacfaf555;
wire                             I958138e39e14c8fc1de83d02091b8f6e;
reg   [MAX_SUM_WDTH_L-1:0]       I3f939889c013f740cc63c981d2ff85b2;
reg                              I83f200ddde413f07bd296b8602aacdc7;
wire                             Idfd5a9e4c4cbd4ba9828220a7d021d28;
reg   [MAX_SUM_WDTH_L-1:0]       Ib0d2fc4f353a82d37bec9aa19a80475e;
reg                              Ib4cec30021700f9f02847c2f1e0fc425;
wire                             Ied5041c527b4f04647dc80932b9ce7c4;
reg   [MAX_SUM_WDTH_L-1:0]       I2f19b77e5bb1b22b3cf5b1ace31ee6af;
reg                              I3cddf5a4ce875cb4e0c2fce7e36e5200;
wire                             If6488c8e84e69a99816842a90c9578c2;
reg   [MAX_SUM_WDTH_L-1:0]       I283f82fd4a9700daca6ff1d16f747a09;
reg                              I9c5d93dc3faea27b0f38898609b41545;
wire                             Ic65f12c4a71f8c3af75f426128b333f9;
reg   [MAX_SUM_WDTH_L-1:0]       I8dc5483fb01a06ad8650e5fd4df30f49;
reg                              I426a2f3c939a72ecff6a6314a19d52cb;
wire                             Ica6cd8bf97c702ae2541f682cc418a80;
reg   [MAX_SUM_WDTH_L-1:0]       I7e3f6b4bff19a0644c12fa4ef3667d84;
reg                              I5919e3d3ea27d29a8093c52a6645959e;
wire                             I73054b5829fd26eb2b09dc585f2c62f8;
reg   [MAX_SUM_WDTH_L-1:0]       Idf2371d30bec7ad5dea346a4a48a6e75;
reg                              I68c4ab26cc7c41ea3f9b8afec502bc42;
wire                             I221be7886d94efc9e1ec553acd79dba4;
reg   [MAX_SUM_WDTH_L-1:0]       Ifd5a3069363cfc42e5a436856eeee708;
reg                              Id4ea7f8c016571cc5a0af8327e2f95b9;
wire                             I33557b5dddc36fe3625bf64e016c1c7e;
reg   [MAX_SUM_WDTH_L-1:0]       I1a4e12577ac5e87d40bdcb54fe55818b;
reg                              If6b109772fc17d898d70f75f538a0fdf;
wire                             Ica7d3d482ec7dde7081b68988f76c9b4;
reg   [MAX_SUM_WDTH_L-1:0]       I1f1b6c20910c4f14999da6c9fdb4c349;
reg                              I930235d80caaa415247c7fb380b3a134;
wire                             Ibf9561c2c5242296a3b607627e7e7989;
reg   [MAX_SUM_WDTH_L-1:0]       I1b0a200eea98f075f059d2a26b00f833;
reg                              I324eeb4bf0e552118536fbd641189af1;
wire                             Id0d621bef47b5c5735a4a999611a1c4a;
reg   [MAX_SUM_WDTH_L-1:0]       Ie0dded072843efc1613cfe7136af37da;
reg                              I839160e07222b1f9f293efe22d68c168;
wire                             I33cee0fcc65354655c9e57b3d43c11f2;
reg   [MAX_SUM_WDTH_L-1:0]       Ia6d6a867ebe63a8926d9affa4c15e376;
reg                              I5244962685ce36dd805a7dc774c05d31;
wire                             I8baad814c6bbc783645f574455b0f2d3;
reg   [MAX_SUM_WDTH_L-1:0]       Iddfc447b0c96056ae6e6434799ea00e9;
reg                              Ib92300e3d61e8a2bcaf0b2f40d4cb18f;
wire                             Ib23a7e23bc223c7f3e83661811493229;
reg   [MAX_SUM_WDTH_L-1:0]       I36d03daaaaa37229d462f4bf5e521f73;
reg                              Id76c8bf8796c329353836a52e1dd74c3;
wire                             I55e8b1c375d49a1a1f044a4a60073d60;
reg   [MAX_SUM_WDTH_L-1:0]       I91e49319831eeee5dc75eac77ed8f8a3;
reg                              Ibb163802022194494881194dc6b49c2d;
wire                             I023853b98208afd9bcb1ff63abb91b2e;
reg   [MAX_SUM_WDTH_L-1:0]       I4e9f03752b041491ae2bc40fbd2b8d43;
reg                              Iedb3b8bfd024408f08a2b377956239af;
wire                             Icd656c959fe941e863db11f02d3c514e;
reg   [MAX_SUM_WDTH_L-1:0]       I9a71e50dac7ad707a4b0946ebc1fe6d4;
reg                              I6cfe7ce048413c7c959a0eefe967885b;
wire                             I06cea262d84c35f3e6a1b6690b82cbf8;
reg   [MAX_SUM_WDTH_L-1:0]       I8220d15825d6bac07d773ff0db2f9795;
reg                              I664a362c93dd438aec485063a6f0c7de;
wire                             I1d7bbe81db5320829eb5b29252fc6cf2;
reg   [MAX_SUM_WDTH_L-1:0]       I6b2dc98acc78a1151dd6670ed981d839;
reg                              I9252e19b54173ae2a9d0815dfc46eec2;
wire                             Iafad27be14640dbdcff055b7e34f6467;
reg   [MAX_SUM_WDTH_L-1:0]       Ie371be4323965591a5786063ba028ce1;
reg                              I2ea93b2142eee9f44c8e7bf892bf02ab;
wire                             Idfd58540bb8d1465514c3c843d303825;
reg   [MAX_SUM_WDTH_L-1:0]       Ic4985251ed9f9120d2232ec96949831b;
reg                              I6772834728b2e641c6e3c14cda255ad6;
wire                             I7c98a5f1ea935e4de159795b5dd795ed;
reg   [MAX_SUM_WDTH_L-1:0]       I6015d64c067415fe216d90a5be409e33;
reg                              Id6a64c33b3beb88abcadc06af18e1858;
wire                             I84b1e71a64cd4d96c44444e337dde784;
reg   [MAX_SUM_WDTH_L-1:0]       If6f304fe091216273270713c6b6e8a6d;
reg                              Ib89f2aee80d36f4e473d1a1046e836dd;
wire                             I609aef4d51d5d190deea41f71ef0403c;
reg   [MAX_SUM_WDTH_L-1:0]       I779ee6daefe3c5c96548dc5e0ba83bd3;
reg                              I78aeec1644701502f6f71c64341274ab;
wire                             I68a99adfa01586d1ad7bdeb282f11d87;
reg   [MAX_SUM_WDTH_L-1:0]       Ieef21b505cc215387f8930888062b767;
reg                              I9a09fda6e73783a7c9a4582fec8121b4;
wire                             I1f68aed9a1379bbbd2c531fc0df392fe;
reg   [MAX_SUM_WDTH_L-1:0]       Icbabacaecbbac74901402e5e5874328b;
reg                              I9db6919efaef0952b84eaf8e71f77777;
wire                             Ib1cbee37b3fad49ab5805647ccf95b7b;
reg   [MAX_SUM_WDTH_L-1:0]       I6ec13a161f7f1a0f57e9ba4998474954;
reg                              I5a4646a8adf0ed43a905fd4ee84d85bd;
wire                             Ibbe9c1e2c9f2c0b00e4be25205a824d6;
reg   [MAX_SUM_WDTH_L-1:0]       I71f9823e92c51be2e9a050d01e63902d;
reg                              I1e3444ee88dc52881397d266f469b45c;
wire                             I6c7e0e56cd76e03261638e924f90377e;
reg   [MAX_SUM_WDTH_L-1:0]       Ia0037030d79400734732f061fd81edf6;
reg                              I3c42e969e5e4b99f1f2eaa01419d4ed9;
wire                             I676d7f8a89fbbef4b067d07264ae427c;
reg   [MAX_SUM_WDTH_L-1:0]       Id796584e3e7af67536a27f7299b71916;
reg                              I9210d06734058f76e7a5a470dbe6e74b;
wire                             Ifcaf093fbbec17632ca0050583df41c4;
reg   [MAX_SUM_WDTH_L-1:0]       Iec938bc1bbad930fade05d74c10989a3;
reg                              I2b35c8fa7c947b3e7691cdcab0c5a7a7;
wire                             Ia358ae5a96e63f3bb5c6bb34f263c387;
reg   [MAX_SUM_WDTH_L-1:0]       I2a7a7c5eabd1623c1c3d4bd93bf18617;
reg                              Id58d1af007bb5858499af71a43e6574f;
wire                             Ib1e4443484bfc289563a8b7d9b1c86b6;
reg   [MAX_SUM_WDTH_L-1:0]       I71cfc7fd85636c5554b9fe9f9ba8e3aa;
reg                              I12e92aa9c9ca2135f7ba879d82ad615b;
wire                             Ib3baee13e51f9fb8c39d04211497e274;
reg   [MAX_SUM_WDTH_L-1:0]       I4c8ae97548bc3dbf3e3621f80c3e0835;
reg                              If32ea54eb47d27e35a81aa4b9e1f7713;
wire                             Ic24de5d8c9148fab7b9dcac9d8996740;
reg   [MAX_SUM_WDTH_L-1:0]       Iaa93c760705c984a0eea90d41a6c049b;
reg                              Ib1ddab09d1a726176414e4a877b66e3f;
wire                             I46489795c1a8e178f1b2d40711655c44;
reg   [MAX_SUM_WDTH_L-1:0]       I2acc73851f8a803e69c0f1865e00f46e;
reg                              Id3838f634ce2d90a19622185391ba868;
wire                             If39c47fd6b6913ec7946018145d31945;
reg   [MAX_SUM_WDTH_L-1:0]       I928333e9cc75d49fa6f7094e49631123;
reg                              Ia3f429c43f23f4f057abed98cfa94748;
wire                             Ie336a92376f51b145c60f935b8fd0f8c;
reg   [MAX_SUM_WDTH_L-1:0]       Idf02dd4b7e8a6958913e6180fec1feee;
reg                              I62b423a6061215d16871bfdf9a9cdbd2;
wire                             Ia6f981e46e3d7ead096d73154e97dca9;
reg   [MAX_SUM_WDTH_L-1:0]       Ib30cc7931858974728d92eb68890449f;
reg                              I17f82f6daa8a92f1da5a1952a558ad7e;
wire                             If7593819b136ad3db74d793e5a0f18c3;
reg   [MAX_SUM_WDTH_L-1:0]       Ia504dbcee6e5894fed83371bf70b2d44;
reg                              Ie0e9f7c1d69d8930f8452d3618512877;
wire                             I0b480fa6fe571ea7d25d13f8f1ba26da;
reg   [MAX_SUM_WDTH_L-1:0]       I32b4e50b8acefe1c108d777da565f4ed;
reg                              Id9de214d84792861772ef396b5b9208f;
wire                             I66ab48b076a0e2006d1f4741e15f3c36;
reg   [MAX_SUM_WDTH_L-1:0]       If9fd1d8c0c13042a6f2d258478b63925;
reg                              I027f018e60dda98666458cb69a6e4be2;
wire                             I9e397fd8cfd4ee1b9cd3cccbd4c03005;
reg   [MAX_SUM_WDTH_L-1:0]       Iccb437017198e4421ab51d74aed779f0;
reg                              I996821515569c215f3f688d91dee8abe;
wire                             I177684367c872f5a3df89c0d2bb95434;
reg   [MAX_SUM_WDTH_L-1:0]       Id10bf2bf52a8f1be9eeafcefd6dd5dcb;
reg                              I6f617bfa2700fb385d425f6b4581f594;
wire                             Icdb37cf629ec16db879e288eba5ef9a9;
reg   [MAX_SUM_WDTH_L-1:0]       Ie590c921147b7252d2605f7712dfe437;
reg                              Id5f8b6b344dc8e629f13e5d157f510cb;
wire                             I225d035b7f8d13e9895ca60f3da8bf90;
reg   [MAX_SUM_WDTH_L-1:0]       I178ed883c28bbf3e1ab05cb95f62b343;
reg                              I579a5dc98f16e0c5d52fc7958586a8d5;
wire                             Ia3572b856ec1a14e316444c2f15ac9a5;
reg   [MAX_SUM_WDTH_L-1:0]       I01971a175615a422d264805252f91f3b;
reg                              I0f2769698735ab28df30370c3c8b56cc;
wire                             I2c927c7ee3628a78f48c6099d2036959;
reg   [MAX_SUM_WDTH_L-1:0]       Ie770c4567f35b40c46ccbda059e6d3a8;
reg                              I9fbc79fd7be52757770dce6e04749b4f;
wire                             I578551b6331fffa97a6d05652e406e3f;
reg   [MAX_SUM_WDTH_L-1:0]       I25975702f0b9c0baf586fe471676dfea;
reg                              Idfe33235c2f93ac311da89ba63e0f1c5;
wire                             I6f301798efb2c67ea363df40f2fe340f;
reg   [MAX_SUM_WDTH_L-1:0]       Id2ef737d910326394b68eaa0833bfccb;
reg                              Ic46d706f6be34cb4133a4128567837d3;
wire                             I744d142b9316b9f8937563c1023882e6;
reg   [MAX_SUM_WDTH_L-1:0]       I577cd1f9ad512ec10f5008165f2e4a74;
reg                              Ibb3c635f2e62a63c9bdb150b3cda7155;
wire                             Id7fa5f9fb6059439297f246cb228cc02;
reg   [MAX_SUM_WDTH_L-1:0]       I1de8f87eb39276e073f5804b1df3b67a;
reg                              I7bdfb2d2b7dd18fc7c0d43b708fb1e35;
wire                             I18e9dd5583f3ac91451a4e75f0d5d474;
reg   [MAX_SUM_WDTH_L-1:0]       I7f8e7928e6caeac14f787d7e0b6a47df;
reg                              I42a1cd616514a1c7384d07095e6b2d70;
wire                             I64afac5bd1ea7a2ab696e630cc3ad162;
reg   [MAX_SUM_WDTH_L-1:0]       Ia7048aa3f949b0b2e54ab900efe01131;
reg                              I19a91106f189ef43ee50edab49d297c1;
wire                             I0b3bfd6ce482cfb20d461862a0bf8f61;
reg   [MAX_SUM_WDTH_L-1:0]       I1fcbb73d165eab038c745fac370fd68f;
reg                              I90088e4928092e62e193039faf154240;
wire                             I16119df9372ce61c0c8600ddba36e607;
reg   [MAX_SUM_WDTH_L-1:0]       Ia822cd52015d599bc45ae7338b4e88e1;
reg                              Ic0fed8f997e03bcca119270589f8bf0a;
wire                             I0957a6c9a87bc89dd9748491807837af;
reg   [MAX_SUM_WDTH_L-1:0]       I56b85e2d5a7259eb50fa983b92d8b160;
reg                              I3ba811abe28766d976a2afd02c22fc76;
wire                             I12f8c91d67e31e11033d5b3b266c659b;
reg   [MAX_SUM_WDTH_L-1:0]       I1d23632f8e8f66a30b4ef6c76aae3ece;
reg                              I66463d17d0fcb691e727568e4d55ae43;
wire                             I690b96154d7717bf62eeb740b10ce6d5;
reg   [MAX_SUM_WDTH_L-1:0]       Ib578de11f0407cfeb0dac68bd5fbf7a0;
reg                              Icf73bfd92fe6265b8e7d9b2439573a96;
wire                             I25b3993479d7cc172ba6a480628b9188;
reg   [MAX_SUM_WDTH_L-1:0]       I08879fb80c58de5fb2bf547ce013c67f;
reg                              I7c3f7076072ee81960c8b0187648eb41;
wire                             I7f3a220cdbf5bf1737690e1719f888e5;
reg   [MAX_SUM_WDTH_L-1:0]       I8f7c4c602b7de5d9a401d3933a7e50a8;
reg                              I68ccb34c409f89f1a2872d64f85e3245;
wire                             I8d068dee7478a9f899c8145ef6d824a5;
reg   [MAX_SUM_WDTH_L-1:0]       I2ab4cc1ef6b743cda8765a22e28fd7a7;
reg                              I069661eba4d8f68a4e5c78e99e9355e8;
wire                             I2286af8d6007a7da5c745d75f407b5d9;
reg   [MAX_SUM_WDTH_L-1:0]       Idc58a89f7d8ee884b198b6e4752ec58f;
reg                              I6cc756f9cb1020c8045872d628b771f8;
wire                             I214f77e05ac2ce4b94d4c5e53675717d;
reg   [MAX_SUM_WDTH_L-1:0]       If9c0f4c64c7648e509077df16c14b7a1;
reg                              I95494fb67de54f6055f54c7568106488;
wire                             I8fc900d4110bc862ad7287255dddf2f0;
reg   [MAX_SUM_WDTH_L-1:0]       I8cc434418203702ad5a21eb4f0340dc5;
reg                              Ibbfab9efcd61f23b09e371554c0778b0;
wire                             If609e068414eed49fbe97f86e2546768;
reg   [MAX_SUM_WDTH_L-1:0]       Iee9d96f800fc848f3c4b6b6901a72623;
reg                              Ibb2a246712268d6d8a0ad0354b8e611f;
wire                             I69177c754e87bc42401bccf54b770358;
reg   [MAX_SUM_WDTH_L-1:0]       I989036e56c9c7386279e83ae83ad4f7d;
reg                              Ie9f5d2f06f60d7f436118f2c92695107;
wire                             I3b121702ca62507c2afda1ed93183499;
reg   [MAX_SUM_WDTH_L-1:0]       Icf23ca0439c76198fe647a0b785d9503;
reg                              I0ee25f335a84b7a190ccd690fccc1fce;
wire                             Id979aeb39d36400b85386a8e96ca5a35;
reg   [MAX_SUM_WDTH_L-1:0]       I406bddf2c4a4b6e6aedb86d72f14994f;
reg                              Ica83129589b16c7392387bcddd9e81e9;
wire                             I61ca2dba668792ee6a83850e2f118eb0;
reg   [MAX_SUM_WDTH_L-1:0]       I5331e97930599788b1df06992c5e4a5c;
reg                              I91fc1c1758eb8c136744c1ef47785b49;
wire                             I7e7f1d73e81031a38992b4f9a3f90717;
reg   [MAX_SUM_WDTH_L-1:0]       I98577e71126ac9bdbe4359101d4d48d7;
reg                              I2bede76feb8d499cef693a3cc0bb95f4;
wire                             I029dbf330bab56469b88cbd602e8e16b;
reg   [MAX_SUM_WDTH_L-1:0]       I696f551b6f96d0f7d27eb685bd374229;
reg                              Ia0d9b7bd503ddeeefe9d0646c1f4e6d8;
wire                             I47ddb6cfe64c5addb3900e193094ac8f;
reg   [MAX_SUM_WDTH_L-1:0]       I1aa256ab19406597846ff353b65224cb;
reg                              I2af1f93bd1d85a66028ef0add7a69962;
wire                             Ibdf7e609b7e42c57450d9d9fdd610881;
reg   [MAX_SUM_WDTH_L-1:0]       I00f1b24291a0e8496e13fe076e377cb8;
reg                              Icc568348313201d6814f92694d7db06f;
wire                             Ia096e8920afb814330e53778c955f8b0;
reg   [MAX_SUM_WDTH_L-1:0]       Ie6f40dc356120aeb6cfa7a3fb5fae8cc;
reg                              Iba815b719f813a245efb2627660634ff;
wire                             I365fd3d16d984516e33a7b68338d0384;
reg   [MAX_SUM_WDTH_L-1:0]       I67e23e6286edc4e01a7ebdace62ce56d;
reg                              Id67d39730eb990c4b125cfa772e27e3a;
wire                             I5e86c33e58b50627d7e69a4200525e05;
reg   [MAX_SUM_WDTH_L-1:0]       Id2c7c6d20146edcca65120c025e25a0a;
reg                              Ib09008d80ae9d6708371c0c40f157656;
wire                             I52ef2681091d643e4ed026581feeb3f2;
reg   [MAX_SUM_WDTH_L-1:0]       Ida1e2d8b0e45e14c4c669c8b9d6947f5;
reg                              Id61b17db82e540f939ed8a4c3b596278;
wire                             I0e30717ed1e983e1c5af25037d5cfca3;
reg   [MAX_SUM_WDTH_L-1:0]       I1fd443d00410d0577eef9f1f26e64700;
reg                              I24868694c2523bb657da19c2e84ec8ef;
wire                             I640e720e6aaa2f8e14b5dacd51cc6e66;
reg   [MAX_SUM_WDTH_L-1:0]       I9ea760f08ba7b84fcaad929a3669450d;
reg                              I9dcf88e53c655bce8190c5e85f5ca777;
wire                             I81f4ac1f01d8170f427ee5ef89e8bd78;
reg   [MAX_SUM_WDTH_L-1:0]       Ia522420603dbde92a49da297554ede5e;
reg                              Ib881ec4b6a6de42dfcb2be830ca39ac8;
wire                             I8319f97640191977a9b89e7639aee739;
reg   [MAX_SUM_WDTH_L-1:0]       I9be575cacaafcc13a0306545be56a04d;
reg                              Ifd2ece02d5ffb0a50d8b151a8fa8e703;
wire                             I21add24f8eed563787b8567fe43947f8;
reg   [MAX_SUM_WDTH_L-1:0]       Ieb9a03ad2c7c7df356477e8b4224ebd9;
reg                              I7da3a787760c42ef510ece8234c020a8;
wire                             I1a772b29d533c44422332cf291d27253;
reg   [MAX_SUM_WDTH_L-1:0]       If7f263cb2fb7fd35682d44c42639bab6;
reg                              I2204fa0d852e56e843393b3959f3df72;
wire                             I8ec002e0ccc2cee9a210b987bf1cccc7;
reg   [MAX_SUM_WDTH_L-1:0]       I5046227e18f800785f8ddfb4a89b1bea;
reg                              Iaee3ca649d20dd29363781e8dcae17c0;
wire                             Ia13212b613a21e983b097fe0adbe59ec;
reg   [MAX_SUM_WDTH_L-1:0]       I73feb8438775bf3faffed6895b6a4638;
reg                              Id8bb7c6409e383793af592892caf23e4;
wire                             Ieeddfaf876af8120f779286b4f60f767;
reg   [MAX_SUM_WDTH_L-1:0]       I6a423d4e11a97d84120a475db8fabca1;
reg                              I96c6b861bfaad7c411db93f1318d6b87;
wire                             If1912201b852f91e8aa0c73439ca7022;
reg   [MAX_SUM_WDTH_L-1:0]       I2098616787bd728bc4af6be5ee094bae;
reg                              I76eb400ed4d1502f7f1864d9556948ad;
wire                             I0995a527d1b13090cf68b771d591c041;
reg   [MAX_SUM_WDTH_L-1:0]       Id9ef21a12edf48e574256ea34fcde992;
reg                              I02155a5c26345ff00d18cec6e2f01592;
wire                             I04bb94f5e9927cb7efa70e68658862d3;
reg   [MAX_SUM_WDTH_L-1:0]       I31ab57596896201ff52990b0641b9511;
reg                              I91e6dcd9fa2efd055125878ab38de3fd;
wire                             I7594f22f889c391838f987765ad478e7;
reg   [MAX_SUM_WDTH_L-1:0]       Ib3dd33a163b0c8153edb4fcc90a453f2;
reg                              If561e078b234a0be8c0b8ade8f5ec0f1;
wire                             I93a25759f720769b941088884bb6db59;
reg   [MAX_SUM_WDTH_L-1:0]       I28496a34b2ee033767fd64f631426b23;
reg                              I0ef01533d6494ce8f092d54c5fb0865e;
wire                             Id518694e3b3a268e7168c17250bfab52;
reg   [MAX_SUM_WDTH_L-1:0]       I0a4ef7fac369df46d1a4b094d7687645;
reg                              I782b73148fd7ed7f9d734baf42b8b5d0;
wire                             Ieaf2b41941b840b3ade630e721e6367a;
reg   [MAX_SUM_WDTH_L-1:0]       Ie7944f3e2adfac325808f8711c0eedcd;
reg                              I2099d6f614a5f7432f6331b1bf56c31c;
wire                             I01a2be56c727d7ca0c5059e8d34919cb;
reg   [MAX_SUM_WDTH_L-1:0]       I58cecb5376f675339028440f0671b0b7;
reg                              Ia8c9228b5d23c91ac06450ab1296dc65;
wire                             I605682c90ff448b91a2e1a82a3cb0c08;
reg   [MAX_SUM_WDTH_L-1:0]       I62f85c1602819e586d9656ba42d263c3;
reg                              I4b76ea8b5d4ed8ccd8ec532889dd6d4b;
wire                             I0a075b833950927c58d8f55264947f00;
reg   [MAX_SUM_WDTH_L-1:0]       I79585885950084095d2ce4a31aa73e4c;
reg                              Ifff6d20dcf891c78ad12a304ca757c95;
wire                             I3b699342f0100a2d56c7013da055fdd6;
reg   [MAX_SUM_WDTH_L-1:0]       Ic3af09106eada35f1d786ed60e314ea5;
reg                              I0dbefebca7ff055a6e9dce2a2c37bd69;
wire                             Ic223e47525ca27261b7db8c1afddadc9;
reg   [MAX_SUM_WDTH_L-1:0]       I81e374d671edb31d060875cdfdcd61c7;
reg                              I8aadd755861e90ac12047f259091ad85;
wire                             Ibb5c74ed3a37c5e244e537e8b8d403fb;
reg   [MAX_SUM_WDTH_L-1:0]       I1e22ea5ecaf87499b7106246a824a547;
reg                              Ia7d21a17d62e7bfb00b83b244201e941;
wire                             I5915ba867f798193c35a4af58e8cabf6;
reg   [MAX_SUM_WDTH_L-1:0]       I0e46eb0f32c91384b07c7b1ba84caf98;
reg                              I6c63fab8059cc3f0c02b0dff5a8cacf9;
wire                             I73ce6acb5ca8a57906440578f4ae15aa;
reg   [MAX_SUM_WDTH_L-1:0]       I562b5f77aedd91f0cb3df00387c7956a;
reg                              I8744fea2c7de33b5308dc9a2828647d4;
wire                             I9cea4e30593a1275f4450adb25b5c5cb;
reg   [MAX_SUM_WDTH_L-1:0]       Id819e47f502c18dca8d1e804d346c1ea;
reg                              I04c99b4d0c54b23a72b698753510a4f3;
wire                             I3dacee8649adfc1a8b2092f5af3cada6;
reg   [MAX_SUM_WDTH_L-1:0]       Ie0586f4b015fd32777d24c2d9856b27f;
reg                              I5de86a27849e73b21e4c40e9e8515033;
wire                             I00537a49036c970d6df97b3917de104e;
reg   [MAX_SUM_WDTH_L-1:0]       Ic28248b41552d2537d0478c23e33e0f3;
reg                              I185257f76b2886cd845e50a01ef5b05b;
wire                             If6ce1f97c23f1d1bf23c283ce37682ce;
reg   [MAX_SUM_WDTH_L-1:0]       I3463cbe0d16b14aa670fda6a0d34e255;
reg                              I1a2c7b5505f4124f945a28565eed6013;
wire                             Ieae92b67815d507df906e1be71d6346b;
reg   [MAX_SUM_WDTH_L-1:0]       I0aac7a09d9253385d34e87bfbb216a79;
reg                              I771d417f6226b04ef016d0943bbc4584;
wire                             I1af89e1ec1210d4d3dafc0927b62afe5;
reg   [MAX_SUM_WDTH_L-1:0]       I305967a657db8531d1ae309fa3e3b98f;
reg                              Icb0a73f2dd46e2195d5efd34fba3a985;
wire                             Ic264e7826b90e379048b094875eeb921;
reg   [MAX_SUM_WDTH_L-1:0]       I0524108ee49eec5fa7861bed35e4ea3c;
reg                              Ia992f7eacefc028526ab4f105e244e02;
wire                             Iea6d4bb1137e579b1605a16c578cbd7d;
reg   [MAX_SUM_WDTH_L-1:0]       Iced1e0b874918a1c66e28752e340a51b;
reg                              I85454620b6568bb7fde468a2e9a5fb42;
wire                             I706d85c9d83bcfc5a2204a67e5c1f84e;
reg   [MAX_SUM_WDTH_L-1:0]       I670e910f74fafccaa9f1a8279fd6ebb6;
reg                              I87557ef641a7b209d4d210498bb15271;
wire                             I6e832b004d0dddf4c3edb682669acf7a;
reg   [MAX_SUM_WDTH_L-1:0]       I02fe6b32b2405fb94afd5d7abbaf0195;
reg                              I28d1125b647b953f2a19ecd6edd8e450;
wire                             Id0f69c70b38b7483a19e32d5982bb4b5;
reg   [MAX_SUM_WDTH_L-1:0]       I5f5304e4b132f816c87248d3ca954164;
reg                              I4a8aa3010248f0bdd3e31822bf2fe0a1;
wire                             I9cb245dceba82553db23cb15854f59f1;
reg   [MAX_SUM_WDTH_L-1:0]       I0ecebe47e1a9ede33c3995945a6ee760;
reg                              Ie1966fd5b564dd6eccfc458e9c6aca2a;
wire                             I978d0157f7403d2f35fa648271f4fbd9;
reg   [MAX_SUM_WDTH_L-1:0]       If425109071b5310e097d2174625b6383;
reg                              I8ad51753f106d0a30cc79bd08e799348;
wire                             I70e5f31e8c4f1aa9a9aa21c28ba20d08;
reg   [MAX_SUM_WDTH_L-1:0]       Ic0f324c7ba05a7cfae9d70b62e30f94b;
reg                              I1c3bf915a6b62d22d04b8c8d92a72a73;
wire                             I3cf2040a93a0184f619ce941c4f910d0;
reg   [MAX_SUM_WDTH_L-1:0]       I35631cbe926290974c90ddeb9b07f231;
reg                              Ie557629e9d52e5fa7435b4fb19e5276f;
wire                             I3278841178f87a4d0ccdf8316c3fb689;
reg   [MAX_SUM_WDTH_L-1:0]       Iceae425f37f3b1194a2ef5cd46d1b6eb;
reg                              I38fc977bb1d52cbc5e02a6733f6a8190;
wire                             I73d0e5f3635c5a2c3f1824c578c07658;
reg   [MAX_SUM_WDTH_L-1:0]       I4faa2187d970078870078c3eff180b4a;
reg                              If84914aaabb020baad2b222f27c9ad38;
wire                             Id1b7ef639fcb74c8fa47fd7ef0cbe96c;
reg   [MAX_SUM_WDTH_L-1:0]       Iec2860f518edf688a9b1b2736ae00835;
reg                              I54c457a658721fa7de175432b340532e;
wire                             I1c83edeea3cd4c32bae64594a2f8b256;
reg   [MAX_SUM_WDTH_L-1:0]       I20e7b48527e4456874d59e50c723c6a5;
reg                              I9036f6cf74a2aecd827c7239da13db70;
wire                             I0b930276a1887380da03c22aa8fb9adb;
reg   [MAX_SUM_WDTH_L-1:0]       Idd60af0dbb02680e11c1b1734f23b895;
reg                              I8825e2665dcee58925a5106a9cbce9ca;
wire                             I63ec886123f0ff76bfa46c2d6b2c5760;
reg   [MAX_SUM_WDTH_L-1:0]       I79cfbb5d5e920bc8cece60565ee0c5c2;
reg                              Ic3311c2f88a7ae151999b2de86d82dfc;
wire                             I32bf44d4f4df42cb664e75ccef06fb34;
reg   [MAX_SUM_WDTH_L-1:0]       Id765a3f659dcdf01cfe23cafdf066f92;
reg                              I3ef7eddb92284b28f97feea52f489aff;
wire                             Iadc0319541fc978cd0efbdf5b3af7078;
reg   [MAX_SUM_WDTH_L-1:0]       If370aaa56b4ba3eee873c99a86577c3d;
reg                              I68728d0cbb3a84370006277186a0829d;
wire                             I9f4036502b40315cfa7d8bb9b83b5806;
reg   [MAX_SUM_WDTH_L-1:0]       I4508376202467dc1bebc69757bd5f95a;
reg                              If5bdbdfa73406a6a9d426920f51fbc73;
wire                             I91dd649eab4a8eb0f8d97553560d3b7e;
reg   [MAX_SUM_WDTH_L-1:0]       Ibf115f80ad72df8599073c05ac58e028;
reg                              Ibd3179c01665a17f9c232196648de8d5;
wire                             Iee09e9c54961c380ff7e1758c84d663e;
reg   [MAX_SUM_WDTH_L-1:0]       I27960a9d3923d053d466955c660a91ca;
reg                              I42c2c03a158ed79ea91ea6b9f9a6f243;
wire                             Iaec27722c40c7cb0c0baaee4d30adc72;
reg   [MAX_SUM_WDTH_L-1:0]       I7c52711e3b71823dd47861341d22adc3;
reg                              Iec064c18b262b95bd6412b1e50e4b5ef;
wire                             I5fe79d8695d426ba54609af4b38bf2dd;
reg   [MAX_SUM_WDTH_L-1:0]       I547ea6a130740e4b0bb85f6c9d3a6549;
reg                              I0470f0fd133851c1241c654abc19992a;
wire                             I8a2b1e09c6f852b0aa4e599e7ef42187;
reg   [MAX_SUM_WDTH_L-1:0]       I0ec19c18ef7da4793427a00a652a9a35;
reg                              I550661edfa7a7b440d43c0840aeed8fe;
wire                             Ie1f415cbb2d3e1d46f2e0e4201fe7ba0;
reg   [MAX_SUM_WDTH_L-1:0]       I640d147f241267ccc89f9ab132d724f8;
reg                              I2f01145e1b41f2f7103c5247bb548a6b;
wire                             I46a75678565a43e0da6b6dc55686c4c8;
reg   [MAX_SUM_WDTH_L-1:0]       I3507152877484394769c12879ce0aed0;
reg                              I34d143e9a6f936b83863a5ebdf8afc43;
wire                             I200bec7d713bc7f05dc3931f20523763;
reg   [MAX_SUM_WDTH_L-1:0]       I382f86490f568ead2dcf51e8bc6989f8;
reg                              Id2f831bc219ca3f43c5c4d69f6724e64;
wire                             I978b7018cd38c7c4f0b6199cc46d258c;
reg   [MAX_SUM_WDTH_L-1:0]       I953178c54a672474dda2f48c70ec21a7;
reg                              Ib708fd61ab7016190a2a7156439201cf;
wire                             I9d298dcd244445c8a047a1ac056fb6a6;
reg   [MAX_SUM_WDTH_L-1:0]       I13b43982093e885ae7bb04a2b61e4eaa;
reg                              I6a2e574a2d27e40faff379b6c26ae51b;
wire                             Ib5de0226d215418202f2cff36b573daa;
reg   [MAX_SUM_WDTH_L-1:0]       I3d7491ac28a4adafbc138d17f08c9111;
reg                              I4be2286baca2745e981a0d153c0f5c42;
wire                             I58e42ededb36d8aaf022e7b42a8fb36c;
reg   [MAX_SUM_WDTH_L-1:0]       I3e0ca15752add87cc01981e7d89d53f2;
reg                              Ib9643265dc8c283d7b0c7afdb19101fd;
wire                             I8017904689642a7e3d82c34839403614;
reg   [MAX_SUM_WDTH_L-1:0]       Id1b152deea3ee894ed5a4c6ff10a6fda;
reg                              I78d7637bbd13c620434d3619e615114c;
wire                             I773d6a848aa20abe6d1ebf8f7d6dad85;
reg   [MAX_SUM_WDTH_L-1:0]       I7df9cc0e3ad69985fe9a3c8f2dec1de3;
reg                              I358ee555d9955cdee436375ff898f4d6;
wire                             I8bafb2d0a6bf186c179ee07ed51a2e33;
reg   [MAX_SUM_WDTH_L-1:0]       I52910c0c2d26095c965d32b85e850d92;
reg                              Ic3961c918c81b14d964e96892b95f00b;
wire                             I63d8a99e826b0d6a5051fb454f15f44a;
reg   [MAX_SUM_WDTH_L-1:0]       I93fd4b4f7d01ec59834f3054fc2eddfd;
reg                              I580e98d4bec3eeeb1642baa425a96099;
wire                             I0b831c8e1d7187024eb93f980cb04f61;
reg   [MAX_SUM_WDTH_L-1:0]       I481b6feb1f1ced501a157b06a4782e05;
reg                              I4cec0a54301908b3f58166a9b0ef1eb5;
wire                             I17867f12563819dd7b89f9079fb0a385;
reg   [MAX_SUM_WDTH_L-1:0]       Ie99b8f3190ee307e743255156b7f7f90;
reg                              Ib7f7c88d83d207bac3daba4658342879;
wire                             I2a2b4eaef143deb9e61110334dc5c2ea;
reg   [MAX_SUM_WDTH_L-1:0]       Iac858597facbc0025a4760eac49531fe;
reg                              I371401ca0c589a1b8fa816beed36ab0c;
wire                             Ieb02d465c1ac76962dd663067ebcd445;
reg   [MAX_SUM_WDTH_L-1:0]       I18c2833554a5b358578e7b6901c91c0c;
reg                              I81f561f223b916600ebc572c05dedde5;
wire                             I6ad4bc4bc7c0f005307199814893faee;
reg   [MAX_SUM_WDTH_L-1:0]       I0cc6945a47b3ffadd1e52e3f71c9728d;
reg                              I7ee36d73f8c69e5e017f4616094d992f;
wire                             If9a814db74759469b79411ed7038c860;
reg   [MAX_SUM_WDTH_L-1:0]       If2807866c5d481cd31c69b67ec537a4f;
reg                              I706d7d2238c5882491d479df0cc40c3e;
wire                             I3d0f05a6136e0c14536830bc53a5333d;
reg   [MAX_SUM_WDTH_L-1:0]       Ib24d495a86e15d9c8b2c8d360445e511;
reg                              Ie28bec241cb36d75c1f2ad846dc5c7d6;
wire                             I1f168715063587b7dfb01e0fefbca615;
reg   [MAX_SUM_WDTH_L-1:0]       Iad2cdac80bc26a0c50335c6467921c94;
reg                              I9fe8aa4f9f74c1f004e5bb536e902ea2;
wire                             Ida3cc6922fe4edded7f2e59b909d6d72;
reg   [MAX_SUM_WDTH_L-1:0]       I18c93f107d0520171864b789ae9707b9;
reg                              I444003b27464f275311d07ae7d4fe016;
wire                             Ic2b81c5409d555402164dd12ae7decc4;
reg   [MAX_SUM_WDTH_L-1:0]       Ifd40aae90a89d2420e43fe4ee533a1a2;
reg                              Ibbe636e1e98bbd4cd97dca56d769d269;
wire                             I8edabaa27753c6f70325108c9c1b12b6;
reg   [MAX_SUM_WDTH_L-1:0]       If46a176f32240b03ae959e9ad889fc2c;
reg                              Ib195ccbfb4411bd3aaece336a5aed65b;
wire                             Ie58289ff961fc431fbf10f78fda337ab;
reg   [MAX_SUM_WDTH_L-1:0]       I5e7b386298be05835cd24554966cdedc;
reg                              Ieafb75c62922cdb3acd95a9614a86efc;
wire                             I3ee219716889ea93423603105de22c6c;
reg   [MAX_SUM_WDTH_L-1:0]       I5258d2bd4ae07dcfe7e022b046800856;
reg                              I5d7018ab259e054ecb48a238f3c03208;
wire                             I957518cfe822b5afcc1f7153e07e26c4;
reg   [MAX_SUM_WDTH_L-1:0]       I14da6601ba08fd3e9a2bcdd20bb43536;
reg                              Iedabb09ffcf910c4dbed2f142dc96df0;
wire                             Id8fb66bc4afa4f7f7f4ca0d7ce3f5543;
reg   [MAX_SUM_WDTH_L-1:0]       I76bbfed1a115c2f503531682cd171185;
reg                              I07b84cae4f002659d68f5c1746416e70;
wire                             I3beb0bdc4242c12a068f7aec11bf022a;
reg   [MAX_SUM_WDTH_L-1:0]       I64f37f25618c6bf5b35e863e3be05a3e;
reg                              Iba31516a82e9d2a5ad1a1c89dfb6af70;
wire                             I629a5a30684270d00605b4fc02eab693;
reg   [MAX_SUM_WDTH_L-1:0]       Iba3b847497a7572624a3a1f172b47d3e;
reg                              If5c42feaf3d586e1f2285b0f3e3a2d39;
wire                             I32aa431be1c47b8c52c3b3f6d371f439;
reg   [MAX_SUM_WDTH_L-1:0]       Ic9885fd472d244d4810bc9ff0971dc65;
reg                              I3f15f6722f339c32bf1dfa41b5b24648;
wire                             I88d8124a68d50e1730a87914ed6b2a55;
reg   [MAX_SUM_WDTH_L-1:0]       I5753bb74c9d925b91c0173bcc320af36;
reg                              I74d5d4a25b6ceba088652dbad9c35bae;
wire                             I474bd0d0a044aae82cfb1afbd3d40f74;
reg   [MAX_SUM_WDTH_L-1:0]       I66cf73ce0a93f90287df52adb628716d;
reg                              I1e3e7019425109b26d4ebc7522074e33;
wire                             I2bcfe7aeef8f2b772605c9ad10a289ea;
reg   [MAX_SUM_WDTH_L-1:0]       I84a477263ea86f2014d28e9ec928fa1b;
reg                              I4f0d4baa740b2f9bea59f4653cc9e8fc;
wire                             Id4a7c3a22060cfcaff64e2a3980dea91;
reg   [MAX_SUM_WDTH_L-1:0]       Idda9e2f9a5e24406700b04e6035dafc7;
reg                              I2df393a2d764f120433f310797abb2c3;
wire                             I6085d7398ccd685c1a60a21e4a15a606;
reg   [MAX_SUM_WDTH_L-1:0]       I694ec5f3a1e7cfc02c1af8369064967c;
reg                              Ib9a2e4c37430ad33531f318a313d4646;
wire                             I203cd1948326fb3fa3dc14423bf3f992;
reg   [MAX_SUM_WDTH_L-1:0]       Id0c6285ee3789c104e483a5626b5827d;
reg                              Ide344589b18aa0332a7114424956b65b;
wire                             I67412169057453e2fb39c3b0760039c0;
reg   [MAX_SUM_WDTH_L-1:0]       If9bc7b1498733ed921b51cb613c2cf53;
reg                              I789b8e58762f722bc0e86e17c2655965;
wire                             I520d93aaf6b72a2ec7c23ae4e253aa07;
reg   [MAX_SUM_WDTH_L-1:0]       Ieeda4b6b301d662ab9be9f6b979bb1f1;
reg                              I243898aa7700f57974ea2834df469f48;
wire                             I34a77904a4a75d2907acd173bf27800c;
reg   [MAX_SUM_WDTH_L-1:0]       Icad98c93196218a7dbd25af042b4a32d;
reg                              Ic65d6b89fc082438b9956504f30a5483;
wire                             I7a4ea8ffce8d52bb241553a681408dec;
reg   [MAX_SUM_WDTH_L-1:0]       I408e198b0eeade8b94c27ab7e04a8776;
reg                              Ibdcf7926e0b7412e4a56d2ae15a4e892;
wire                             I8e89fb1ed1d604bbf0177e0c61da6e94;
reg   [MAX_SUM_WDTH_L-1:0]       I24b90526a93dc177a5d23b61d20f8797;
reg                              Ie552917ecc454608adca6dbc4d9153ad;
wire                             I5d2148b5809cd169c41663caa441c464;
reg   [MAX_SUM_WDTH_L-1:0]       I4da324410e88d8c9738949c287e7bff9;
reg                              If3b234f8485412e76e5cc497b7c3a6f7;
wire                             I5bb0ab59e3468a9a95b65bfe58acd6a5;
reg   [MAX_SUM_WDTH_L-1:0]       Ie24b89ee61bddac2f2bbf1b8b5dd437f;
reg                              I67c58e4de1a3413b77529f5374201308;
wire                             I3e9c216d05b6a9c1040616a42af371ff;
reg   [MAX_SUM_WDTH_L-1:0]       I27b99df87eefd6fcd484ec321bb73dc7;
reg                              I9ad9a905418216c83643eae11965f330;
wire                             I4902647240aca7d98844546130944322;
reg   [MAX_SUM_WDTH_L-1:0]       Iaac7f8ca30f4e74e1ae5016a222673d7;
reg                              I2f3232289260297dfb0cb36e42e459be;
wire                             Ia4c22694be7c5db34c1b875db1e91ff3;
reg   [MAX_SUM_WDTH_L-1:0]       Id3076c8e12f28723096148d8cf91a13d;
reg                              I58525519bd3b6773ec9ebabdf2764f69;
wire                             I0760280d5f5f23d9e06752908f0bbd96;
reg   [MAX_SUM_WDTH_L-1:0]       Ib2e36c2d0a51f5b953b9f368f11bb295;
reg                              I0e369759d6a2e5df5cd4fe6765ef8436;
wire                             Ic807e0ddc985cffca6a389b468aeae49;
reg   [MAX_SUM_WDTH_L-1:0]       I9ef5138c78fee50aeb2568def8bc62a0;
reg                              If155fcdeb6ebdce7305bf57a5e8fc426;
wire                             I9e3643f805ebd6623b9ab7ab41c41ec2;
reg   [MAX_SUM_WDTH_L-1:0]       Ic1cac944a0ed80e5b6e3821e8451045d;
reg                              I53e38457ad9a8a8244c9a2dd06034f60;
wire                             I0dcf2ac5c06f517ea62c1ccd5acd9298;
reg   [MAX_SUM_WDTH_L-1:0]       I915f18e8333d52f6ec4162fe35317d17;
reg                              I0cdf5ba9765cb28f2718129218794ec3;
wire                             I26879becf6ee094c9b8b4969c9377af7;
reg   [MAX_SUM_WDTH_L-1:0]       Idbcf9e41a431a42028cc99d6be0c46da;
reg                              Ic8e633425dff5441ceaa669bdd924077;
wire                             I3daa291236c162f58fdb9587a880dddb;
reg   [MAX_SUM_WDTH_L-1:0]       Ic46dd35355bcd4470886fbd416b3c75c;
reg                              Ie7efb37f21bcddfe6cb7969533bbaca7;
wire                             I2e150157b54bedd2bc6d31435e29af0e;
reg   [MAX_SUM_WDTH_L-1:0]       I0765c8beae32257c6c37dabd94cbab7c;
reg                              Ie5a9f440574d20f6047c0ce556bc8477;
wire                             If392bba16edcc39c846dc23bdf59f976;
reg   [MAX_SUM_WDTH_L-1:0]       Ibc002286423e5ddf50b8ea25ea1b3377;
reg                              I8fb0748ba8138a9188a557fcf752a055;
wire                             Id0838a2f54127e6e86536294821b8fd2;
reg   [MAX_SUM_WDTH_L-1:0]       I714b85ebaccb1e11d16d53cf6bcf65b9;
reg                              If6261c7d9d9c1b95edf08322eac2332e;
wire                             I3d11d3dc5ad053fd7a82b00d4ab4b180;
reg   [MAX_SUM_WDTH_L-1:0]       I864ca16e4e93b435a94fb012d995c7e5;
reg                              Ib9f5522d41ddd9087096bb10ce7f5e23;
wire                             I1f67b8b8a325071662e006b730b1cc8a;
reg   [MAX_SUM_WDTH_L-1:0]       I227ef7de18494a9f62b2e8cf37687840;
reg                              I686a59acf3c8d19e90c2060b7db4be8f;
wire                             Icd7c05e9200f346555aa6b82827ad164;
reg   [MAX_SUM_WDTH_L-1:0]       I535a78cff546aed9fbd1d79827d56fe6;
reg                              I73ba52dc87f86c76035540575994a224;
wire                             Id136b4b678027d89c31614cd5baa6282;
reg   [MAX_SUM_WDTH_L-1:0]       I90cf52bd1332ea1b955e8c193b670218;
reg                              I5947a59182e394e4b2f84b68ffd7bccc;
wire                             I08dad437a9b452f65231279ae25ab7e1;
reg   [MAX_SUM_WDTH_L-1:0]       If7dc2cec6ded3b32d42281d08e871513;
reg                              I006c14dc1c5be7dd3c5e1e5dcce08c21;
wire                             Ief01dd5ab84a9f9b05e48b07e0d1ed54;
reg   [MAX_SUM_WDTH_L-1:0]       Iee43875ccb00a79e67acbd3e12cb516d;
reg                              Iee841700cb259de93cbbfb47e828e1f4;
wire                             Iba8886370777ea357fd7c1e13bf03cd2;
reg   [MAX_SUM_WDTH_L-1:0]       I7aaad9fdd239670e028a896695c01216;
reg                              I71e36dabaef7951e59fc8b08da50003d;
wire                             I9e1e97a64e15a82443cc946178c11d52;
reg   [MAX_SUM_WDTH_L-1:0]       I4a992ed2550a3c5b346158ffe18c255d;
reg                              I323df8d18a73cd3947512f8a2c41b323;
wire                             Ib830e17254cac0158be2b443e3dd4d43;
reg   [MAX_SUM_WDTH_L-1:0]       Ib2eb28843cf201e8c6f8900b7029d42d;
reg                              I30604b84bad8b4bba6d340cf020ca901;
wire                             I819741033c6737000bcf4a07a78e0938;
reg   [MAX_SUM_WDTH_L-1:0]       Ic9a5b2c8aee24c3fbc7e92b8fdaed5dc;
reg                              Ib436620d6352c9ad5fa1d1fb5083de7a;
wire                             Ief41b57c092906a598c1cdcfea9b1062;
reg   [MAX_SUM_WDTH_L-1:0]       I6996efa8115f38da03518dcb7dd42a4d;
reg                              I0722db2c7497d82a0ee09a109f698250;
wire                             Ibea5db121c78f1b6d5288231ef59d04b;
reg   [MAX_SUM_WDTH_L-1:0]       I1c4bf7954b4bd5f4e9c176a3ae1fc28a;
reg                              I34fe1fee7604351d37636552ecb32d8d;
wire                             If9d3ee7956572ceb26e7d60077de7e00;
reg   [MAX_SUM_WDTH_L-1:0]       I55d0fd8eda9c128cacdebab55a8dda5b;
reg                              Ie9ca773a78e9592fc49a7c590a3afee1;
wire                             I46fa901f3606f4d2ef11e13cdf029826;
reg   [MAX_SUM_WDTH_L-1:0]       I02fcd92b426929f24b9a8c063a56c0ed;
reg                              I023b8de48fefb0b45bed81ada503d779;
wire                             I9918607fc0fdd746a6830800696a9439;
reg   [MAX_SUM_WDTH_L-1:0]       I3202a0ce45afe072eb955cd6e0789cd6;
reg                              Id0ac1f9bcd5fa52b3b0536f0c831d504;
wire                             Iac50ab3381392442d8e7f18bd9ecacd8;
reg   [MAX_SUM_WDTH_L-1:0]       I06c82466a2ca646abb62bcaad3d63748;
reg                              Ic5c3ce39ad2fd88b6a26e639e390155d;
wire                             Ie8bd9deffa3345851a9ff645b5bd1ddf;
reg   [MAX_SUM_WDTH_L-1:0]       I23af695cf96a03638f0c1ef719d8d530;
reg                              I80a34c662ed81f7d38d3055d470a1d1d;
wire                             Ia7d6b9edd50a4046aab863855f9491ee;
reg   [MAX_SUM_WDTH_L-1:0]       Ie20b7fc4110631c1da7de4c7f38e2581;
reg                              I0552127e741bcac86d4ef3994bf8830a;
wire                             If8c22f4e0850faaa35f617a99c827f84;
reg   [MAX_SUM_WDTH_L-1:0]       Ic6983ef65e0de21992fa0b90ddbdce9d;
reg                              Idef88c7c7169dae7b6d14e0edb17f47d;
wire                             Iee22d62b28aee7dfc6c9304c92214e55;
reg   [MAX_SUM_WDTH_L-1:0]       Ie7c2317cef621a89ad24c8b5bc79a39c;
reg                              I6f2e27ee85aad612520efe0e53f05aac;
wire                             Idd235ad7cda4d67de5992f50db3b8de3;
reg   [MAX_SUM_WDTH_L-1:0]       Ic58955d8604cb1a6a20a199372d44774;
reg                              Ia9afdb2578f40035f59aabad30a7e156;
wire                             I6bb6fc0f5773f1386ac5af0688f224db;
reg   [MAX_SUM_WDTH_L-1:0]       I8198473d2a666821cdf398dcf1b0fdc1;
reg                              I3c07ba2d2d09f45d52fbfe66bc54975f;
wire                             If44d50ac2bf54fad8236b3fcd9484792;
reg   [MAX_SUM_WDTH_L-1:0]       Ic60bdcbc8a55bc760e52c37aa3030001;
reg                              I77a2d8cfbb2e6f050545e2865b514205;
wire                             I9039a46d1a19d43e6c1cb3f0c162efb1;
reg   [MAX_SUM_WDTH_L-1:0]       I987cca9a9fcbe4b617a7e524476431be;
reg                              If126c59dab3d743d2451279fc184182d;
wire                             Ib3c48b1a31a7198cc8d4fdd10d0c2db8;
reg   [MAX_SUM_WDTH_L-1:0]       I765c7209f3c7173362057fdb60aab732;
reg                              If745dbf2f0d756857eff51da036067fe;
wire                             If37efa97b30f1c80267e986fc90f759b;
reg   [MAX_SUM_WDTH_L-1:0]       I2c117c8ea4060a5094453cc6140c9bb6;
reg                              I22231ac2204ad703262885231f7451e8;
wire                             I42e35cda79f11acac889996660ec32ab;
reg   [MAX_SUM_WDTH_L-1:0]       I56a6be4115d52bd49fc003b164fbcdb0;
reg                              I4e1e119c87f56b39ec6ddab9b160430d;
wire                             I0ac3076614fbc543f41c76c6be389a37;
reg   [MAX_SUM_WDTH_L-1:0]       Ib834a7e4f3a491e351e2e49d809d2448;
reg                              I9d9cc96988bd0af2b2c8682af3779794;
wire                             Iefae454b50cfb5b83c8016d5826e7670;
reg   [MAX_SUM_WDTH_L-1:0]       Ifdcb28209b39b8d99c2eb00a72921a75;
reg                              I027210d36e2ae38a39746ac6fde3129a;
wire                             I86cd5db563b397776c52a89f0b44e442;
reg   [MAX_SUM_WDTH_L-1:0]       Id721a94e50637fa39c5bf6124ecfae6f;
reg                              I28e32abf786d964b95d72bc17425a90f;
wire                             Ibbf7f6c104c9f3163fc8d6b8a33ff5fe;
reg   [MAX_SUM_WDTH_L-1:0]       I72ee7b62c165dc693cc6b5185970f7f5;
reg                              Id29266756e91fa3c40480f9cf22f1671;
wire                             Ife8ac54e4431329086b20d2111eb4f28;
reg   [MAX_SUM_WDTH_L-1:0]       I564ae36637e0cd6a8a06289e95823572;
reg                              Iad31d6f7d366c849222593883210e817;
wire                             I38c2a0e463853ac84b1f4e5c92f44243;
reg   [MAX_SUM_WDTH_L-1:0]       I085e99650c86078bf02f1b2aed141add;
reg                              I495d2cfe02637adf0bde6dd48201cedc;
wire                             Ib73515d47a61e4a795005e8ae6bb2968;
reg   [MAX_SUM_WDTH_L-1:0]       Ie4e63cba44dee9885eeae32cc844c3f5;
reg                              I544225b6c571710d59f804f082f475c8;
wire                             I48b52a0f686c64c91c6ef4b1ca47593f;
reg   [MAX_SUM_WDTH_L-1:0]       Ic054b062712da78ddd4a148bafeb1a0d;
reg                              I6f7ff2aeffdfe5bd4090ecd655ff5aa2;
wire                             I9ed8d0fadbdab4e176b2d03549e41c91;
reg   [MAX_SUM_WDTH_L-1:0]       I81b01fc018ad1c79ec03a123763e95d9;
reg                              I1783da96203ac6a00cd2e8f2dfe1ac34;
wire                             Ibed24a9317d456b1a27bf71649c9a751;
reg   [MAX_SUM_WDTH_L-1:0]       I1d38ff144c3dcfe4c04778e50a044d5e;
reg                              I00ae9e980c05d6d55570d92582a80410;
wire                             If6b0b5b913b2f16e0354a62459f87487;
reg   [MAX_SUM_WDTH_L-1:0]       I2e31a90886f87907d19d0c034caeee9c;
reg                              I86282458466a079a1063e068011d58eb;
wire                             I6cf5556c5887ad4d2f85b26aefe2aabf;
reg   [MAX_SUM_WDTH_L-1:0]       I7c48130cd79566b1f1e30b7c709ee5cb;
reg                              I7dcde2729bcd8e63b86dcac06325887b;
wire                             I4fa8769d910cc70e158a0b649ce1e1d4;
reg   [MAX_SUM_WDTH_L-1:0]       I3868c6ed60d1f0ef9d3ad98e91931acf;
reg                              I31ca3f6f5d61b73718bbd9c19f7fd53b;
wire                             If25316f70adbd92abb74b4338c63d7d0;
reg   [MAX_SUM_WDTH_L-1:0]       I7fa57873a108e5894f837bdf45979b8d;
reg                              Ie01688869a15f6b506bc3fbdea78b6b0;
wire                             I38b3f467871a1646a7694cc6433b5c8b;
reg   [MAX_SUM_WDTH_L-1:0]       I59d4025a86d065a84741dafb86b50cbd;
reg                              Iff748fa3440e5d0f80969f64b10eca98;
wire                             I0c7ee025ebd05956c96fd50885d627c6;
reg   [MAX_SUM_WDTH_L-1:0]       Ib28a3fb3dcdea36c883c88b017fefa56;
reg                              I85018196561b6ef22994dfff7e3a8b80;
wire                             I680660d6ba504eb445d2588ecfa046bf;
reg   [MAX_SUM_WDTH_L-1:0]       I91e4dca55e1a5d1d8ddee5c3bd1048bc;
reg                              Ifff25101d23e8e0ac43d5f0507a34217;
wire                             Ia861785bea48073ffcabfd97a16890de;
reg   [MAX_SUM_WDTH_L-1:0]       I55dd62b8ff91323075533e896207c1e5;
reg                              I261ed926e2e82b283ac24970f546a5fe;
wire                             I8619e41804844cd4d98818cb8387c3a7;
reg   [MAX_SUM_WDTH_L-1:0]       Ia30ca84355bb976cd045e969b2862856;
reg                              Ibf081c14165822b88553a913ba320016;
wire                             If916ac75b729dfffab3cf6b0029197ce;
reg   [MAX_SUM_WDTH_L-1:0]       Ifa1359651fd7e160301261bdbb81b02c;
reg                              I595bd58339ea7427b88385a62835aab6;
wire                             Id4f85daa963c656cff69ca2a821247fa;
reg   [MAX_SUM_WDTH_L-1:0]       I0b465f693268f6f56f52d41165bf66ef;
reg                              I41b82d4c805471097a0dd4f85615f990;
wire                             Ic39575e662d7843dcd7418a7e8cc4a75;
reg   [MAX_SUM_WDTH_L-1:0]       I3deffa3a53b31688f28dfbfa66571d0c;
reg                              Ie07ed8367e7b83324c539bddcb3b1dfd;
wire                             I7c445b4e53ebe960faa00a46e00d66b4;
reg   [MAX_SUM_WDTH_L-1:0]       Id40c9857a5bb6c8cdc616fe68d8dc39d;
reg                              I67ba6804ea940c34c7c588832272581e;
wire                             Iede71af4d6ced16d85e2576f035cc712;
reg   [MAX_SUM_WDTH_L-1:0]       I26754124b13858a3b925cddca5cd8c5b;
reg                              Ifb2d4794b0630c3cdecb6cd2d2b1b384;
wire                             Ifffbd3dc45d11e43be5de5a276300bd4;
reg   [MAX_SUM_WDTH_L-1:0]       I2ebc1a7d32a5457de4d35b6bb25507d1;
reg                              I9c6dda8e9e0d7e69032a1fb40684c87c;
wire                             Ib7be21d644d545e6671098d3d8622fe0;
reg   [MAX_SUM_WDTH_L-1:0]       I77bf5b03fa300d1dbf8df5ca4acbed14;
reg                              Ie7d857b468dedb6b7a73fe918332ff1d;
wire                             I1bcc55c2c22b349f421eac34341487c4;
reg   [MAX_SUM_WDTH_L-1:0]       I6c1c1e404f92fc80495e8e5d187934a6;
reg                              I34662a12c505be8abbe01cb690d117d5;
wire                             I5117b588204bc017b2a94a6e1097df82;
reg   [MAX_SUM_WDTH_L-1:0]       I126a2b15cdc34d88d17ebacb3681625f;
reg                              Idc13433074453a726e7a35789d7d27d2;
wire                             I7c6e35ef749c858168d55bcabea9078b;
reg   [MAX_SUM_WDTH_L-1:0]       I9c5ec8e21febe3ebe00c53ac8b21d1f1;
reg                              Id16d40761b18218d4270c00db6d4eca2;
wire                             I84a9bd349a6cd85859437ad4f9e70693;
reg   [MAX_SUM_WDTH_L-1:0]       If27eaa7cc4d1b5d2b7a962b48f0919df;
reg                              Ifac93c987a8fb9726d85b77a2e4c8bba;
wire                             I27b66137a39cb30b8059289cf98f8a19;
reg   [MAX_SUM_WDTH_L-1:0]       Ic15f443512d68537f9764a3ba88334f6;
reg                              Id742302a78483bbb2852b002262ed33d;
wire                             I89b31cd7510ff82f89398b8682f040f7;
reg   [MAX_SUM_WDTH_L-1:0]       I47b266262fb5a98f66706f460f1248e6;
reg                              I2f87df8d48fe83aa0ce493d69aaa3d88;
wire                             I801f6e47b9e4f6b6acfaf6f8369ea217;
reg   [MAX_SUM_WDTH_L-1:0]       Id301f31702270a4f8e9964e3a75e3d62;
reg                              Ic4bb880cb9f8d5a6d1cbbdf7cd205470;
wire                             I6f7db7eb1e5bc6d08ea9059ef7c31949;
reg   [MAX_SUM_WDTH_L-1:0]       I097ba3ae5a0232ae6aa35478635640b3;
reg                              I369ea36c9da8f4c9b93ee70f8d4c149f;
wire                             Idd01178431a1c4a53be45095dc897c33;
reg   [MAX_SUM_WDTH_L-1:0]       I3b65eb49005aee57f61279c5a172d158;
reg                              I17f6c250d2d07a58ddde6d232a1ab5de;
wire                             I64ae03b30dd467619e71498ce8126df4;
reg   [MAX_SUM_WDTH_L-1:0]       I8573059885be4373531275502affd59d;
reg                              Iba5b23512434eb51ec8679a798273551;
wire                             I36eba1bdcf4eac1c5c4b458515ed3f6e;
reg   [MAX_SUM_WDTH_L-1:0]       I627f9d9ac0c07ded7306fd14773fbee4;
reg                              I91a06282a09b01980f2e7be4ecd3a982;
wire                             Ibb1a5ae8240913132795df9605e82ce8;
reg   [MAX_SUM_WDTH_L-1:0]       Ib559f45098803b21622fa96ade885abc;
reg                              I1b928fa95275de94960b3e2b4d67338b;
wire                             I597865149cd8d3e173f8aed514cec357;
reg   [MAX_SUM_WDTH_L-1:0]       I10e294379879538ecbf65fd423e7355d;
reg                              I6488c30acdb3b47d4d4ee7b5947abdfe;
wire                             I667f0a049c87ac48820b60b2346de1c4;
reg   [MAX_SUM_WDTH_L-1:0]       Ice861034cd3b2f3847f325dbc9f52d08;
reg                              I29a436013f98b750df592eb7d26d0d1e;
wire                             Ieb1c4ec26a969a2c1cb60e0d1c67b5cf;
reg   [MAX_SUM_WDTH_L-1:0]       If201eea7e0023bb17fe41dbb4b5ec076;
reg                              I6fb12e6f50ffa6e94c9d43a22681702c;
wire                             Id3293a3ac3bb53134fade82ddb8aace1;
reg   [MAX_SUM_WDTH_L-1:0]       Ib15f9bf401d734008d6a2b9a00c572d1;
reg                              Ib3f42f17505d5c091c8c924bbc26d117;
wire                             If7ed4187de370efdc1b9798bb6b05232;
reg   [MAX_SUM_WDTH_L-1:0]       I581f4e137ec21e639eec32a1675f4750;
reg                              Ia4c22a118187d5b2dd154a4371dc06d1;
wire                             Iefc40b941a682059aca6ac8abffe1cfb;
reg   [MAX_SUM_WDTH_L-1:0]       Ib7ff7b93c88fc8d9bcd915f0c678acff;
reg                              I1a87822c50f6a0ac5a5e96021ad49fb3;
wire                             I746ebc4b00c09f116eb087dfed4bf89a;
reg   [MAX_SUM_WDTH_L-1:0]       I34dc9dff97e78a2d711f75675944b0d1;
reg                              I6addbc7c163ce97b3482277e76c5feaa;
wire                             I69683a0683ab00462065f6c3069fb6f3;
reg   [MAX_SUM_WDTH_L-1:0]       I8bc35065fe56bb75e6595937aaf9ef2a;
reg                              I124c4374f19808abbdc401a3b85aec67;
wire                             I183ad57174d779bab96973fc5ba5efd9;
reg   [MAX_SUM_WDTH_L-1:0]       I1822ab8ed690d872380ef820dc4282fe;
reg                              I162653d33938a4553978b08df208228b;
wire                             Ic4e5558ac995583236747a83b3f54f33;
reg   [MAX_SUM_WDTH_L-1:0]       I1a1965726584c6c91a7e20de63f0fce3;
reg                              I291a3bbec5669b8958c0ded154af1f89;
wire                             I12899b73e235f01bce4137c479f6b300;
reg   [MAX_SUM_WDTH_L-1:0]       I08c5dcac6674c1671b85d07a55a005b0;
reg                              I53a1d11cce6e036ba3a23dcc29d1cc3e;
wire                             I8dc3438a0d2b1c000f2b581f9a7ee588;
reg   [MAX_SUM_WDTH_L-1:0]       I40d67287bf525ab2696c30755d6babd5;
reg                              I5fda5f3c582bb88cb7de87298d15194a;
wire                             Ia589b25714c687f50bfa26ead5cfae55;
reg   [MAX_SUM_WDTH_L-1:0]       I60dc8e5b6204e3a5fa32e79c5cceae94;
reg                              Id3933d661bcebbc3584c9e437c96c89d;
wire                             I7e4263d478638c2f3127394328deea11;
reg   [MAX_SUM_WDTH_L-1:0]       I0074b447046d75787aa872d8167171aa;
reg                              I0d38a30070a5ae3e879c357c3dde88ea;
wire                             I1c432aa61cf7d02567ef990929a15696;
reg   [MAX_SUM_WDTH_L-1:0]       I384965816ec3b915b9b623ad68fcc4c9;
reg                              I928993ece796543b23fb83df8c250845;
wire                             I64531ff978fb8892605f2b0dd8422873;
reg   [MAX_SUM_WDTH_L-1:0]       Ic0e2656bee7174384f7f952dbb9da619;
reg                              I226f8490438d72f58c43377c8e60fc34;
wire                             Ib8c44be17e150cbd0b49d41c060f95f1;
reg   [MAX_SUM_WDTH_L-1:0]       I4cc3b0546ddc14d78da59e4981a77b58;
reg                              Idaefaba16ce80e24f16df683cc83d759;
wire                             Ic45b89f2b51ee014d9a0fb19a7ed7619;
reg   [MAX_SUM_WDTH_L-1:0]       I7b680caf7d0d94114fae1d96ba374e68;
reg                              If1da75cd8208f606c1b121f441685cbb;
wire                             I338e32162153b4ed5d991c44c38aca27;
reg   [MAX_SUM_WDTH_L-1:0]       I7f8986a922c03b6afb5786cd2e1d5288;
reg                              Ib63f66960a3981879aad950588ea14be;
wire                             I06c60ff1b8b447112b28f71eb9e3944d;
reg   [MAX_SUM_WDTH_L-1:0]       Ie7814643e3833736c0f54b39f91fe792;
reg                              Ia2c2ecedc809186e3f9224a9aa4bf385;
wire                             Ic2cc5a2da05052c4a68cadde2745b44e;
reg   [MAX_SUM_WDTH_L-1:0]       Id1f0c95b85ee041818da4fd9b5466c7d;
reg                              I1fc189d6e8a90cc0033c6e690916de83;
wire                             I8073ab2d9dc1d68d0bb4694ff206995f;
reg   [MAX_SUM_WDTH_L-1:0]       Iefa8421c0c908de69fccffbe22f40911;
reg                              I7fa18d2c7159b9fda8957384ebca5700;
wire                             I6aec90f4d15da8590fe767c4facfe19b;
reg   [MAX_SUM_WDTH_L-1:0]       I4319bf1bbb31debc7f58157b75025134;
reg                              I7ea0274f5b34aac64a17fa9171201a5a;
wire                             I39a8cf4c424841d2b367cb3a1207fe03;
reg   [MAX_SUM_WDTH_L-1:0]       I4a349021efeeda16b646979a959bff6e;
reg                              I8d26db6f54d068f798e2951701aebed1;
wire                             I031f3e2575360f675bed8e87a71755d7;
reg   [MAX_SUM_WDTH_L-1:0]       Iaae0c136077ecc36fc382a76abd550e7;
reg                              I8fb8a6e1ab4647e8e1dda4da8b3ef3c6;
wire                             I40feba64660df64a02c3df651a2ca26c;
reg   [MAX_SUM_WDTH_L-1:0]       I4a442564148493664046e7b38cc6cfe4;
reg                              Ie4821dad77dec0567d64f7c1de7710af;
wire                             I985f121a0212a4d64ca4a47c1c210b40;
reg   [MAX_SUM_WDTH_L-1:0]       I12cc5eec3de8ceb3ca084194d430d9a5;
reg                              Ic4d741a90fcc86f31eb3567d028eb27f;
wire                             Id4ce64c9f467d1b1c4bc9099ab855db2;
reg   [MAX_SUM_WDTH_L-1:0]       I56db71b7df11c35080cbaee80c389c59;
reg                              I1d2641b8888a0f7b4b78cae16779da75;
wire                             I01c6d49bf9698d7621a545481b129692;
reg   [MAX_SUM_WDTH_L-1:0]       Ifd1431230378775456efa4bdd5bfc397;
reg                              I48badf0536ab133751d4be1e0450fd81;
wire                             I73164ee0df8db9282850f1b325afc7ae;
reg   [MAX_SUM_WDTH_L-1:0]       I6f0cef6d870e38e5ba192463a3920818;
reg                              I043ba9e5157ad18a4e466df0540b79ba;
wire                             Ic985d004f7feb36aaa6415dc7365e617;
reg   [MAX_SUM_WDTH_L-1:0]       I3ee87c05f23571b687611fdce84a1b91;
reg                              Ib9760b69084b2d4a3a93126e5da0f20b;
wire                             Ia09ac88781a570aead25d43447ff9afc;
reg   [MAX_SUM_WDTH_L-1:0]       Ide521f7523b897bb6fb747202f730ac5;
reg                              I4978a011cb09d68ac2850e1f515d7e88;
wire                             I17cb6dfd1374c74d63862703fa6665ce;
reg   [MAX_SUM_WDTH_L-1:0]       I314b64e5fbbc14807fd7fe3c7bca101f;
reg                              Ib09ea18232dfca23f3f139438e6cb800;
wire                             I6c05d39d4c7a50f019474562f741e591;
reg   [MAX_SUM_WDTH_L-1:0]       Id5ad2e12b160bc6a9f96f2524f849c8e;
reg                              If29c61ebd2b452efe995c212a76a77a0;
wire                             I413638a340bf1e686e718453f1b243b6;
reg   [MAX_SUM_WDTH_L-1:0]       I2b2bf6d4e879b8f53b02f94f1e964344;
reg                              I60fa2e2b5dd8b0a99612d2f2f6c5c740;
wire                             I904a05d4a23c6d15438654f937811877;
reg   [MAX_SUM_WDTH_L-1:0]       Ic60cb038b4b90d8035059b1e06f8d765;
reg                              Ifc9b6cc64f5bf8bc685911bb28884a0e;
wire                             Iab36b17e472fde9a92c4dc5ebb75ca6c;
reg   [MAX_SUM_WDTH_L-1:0]       I707e2d6d9807076bfc91417fb9e198e6;
reg                              I1aeaa36994ba29298931735d5a1237e0;
wire                             I4d265ef808b1e19fb1dcef26a6dd4204;
reg   [MAX_SUM_WDTH_L-1:0]       I49f5797b92e17562e6dfde42c20c7a37;
reg                              I415ed6a9802acf39be10b220ddb3ff66;
wire                             I535542d9580a449d24a712ef814d5e58;
reg   [MAX_SUM_WDTH_L-1:0]       I0a9f0274dc61d574c40e0e2048fb0b9e;
reg                              I1c06321ed28c991ad2aa8a3725769dee;
wire                             I82298047310dc4da0ea3762c6a48e07f;
reg   [MAX_SUM_WDTH_L-1:0]       I53ae3de5769255a9e69a2ae690d44ba9;
reg                              I198d5b5bf8f39f9bd6b2f4c993fd58ca;
wire                             I761dfdefbc96fec3c2ac79f0a1de18b7;
reg   [MAX_SUM_WDTH_L-1:0]       I1390f0ff082dbff11a64cdfcbe1b681d;
reg                              I3bf64d0a85c83de954a286e6afa8f727;
wire                             Ib68e4d694df8e44519916724104f7962;
reg   [MAX_SUM_WDTH_L-1:0]       Id2f8816659d3881ee1b1d14668a53a08;
reg                              I897c7fc822d490f69b531a8f749815f4;
wire                             I3284ce21b5d114a7127917f8b261b21a;
reg   [MAX_SUM_WDTH_L-1:0]       I286bacc5a8a77b89cb99dbb00962555b;
reg                              I6c7cb10db83156b49d46fab38d0f9fc5;
wire                             I30b857065185101e8e4cb0270e747cae;
reg   [MAX_SUM_WDTH_L-1:0]       Icda8e8a6ba7607752ed282114a542b67;
reg                              Ie47af3b071351ec683abe28b7fe2b642;
wire                             If9be63889327fc1b68abc628c9a0a78d;
reg   [MAX_SUM_WDTH_L-1:0]       I2da4a59f9a6bd71af95790a75b172df0;
reg                              If2dd4df3af6446c05da4afdaa7e92cab;
wire                             If0c3ec1e3a80a23b2506621ec2d9f02a;
reg   [MAX_SUM_WDTH_L-1:0]       I1bcf01b7fde13919f5d7c4df4483e61c;
reg                              Iabf085ea078abe8748810e81a6d03cac;
wire                             I2842882109b7ef022421ab185471ab33;
reg   [MAX_SUM_WDTH_L-1:0]       Id5f000c37734979d057f7887739a5615;
reg                              Ia2ae348906a599a4d327ff1419315afb;
wire                             Iecb13253abbfb0a891a4e526f05841f3;
reg   [MAX_SUM_WDTH_L-1:0]       Ibccd7142ba951dadbeca13178458bb3a;
reg                              I18df34aea04ea7dc99fc918892bf8f0e;
wire                             I899cefdf3938be01e93d011e046c1e49;
reg   [MAX_SUM_WDTH_L-1:0]       Ic1fe6b93bc8d517686ba430d3d1fe7ab;
reg                              I910749abcd809e1c730f27fb5e1ddab1;
wire                             Ib96a9bf253b178aa920a63c8493932fb;
reg   [MAX_SUM_WDTH_L-1:0]       Ib1c8d1d733e91f052f6d6824e734b1e3;
reg                              Iae95ea2f32f53a5060c0199c8196d681;
wire                             I5f534382562a3394100cdadb3ad1e0be;
reg   [MAX_SUM_WDTH_L-1:0]       I08348d0a177e264af1a4769422878a06;
reg                              I8c3d927ec93e73c5bca489a2f2b43f55;
wire                             I137e343ba2386bbe31813bbe37e87dd9;
reg   [MAX_SUM_WDTH_L-1:0]       I2d2c2997dcc5167fc6ddc1e90f0ebc49;
reg                              Ib41ff881898782965734bb0cc333be79;







/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic05b492587d8d5083e8570900995293a;
reg  [MAX_SUM_WDTH_L-1:0]        Ic93835a022c46b7aa00a465c407d7da2;
wire [MAX_SUM_WDTH_L-1:0]        Ibee9ba58404f1adb9e4e8e6f822a38c1;
reg  [MAX_SUM_WDTH_L-1:0]        I2e30088bf29cedd7debc15b1e6ec4ada;
wire [MAX_SUM_WDTH_L-1:0]        Ifab38317b76e52f9d9d64bed976e2cc5;
reg  [MAX_SUM_WDTH_L-1:0]        I38f512bfb84094d1e92a10a345d5505f;
wire [MAX_SUM_WDTH_L-1:0]        I86195d9a1da88ffc163298c54401039e;
reg  [MAX_SUM_WDTH_L-1:0]        I1e878f00f056f637625cb013a93325a8;
wire [MAX_SUM_WDTH_L-1:0]        I27c02895bfd59c762d5c7a725aa5cefd;
reg  [MAX_SUM_WDTH_L-1:0]        I25db27464b31fee41ccd7a3cfe4d403e;
wire [MAX_SUM_WDTH_L-1:0]        I60de515e03218ac363566ce7b92f5034;
reg  [MAX_SUM_WDTH_L-1:0]        I19417a224c5cdf1211e9790aa29c4c5c;
wire [MAX_SUM_WDTH_L-1:0]        I9b75e7451fbf27c3645bebbdba234996;
reg  [MAX_SUM_WDTH_L-1:0]        I16dcafa854ea9c67d8a080feb2ba9166;
wire [MAX_SUM_WDTH_L-1:0]        I056c79002bbba10ddee2448e36dc7478;
reg  [MAX_SUM_WDTH_L-1:0]        I7f63338eee2663fbe61fffd248433310;
wire [MAX_SUM_WDTH_L-1:0]        Ia5db5f66b7fb04e2344abff9b4f75404;
reg  [MAX_SUM_WDTH_L-1:0]        Icb1e3c56c8729c32d43c69710e345db2;
wire [MAX_SUM_WDTH_L-1:0]        I250898de23a8793f0c21eb333d61af53;
reg  [MAX_SUM_WDTH_L-1:0]        I6ece8e3c1e89613879336936f77d732f;
wire [MAX_SUM_WDTH_L-1:0]        I1320273c298c7953b3227b58439b54c4;
reg  [MAX_SUM_WDTH_L-1:0]        I72a646ae7e32a16af0f5930a6e95b36a;
wire [MAX_SUM_WDTH_L-1:0]        I49a036af196fb318309a43c150540a2c;
reg  [MAX_SUM_WDTH_L-1:0]        I7e72d119dd93a6ab05a23fde0a865866;
wire [MAX_SUM_WDTH_L-1:0]        If115c3e5f121363c2b8a6c14905aebe7;
reg  [MAX_SUM_WDTH_L-1:0]        Ied4fdf5805039cd2fcd042fd13755fdc;
wire [MAX_SUM_WDTH_L-1:0]        I5fcd95690fb291f9b95996e687de022c;
reg  [MAX_SUM_WDTH_L-1:0]        Id44c2293b765cff450dd1d747c47c1f3;
wire [MAX_SUM_WDTH_L-1:0]        I5f6f8a4c5c5ab4cf1f9c496795c41ce8;
reg  [MAX_SUM_WDTH_L-1:0]        I8f4ed02f7aeb823b745040f7f3f43ac7;
wire [MAX_SUM_WDTH_L-1:0]        I775180b845280ec240e4adf20605b8fe;
reg  [MAX_SUM_WDTH_L-1:0]        I6488b9b8f405d7d81a4874fab2678102;
wire [MAX_SUM_WDTH_L-1:0]        I642fe2c7978d7229d660431061a6f781;
reg  [MAX_SUM_WDTH_L-1:0]        Ifff612d16828ec907a348479e19ddf31;
wire [MAX_SUM_WDTH_L-1:0]        I3ce66aa6048542c81a89c28e80412e70;
reg  [MAX_SUM_WDTH_L-1:0]        I268262076f22bc6b1507bc8f91b98a0a;
wire [MAX_SUM_WDTH_L-1:0]        I436fc89b03a41f35b8d2ab89464d07c0;
reg  [MAX_SUM_WDTH_L-1:0]        If1f732841adb7c0cad1ba37c0f5fd517;
wire [MAX_SUM_WDTH_L-1:0]        I67861da88ed0edc52bb876287fc60261;
reg  [MAX_SUM_WDTH_L-1:0]        I0df8a24f31c027756d248c3bd1b9bf7b;
wire [MAX_SUM_WDTH_L-1:0]        If51bec96c3139419947f0442b0ad7281;
reg  [MAX_SUM_WDTH_L-1:0]        I8ef901e733b12e76412eb36684e2b575;
wire [MAX_SUM_WDTH_L-1:0]        I5e126994711cd1782fcbd2fb3eec3cdc;
reg  [MAX_SUM_WDTH_L-1:0]        Ia48916a02f68b1b8f5fc7fece04677bb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I44d2fe323e921ba0fd66c82a792302e1;
reg  [MAX_SUM_WDTH_L-1:0]        Ia37409944d9fdd3b16e7007e13d82a79;
wire [MAX_SUM_WDTH_L-1:0]        I875b53feb16dc1ac263e9d1c2552dd38;
reg  [MAX_SUM_WDTH_L-1:0]        Idd65f149afe9d5f63ddaf34b82b11e95;
wire [MAX_SUM_WDTH_L-1:0]        I651f168318d2ce4746ade3230e052ace;
reg  [MAX_SUM_WDTH_L-1:0]        If2886d560854faed32ebd8e33d868973;
wire [MAX_SUM_WDTH_L-1:0]        I00a65dc6a94fa280ec3aac7b04fd4aba;
reg  [MAX_SUM_WDTH_L-1:0]        I77778118bb3ea900c080754ff4c49c26;
wire [MAX_SUM_WDTH_L-1:0]        I38f5eb8d994476d2edb5fd71b7636452;
reg  [MAX_SUM_WDTH_L-1:0]        I7292ed752d8741594d757730950feea4;
wire [MAX_SUM_WDTH_L-1:0]        If0d9102fbff225bd3ef4f4e1aab2811b;
reg  [MAX_SUM_WDTH_L-1:0]        I68cfd7868e061793ee8a41e69e80219b;
wire [MAX_SUM_WDTH_L-1:0]        I09734a3840b1b01a467b075c65608f3e;
reg  [MAX_SUM_WDTH_L-1:0]        I667ead814b303fca64ef047bb8246b19;
wire [MAX_SUM_WDTH_L-1:0]        Icec563470fe1bec10dfa8d36561f6ed7;
reg  [MAX_SUM_WDTH_L-1:0]        I4f25c7edb12e868cb5532e42b4ba5133;
wire [MAX_SUM_WDTH_L-1:0]        Iaa82bbd78ea7acbc1949f7db44d339eb;
reg  [MAX_SUM_WDTH_L-1:0]        I5aed2d82717f359bb5ac5a0ab91b7beb;
wire [MAX_SUM_WDTH_L-1:0]        I1bf879a8671257cec876577804bd6ffb;
reg  [MAX_SUM_WDTH_L-1:0]        I92835fd54631deaefa7b214e2c4b9bff;
wire [MAX_SUM_WDTH_L-1:0]        Ifdb571f08bb8fc78631b0af95d6f5b68;
reg  [MAX_SUM_WDTH_L-1:0]        I67e067da565635fcff166e3a7d0c446b;
wire [MAX_SUM_WDTH_L-1:0]        I06117d4a9cec69582f336796f82af871;
reg  [MAX_SUM_WDTH_L-1:0]        Ifdb0f307b1b9458c0487a1574ccc094b;
wire [MAX_SUM_WDTH_L-1:0]        I23178a40d717727916e4c44fb8ea7de9;
reg  [MAX_SUM_WDTH_L-1:0]        I5c6b7d143e42fd3b8bcdb7d7ed4da2c2;
wire [MAX_SUM_WDTH_L-1:0]        Idd1454bc7f85ca3c184a20fd0864c666;
reg  [MAX_SUM_WDTH_L-1:0]        Ie679a21d0136a08cc5e6526e9f8d1843;
wire [MAX_SUM_WDTH_L-1:0]        Iee01a4b6a910ede0b61e2465d7d5d696;
reg  [MAX_SUM_WDTH_L-1:0]        I611942a72a5e12f6afaea6bde6699ef6;
wire [MAX_SUM_WDTH_L-1:0]        I383d6b1028ae1e4e2ea40cfa22043d72;
reg  [MAX_SUM_WDTH_L-1:0]        Ica9883c97f823a4491cbee5b45c43590;
wire [MAX_SUM_WDTH_L-1:0]        Ifde4b0c41d42daf9b134ee6c05db336a;
reg  [MAX_SUM_WDTH_L-1:0]        I8e6addfc61f5bfb7af74fc2993639565;
wire [MAX_SUM_WDTH_L-1:0]        I9f0b1952f54a14726de1d31a2302a95f;
reg  [MAX_SUM_WDTH_L-1:0]        I9d53619f10e2a426f7297bbf7c81158a;
wire [MAX_SUM_WDTH_L-1:0]        I3991c8d4f24af7dfb52a65f70c3ab2d5;
reg  [MAX_SUM_WDTH_L-1:0]        I8a055c27778913287ad951183fa0d4d6;
wire [MAX_SUM_WDTH_L-1:0]        Ie928ef6ba83900dca8b150428d713448;
reg  [MAX_SUM_WDTH_L-1:0]        I8f6ae5c80bb2f50084b5f5ee5ab0ffc3;
wire [MAX_SUM_WDTH_L-1:0]        Ic085f1faeb81e3027f909a7bd890d359;
reg  [MAX_SUM_WDTH_L-1:0]        I3db8b3a342e8e2f13a448246aa001c2f;
wire [MAX_SUM_WDTH_L-1:0]        I159df37fedc1447f6766308aa58ff70c;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbee0996ea0f5e16b1f711345be7f2ae;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I53491740a9877fcff56e6a3d8ac61643;
reg  [MAX_SUM_WDTH_L-1:0]        Idb777f1eb4c3cbba103b9b43f948ccf9;
wire [MAX_SUM_WDTH_L-1:0]        If9eba70be918197cc0bb2974f04c0687;
reg  [MAX_SUM_WDTH_L-1:0]        Id5e46b1f8844c7587f99d22170581a24;
wire [MAX_SUM_WDTH_L-1:0]        I2a30d44d2006f17582bb431e397d3874;
reg  [MAX_SUM_WDTH_L-1:0]        I67aadabd3cf49456cace7392a1e7a35a;
wire [MAX_SUM_WDTH_L-1:0]        I4b64bd561b279a17da4758a188a2f395;
reg  [MAX_SUM_WDTH_L-1:0]        Id5635595d6b7b6dd7e6d510a27ad6702;
wire [MAX_SUM_WDTH_L-1:0]        I93d5297fada8dfdcffed4b7b56ef9c43;
reg  [MAX_SUM_WDTH_L-1:0]        Ice783314a4868f0bba8bc3c5e3b65ae4;
wire [MAX_SUM_WDTH_L-1:0]        Ic6e5118343e784f89cd1d3ba03309f20;
reg  [MAX_SUM_WDTH_L-1:0]        Ib2d9b7f58cf571b904be02e6073f9b94;
wire [MAX_SUM_WDTH_L-1:0]        Ic5d76ee2f693c012e26dc17acb0086e2;
reg  [MAX_SUM_WDTH_L-1:0]        I61b6effae91ae4bdcce4550eb5cf0796;
wire [MAX_SUM_WDTH_L-1:0]        Id4ad545c42b5e4c8d5383568ad1e2013;
reg  [MAX_SUM_WDTH_L-1:0]        If5cf6e81b0e3b77f6a45f2555201acc2;
wire [MAX_SUM_WDTH_L-1:0]        I3a6030885679b87e44a54cdac13681ad;
reg  [MAX_SUM_WDTH_L-1:0]        I62fae5bf51588f28c3521715b834909d;
wire [MAX_SUM_WDTH_L-1:0]        I0791083d118ca9bf64108ec397af3d04;
reg  [MAX_SUM_WDTH_L-1:0]        If5cbdab78a4cf86b6285a400d0e0ac90;
wire [MAX_SUM_WDTH_L-1:0]        Ic683598c8ec40f18eed02cb89e8a8270;
reg  [MAX_SUM_WDTH_L-1:0]        I6e481cc49441c08bcd9fdcabbe90a000;
wire [MAX_SUM_WDTH_L-1:0]        I1fc9bb5cc8d38dd67592141a4dbf2532;
reg  [MAX_SUM_WDTH_L-1:0]        I3aa663be3dd604564ef68b9a2b9d7319;
wire [MAX_SUM_WDTH_L-1:0]        I7ec34dc5c899abcd284ccd637fccf4ba;
reg  [MAX_SUM_WDTH_L-1:0]        I8031632ee8700c63c207e2d6a6bdb630;
wire [MAX_SUM_WDTH_L-1:0]        I2d43f4939c3509b6e7e540d3da880c35;
reg  [MAX_SUM_WDTH_L-1:0]        If9be2701858da0bdffbf2dff7bcfd7e1;
wire [MAX_SUM_WDTH_L-1:0]        I385df2a645f7269a298cbadc418a54b9;
reg  [MAX_SUM_WDTH_L-1:0]        Ief209532f4cbf1c6a41bea414577f825;
wire [MAX_SUM_WDTH_L-1:0]        I5f90162de7034f414b502958f5ec9b3a;
reg  [MAX_SUM_WDTH_L-1:0]        I1c8953ad3f64f3c3cc506808aad29dab;
wire [MAX_SUM_WDTH_L-1:0]        I74353ed1bcc55b22f5d1f406b5069eaa;
reg  [MAX_SUM_WDTH_L-1:0]        I1b519d88bbf86cfb080a50ea0480a128;
wire [MAX_SUM_WDTH_L-1:0]        I6c28ab1bc42131e4ff3fa98c97990c37;
reg  [MAX_SUM_WDTH_L-1:0]        I5b8258f35d889071109216b464abb2a4;
wire [MAX_SUM_WDTH_L-1:0]        Ia7c2ca9384d0415bbfe92f719a8a4a2f;
reg  [MAX_SUM_WDTH_L-1:0]        Id9681d4e0e4d375f9279de115a4337a3;
wire [MAX_SUM_WDTH_L-1:0]        Ice3a20a00f8742bbf47a043b84964ee3;
reg  [MAX_SUM_WDTH_L-1:0]        Ib42144ece00b82debd70011724a29c91;
wire [MAX_SUM_WDTH_L-1:0]        I22bdaa7e1b37f335d3fb2232df587cfd;
reg  [MAX_SUM_WDTH_L-1:0]        Ic5717058a1815f63f164de1b1defe8cb;
wire [MAX_SUM_WDTH_L-1:0]        I1c41347158d76f8b81dfa334e99d07ed;
reg  [MAX_SUM_WDTH_L-1:0]        Iea41672f012f225d64d9c75b198c812f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3464039cbf8ed089ae1894998c1e156b;
reg  [MAX_SUM_WDTH_L-1:0]        I7a070bd014e1d2c5e55e5fcba88a5664;
wire [MAX_SUM_WDTH_L-1:0]        Ie7409851212f99a429d94460669686b8;
reg  [MAX_SUM_WDTH_L-1:0]        I4a0a8b28429b708363458c74230b0fc2;
wire [MAX_SUM_WDTH_L-1:0]        Ia575bcac8f127884a151a3a323763614;
reg  [MAX_SUM_WDTH_L-1:0]        If585e4075ac1740f3b141ae6a50200f7;
wire [MAX_SUM_WDTH_L-1:0]        I2a193624be6cb259f18ece3546c7ad21;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1a68cf09bb21a1629369fde87f51bea;
wire [MAX_SUM_WDTH_L-1:0]        If40ad1197633c486c3aadfa277f9ab51;
reg  [MAX_SUM_WDTH_L-1:0]        I72b8547125d0ad6c1ad39a68b55c818c;
wire [MAX_SUM_WDTH_L-1:0]        I629ddfee3e7d36b93b743e69b4c817d6;
reg  [MAX_SUM_WDTH_L-1:0]        Ie14ba4a8657740f9a8d057258db2cb09;
wire [MAX_SUM_WDTH_L-1:0]        I3469ef81705fd1534d6e5eb194f1e4b4;
reg  [MAX_SUM_WDTH_L-1:0]        I27490a69fb2a1f6f298639254c37cf9e;
wire [MAX_SUM_WDTH_L-1:0]        I832d0a2832b2c665f1261b07ac6f9f2f;
reg  [MAX_SUM_WDTH_L-1:0]        I49b9c212fbe74a5dd8b087e417296186;
wire [MAX_SUM_WDTH_L-1:0]        I3c2aa289ff967b044d6a37f75f048ec8;
reg  [MAX_SUM_WDTH_L-1:0]        I0a8e6f5cc8b6ea599b7605abe6479bec;
wire [MAX_SUM_WDTH_L-1:0]        Id2ea09c8febd9e18d231a5b069beb3cf;
reg  [MAX_SUM_WDTH_L-1:0]        Ib6d94b34d3886717e4016fec196f277f;
wire [MAX_SUM_WDTH_L-1:0]        I7b80623d743adcc50430ab9c8591ff29;
reg  [MAX_SUM_WDTH_L-1:0]        Id7e53d36da7171e036ebfc984dbcea6e;
wire [MAX_SUM_WDTH_L-1:0]        I05750cd7c98f3c9726b8bbf5cdc76844;
reg  [MAX_SUM_WDTH_L-1:0]        I2ec254d80fd0683d782302cf3839559b;
wire [MAX_SUM_WDTH_L-1:0]        I389c717754a30812dc8ae3c8dffa20fb;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbedaef61051d5df82cd6d55e05c80da;
wire [MAX_SUM_WDTH_L-1:0]        I8f151f04b124fa5023d7be59c9a43519;
reg  [MAX_SUM_WDTH_L-1:0]        I501336bb7ba172c05dd5840036e6228c;
wire [MAX_SUM_WDTH_L-1:0]        I29a6f7a5b1c0bcc988363bee48b6cdc9;
reg  [MAX_SUM_WDTH_L-1:0]        I8e5c4c6c63e42054359cee697cc0d026;
wire [MAX_SUM_WDTH_L-1:0]        If35ed918a1a2b59c5e0ba5f3e0a1a6f0;
reg  [MAX_SUM_WDTH_L-1:0]        Id3daa6db921871b752bf92366446afcc;
wire [MAX_SUM_WDTH_L-1:0]        I0816b1444f89b9c61ccfee1d16a72c1a;
reg  [MAX_SUM_WDTH_L-1:0]        Id8367ec60787bfad0da8aa76c6ed8ddb;
wire [MAX_SUM_WDTH_L-1:0]        I4a292e7bcef3cdaa716ceb101685471e;
reg  [MAX_SUM_WDTH_L-1:0]        I533649312ec995f1f9e514c59a8675b1;
wire [MAX_SUM_WDTH_L-1:0]        I1d6b3fdfa7d64dc0761ebcb6ad076bff;
reg  [MAX_SUM_WDTH_L-1:0]        I0621d0b2c83e70b4afd65eb9dca4b514;
wire [MAX_SUM_WDTH_L-1:0]        I3ce8fb414e9fa103854658db43291eb0;
reg  [MAX_SUM_WDTH_L-1:0]        I2ae01892a3cd0432618d7280b31daddb;
wire [MAX_SUM_WDTH_L-1:0]        I01d190427900b3cef55d978630d6e035;
reg  [MAX_SUM_WDTH_L-1:0]        I5ed8a2f30bd2ea269341c2267ae3fe83;
wire [MAX_SUM_WDTH_L-1:0]        I59a613f178a100a88f479d85e5f01cbf;
reg  [MAX_SUM_WDTH_L-1:0]        I2c819e7f62c0dc0aac650074b203163b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ife0377dc8109d89213ab27df5304e1e0;
reg  [MAX_SUM_WDTH_L-1:0]        I30e20b58913d6fbe5817e1956ba8e570;
wire [MAX_SUM_WDTH_L-1:0]        Idb55c5acb92ff1b590670da114d3c668;
reg  [MAX_SUM_WDTH_L-1:0]        I1b922bed7f3c4a6705f3ce7a885a68cd;
wire [MAX_SUM_WDTH_L-1:0]        Iefdc7b1d3aea42c3ddf9645510803a98;
reg  [MAX_SUM_WDTH_L-1:0]        I2f65f0917713ecc8585392d3b557c1bf;
wire [MAX_SUM_WDTH_L-1:0]        Ieae82f715fb1dc2d6d173f82b1547c35;
reg  [MAX_SUM_WDTH_L-1:0]        I3301533e7d9e527118a67c462f1b4357;
wire [MAX_SUM_WDTH_L-1:0]        I18a9e19a2c41be29621e5da6a2b08e3e;
reg  [MAX_SUM_WDTH_L-1:0]        I52a88bdb1f03da82730f7579b7b5305d;
wire [MAX_SUM_WDTH_L-1:0]        If4bfa23dd5ba282c7c9445769eb865f2;
reg  [MAX_SUM_WDTH_L-1:0]        I644c730662b3725d26cd46fb46106104;
wire [MAX_SUM_WDTH_L-1:0]        Id9717e06ce4a9b03b8430559671918d7;
reg  [MAX_SUM_WDTH_L-1:0]        I3da3e36c76c4123bec6879bccb39e933;
wire [MAX_SUM_WDTH_L-1:0]        Ie54acd665004eec584ab9ff50df3961c;
reg  [MAX_SUM_WDTH_L-1:0]        Iebde55cddc8170f7dd8855ea55eff0ce;
wire [MAX_SUM_WDTH_L-1:0]        I16c418af5cc92780b28cd56e8baa825a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie673e2d92a7090b2fa1c5e14a2e03be3;
wire [MAX_SUM_WDTH_L-1:0]        Iddb359180e3925dcf7081ba0560c27da;
reg  [MAX_SUM_WDTH_L-1:0]        If90afe75714f8660ad0eb9f9ea06cd6b;
wire [MAX_SUM_WDTH_L-1:0]        I354ac9e0f361928cf5cc7aaf22fd9622;
reg  [MAX_SUM_WDTH_L-1:0]        Ifd96e3a6e0050c30a4308328cfecb21f;
wire [MAX_SUM_WDTH_L-1:0]        Ibf2b259738d54319e3af570db254a79f;
reg  [MAX_SUM_WDTH_L-1:0]        I68b92cc2d83e9a718edd2aea82314016;
wire [MAX_SUM_WDTH_L-1:0]        I07150b2eb1a5818fe98aa210cb6e8221;
reg  [MAX_SUM_WDTH_L-1:0]        I6bdbb92363f0e072ed04654e9aad17a5;
wire [MAX_SUM_WDTH_L-1:0]        I5dea5fdbd4e09be8fd264360ae399b32;
reg  [MAX_SUM_WDTH_L-1:0]        I87a4267db59b97ef1b9bca8743cb0322;
wire [MAX_SUM_WDTH_L-1:0]        I9c52550c142c131371199bbf8bc08c01;
reg  [MAX_SUM_WDTH_L-1:0]        I44eacb2bea725efab7c0dd560279f0f8;
wire [MAX_SUM_WDTH_L-1:0]        I72d86068a1d9bdfe04f6ebe9afcf980f;
reg  [MAX_SUM_WDTH_L-1:0]        I87a2736466c5ee62b7cc55f17e715ffa;
wire [MAX_SUM_WDTH_L-1:0]        I412dfb474dbd41f407bbd57b0dd75a4e;
reg  [MAX_SUM_WDTH_L-1:0]        I7a66c7713ba126fdc24940cd92f7e10b;
wire [MAX_SUM_WDTH_L-1:0]        Ie759523643b0c4becb96025e66635b3b;
reg  [MAX_SUM_WDTH_L-1:0]        I1f11c579f34c41aade41c53f53468057;
wire [MAX_SUM_WDTH_L-1:0]        I1ef0aa04ba8b896c7ca95c10513b0ecf;
reg  [MAX_SUM_WDTH_L-1:0]        I651a438f70583d476ae10f066e035435;
wire [MAX_SUM_WDTH_L-1:0]        I880964445bdadb87455b7f8a865fa0e8;
reg  [MAX_SUM_WDTH_L-1:0]        Ibdf17fa73794c846e15fe0a915b071e5;
wire [MAX_SUM_WDTH_L-1:0]        I145bec82b2f3234d2299ea32c9cd32ef;
reg  [MAX_SUM_WDTH_L-1:0]        I76d3221fbcefc0ee08655f7ba4919f3c;
wire [MAX_SUM_WDTH_L-1:0]        Ib045b4ad82a55c17dd36f29467d49f36;
reg  [MAX_SUM_WDTH_L-1:0]        I3458f69c90ea8b20b3d1f67e9a13ec2e;
wire [MAX_SUM_WDTH_L-1:0]        I7a195d3fb06596483191024720bfae2c;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2d6e9e1e92a30c7028af50ddfbb9bf9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib84c4b8d94ce1e35ab220224ffedf4e5;
reg  [MAX_SUM_WDTH_L-1:0]        I66c91b5133d9812a03daecc0b14211f8;
wire [MAX_SUM_WDTH_L-1:0]        Idd54eedf955c30f097484bd789eaa3d1;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb5986949e88167526d9fcfe07b417ca;
wire [MAX_SUM_WDTH_L-1:0]        I123677fa899ce173a83101d91990014a;
reg  [MAX_SUM_WDTH_L-1:0]        Iedada801ca6cd173ee523ef335e91ff6;
wire [MAX_SUM_WDTH_L-1:0]        I26617d3c93a1f4069ee6fb732264d935;
reg  [MAX_SUM_WDTH_L-1:0]        I4e2722e547586da7565b2d91a7fc91e7;
wire [MAX_SUM_WDTH_L-1:0]        I00410cf0d9a85b1fa2f70212bed15642;
reg  [MAX_SUM_WDTH_L-1:0]        Ib321a8ceda62c64ab25dc1c718301bda;
wire [MAX_SUM_WDTH_L-1:0]        I28f355e643584a4ab8d55777aa26fa78;
reg  [MAX_SUM_WDTH_L-1:0]        I58daeebec4873e6c1c07c090ff81235c;
wire [MAX_SUM_WDTH_L-1:0]        Id21bc865cd2de83bced952fb9c25f11a;
reg  [MAX_SUM_WDTH_L-1:0]        I3f103fbbe49c86c9db46129bd4632cab;
wire [MAX_SUM_WDTH_L-1:0]        Ib6fbb4e2ef502ae86dc697dccfe035a8;
reg  [MAX_SUM_WDTH_L-1:0]        Id6697ca17f1bd6ddd112951b9d89a8ea;
wire [MAX_SUM_WDTH_L-1:0]        I2b0c304769c917cc6acc0855ada30c54;
reg  [MAX_SUM_WDTH_L-1:0]        I445ede2983c7470b4418a2ec0cbbd5e1;
wire [MAX_SUM_WDTH_L-1:0]        Iba61bc5c2e1230784d619375b7c756b4;
reg  [MAX_SUM_WDTH_L-1:0]        I034e56cd77ee400ed81b78177b202930;
wire [MAX_SUM_WDTH_L-1:0]        I613acad8a236e9deeb6967de9c067a48;
reg  [MAX_SUM_WDTH_L-1:0]        I08edadbd9366786f96b44268d096b4aa;
wire [MAX_SUM_WDTH_L-1:0]        I427eb014c821ba5108aaa6ebbd8bc23c;
reg  [MAX_SUM_WDTH_L-1:0]        I8f86a7af86eb04c5df18e09888cdce7b;
wire [MAX_SUM_WDTH_L-1:0]        I9b3fc0250b26e6faa2b7b44e863ff3f0;
reg  [MAX_SUM_WDTH_L-1:0]        Ic00d037a11f8a27ab34e4daab8c9c2e6;
wire [MAX_SUM_WDTH_L-1:0]        I79c12183f8bb94f4a3ce466570eadb80;
reg  [MAX_SUM_WDTH_L-1:0]        I4d95ceccc6c3ad37f13c98339c59e5c4;
wire [MAX_SUM_WDTH_L-1:0]        Id4ba2f12931de7439cd52eb15b0241eb;
reg  [MAX_SUM_WDTH_L-1:0]        I1ea967d377f462a0e06d7d0d4d95b342;
wire [MAX_SUM_WDTH_L-1:0]        I430558329b5398ffd51855414df8ba17;
reg  [MAX_SUM_WDTH_L-1:0]        Ib0feec63123e66bd6ad6935e9b7fa6bf;
wire [MAX_SUM_WDTH_L-1:0]        I4eacf5b6fddf6cb1dad592392eeef166;
reg  [MAX_SUM_WDTH_L-1:0]        I7d120060ddae9ff8f7206b3ef63eda50;
wire [MAX_SUM_WDTH_L-1:0]        I64921a58b87a14a3d6d02647f5c4a496;
reg  [MAX_SUM_WDTH_L-1:0]        Ib47f8f72386e2e65a88fbadd3a705225;
wire [MAX_SUM_WDTH_L-1:0]        I9a93abf3585f9f937118adfdacdd8736;
reg  [MAX_SUM_WDTH_L-1:0]        I4e0efc35346e2934f5bb4c34a4bc5f90;
wire [MAX_SUM_WDTH_L-1:0]        Ib368c9afabdccf356ff389540397e3e9;
reg  [MAX_SUM_WDTH_L-1:0]        I3ca1014802f58087e3434a1e0df19c01;
wire [MAX_SUM_WDTH_L-1:0]        I939d31990dc2265d78b3d5b9a031f0df;
reg  [MAX_SUM_WDTH_L-1:0]        I688a3879b7be1544e6f94b4221c03213;
wire [MAX_SUM_WDTH_L-1:0]        I3ded8a67a0163feb95cafacb2c539412;
reg  [MAX_SUM_WDTH_L-1:0]        Ic22988138610c8671ec342f65f34c7ae;
wire [MAX_SUM_WDTH_L-1:0]        I20c10afd04ed128ce31162ca3c1a89fa;
reg  [MAX_SUM_WDTH_L-1:0]        I0b85fdd83569e5cbb7d71eed50cb32fd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I71db9043fb2adee1e96818330469e51d;
reg  [MAX_SUM_WDTH_L-1:0]        Idf55390c11e5b41ebc2a28e0af109913;
wire [MAX_SUM_WDTH_L-1:0]        I64112bb2686f6348b7caaf3e0cf6a4aa;
reg  [MAX_SUM_WDTH_L-1:0]        I6b48935ea25672ee9a42f49eae9e519f;
wire [MAX_SUM_WDTH_L-1:0]        Ib4d8b49de697e1a70b07e76e836872b5;
reg  [MAX_SUM_WDTH_L-1:0]        I6a9e6c39c20e45773dab7823a7ff9486;
wire [MAX_SUM_WDTH_L-1:0]        I67dd716c2039d45a57fe94847cf2eef5;
reg  [MAX_SUM_WDTH_L-1:0]        I42907182010c5889ddb7a700ead16525;
wire [MAX_SUM_WDTH_L-1:0]        I60558c2a8261a6c4a06491a95c40dfec;
reg  [MAX_SUM_WDTH_L-1:0]        Ib6c26f3e3358cc2ed6fbda83eabd4bd3;
wire [MAX_SUM_WDTH_L-1:0]        I37e4ed1440968cf86567341f4febf6a7;
reg  [MAX_SUM_WDTH_L-1:0]        Ia50d85808790790450f87a5246874b3f;
wire [MAX_SUM_WDTH_L-1:0]        I369a541788e6ec2dbf5a29a93b8e9379;
reg  [MAX_SUM_WDTH_L-1:0]        Id4a1744702d7808a80bc40697c864765;
wire [MAX_SUM_WDTH_L-1:0]        I7fcf3847a6884d9e2cb216ac22cc6eea;
reg  [MAX_SUM_WDTH_L-1:0]        I0cf3d2f3e6793a2dcf15949da16ad28d;
wire [MAX_SUM_WDTH_L-1:0]        Ifc34e5240f1440c3a0415cc944241208;
reg  [MAX_SUM_WDTH_L-1:0]        I90bd9107f4c931fa1ccb92998ea8cdeb;
wire [MAX_SUM_WDTH_L-1:0]        I7e7a9c6ba8c0e7b945fc5cbc7def9c6b;
reg  [MAX_SUM_WDTH_L-1:0]        Ida1c729e6bfcec2c31a92aa9002f2c68;
wire [MAX_SUM_WDTH_L-1:0]        I8ea9c190206ea186295c33528d45551c;
reg  [MAX_SUM_WDTH_L-1:0]        Ib848feeccd0ea78ebc8ba8368534c3d1;
wire [MAX_SUM_WDTH_L-1:0]        I70f9d851136c9e8fb264fb43d6ebeb61;
reg  [MAX_SUM_WDTH_L-1:0]        Icc11970bbae3adcfa33a0e5dba3e78f4;
wire [MAX_SUM_WDTH_L-1:0]        Iea50b0ab0e00bfce47e6fdb129ea4cae;
reg  [MAX_SUM_WDTH_L-1:0]        I86bb4ef4bdd7af8861280ef30fbeeeea;
wire [MAX_SUM_WDTH_L-1:0]        Ie74b8877e9a7df32f3f5674aab1300af;
reg  [MAX_SUM_WDTH_L-1:0]        I7e0c259c6c7bacdff5edc44a22e005ba;
wire [MAX_SUM_WDTH_L-1:0]        Iaa3d8acf714f23e5059aa21cc1c36dd4;
reg  [MAX_SUM_WDTH_L-1:0]        I897ddba059b27f7ed009b0cb70cfb46f;
wire [MAX_SUM_WDTH_L-1:0]        Ic98698807ac6942eaa491de5a2a523c0;
reg  [MAX_SUM_WDTH_L-1:0]        I4496243eb0542a514b551b4d09bffd7d;
wire [MAX_SUM_WDTH_L-1:0]        I3579622172c0ccdf3eeb3bd490b2e6db;
reg  [MAX_SUM_WDTH_L-1:0]        Ic931fb08b2e8441321ebdeed84576a0d;
wire [MAX_SUM_WDTH_L-1:0]        I1369d79bd170cc9b7ed0352e0701261b;
reg  [MAX_SUM_WDTH_L-1:0]        Ieb6af5390b98e893ee05a939c16d2ffd;
wire [MAX_SUM_WDTH_L-1:0]        I16196f7cfe21843797e1f3ef19b09048;
reg  [MAX_SUM_WDTH_L-1:0]        Ic2a54bad4c5a8885dd24b8687c6db0de;
wire [MAX_SUM_WDTH_L-1:0]        I20e403ad09d5eeb59020f7fe3b683432;
reg  [MAX_SUM_WDTH_L-1:0]        I6ecbad763d2b48b78a0584beaefc78ee;
wire [MAX_SUM_WDTH_L-1:0]        I8d6ef29e41c3ef0fe66820e77c486591;
reg  [MAX_SUM_WDTH_L-1:0]        I20556d23c873c71c7ebc8a961bf40251;
wire [MAX_SUM_WDTH_L-1:0]        I77fcee77b0cb1c65ca313526461231e4;
reg  [MAX_SUM_WDTH_L-1:0]        I79012e6351e6320c22437aa216ea4df1;
wire [MAX_SUM_WDTH_L-1:0]        I40c64a3c54b15800ed725dfce5144f17;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf74ab9af877d27c3a6f3881f00ddaf1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I57bddc5d3b9daf16fa9c2eaa3a148a03;
reg  [MAX_SUM_WDTH_L-1:0]        I843d35db35d7b42a87ce78d3772cec2f;
wire [MAX_SUM_WDTH_L-1:0]        I5d3dc544f4e02f31e8dbc2b399afa89e;
reg  [MAX_SUM_WDTH_L-1:0]        I2b1398b4bfd374d7221b0a68da28e979;
wire [MAX_SUM_WDTH_L-1:0]        I0bc53eebdddc25c9c1423068bbe7a2a1;
reg  [MAX_SUM_WDTH_L-1:0]        I6f615d6e74b0c02f8e4265523ad16404;
wire [MAX_SUM_WDTH_L-1:0]        I23429a89ac40e62e5b13ec75e348e432;
reg  [MAX_SUM_WDTH_L-1:0]        Iae8a98dd4a7cbfbc56c1404b6a2020af;
wire [MAX_SUM_WDTH_L-1:0]        I417ae67e3ed05fb6ac8b24bcba692a83;
reg  [MAX_SUM_WDTH_L-1:0]        Iad53375a54d01c559c74981bf279dfb5;
wire [MAX_SUM_WDTH_L-1:0]        I5edf732eb5451f0f84087b8ccccab387;
reg  [MAX_SUM_WDTH_L-1:0]        I5db1307f922e0c742d7d9f3a79a4a4f3;
wire [MAX_SUM_WDTH_L-1:0]        I26833c93cc1b8be86febb45560ae4707;
reg  [MAX_SUM_WDTH_L-1:0]        I9f78172ed5bf73752196f9a8810005f3;
wire [MAX_SUM_WDTH_L-1:0]        Iab7fe9d9176e8ceb00b7d04116dc0236;
reg  [MAX_SUM_WDTH_L-1:0]        If85a22d670d47f491dd7568d0453ba1d;
wire [MAX_SUM_WDTH_L-1:0]        Ie66e4f53df7e0bb44442a3c74883ab30;
reg  [MAX_SUM_WDTH_L-1:0]        Ib9e529170b2896e930a839295796fd31;
wire [MAX_SUM_WDTH_L-1:0]        I591dd226d239200c681a1aac16849d31;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7af536846bac40c1f221d1f72c6c25c;
wire [MAX_SUM_WDTH_L-1:0]        Ic572d19feb1b9d45cb81aa0aeee01340;
reg  [MAX_SUM_WDTH_L-1:0]        Ib0eb61a2cb831dd35ce9850994e7c2da;
wire [MAX_SUM_WDTH_L-1:0]        I31306ed55c012f4e3f3da72bc404d6ba;
reg  [MAX_SUM_WDTH_L-1:0]        I89d338f59960af7a47595d6afa206abc;
wire [MAX_SUM_WDTH_L-1:0]        I374c888e91b747a2a6b58649c4a1969b;
reg  [MAX_SUM_WDTH_L-1:0]        Ib3c1176eb8991e3e85855a9fe845c303;
wire [MAX_SUM_WDTH_L-1:0]        Ic71fea427a788b416d088a44f2600c51;
reg  [MAX_SUM_WDTH_L-1:0]        I93073d05d509b821a743998cf32c58ee;
wire [MAX_SUM_WDTH_L-1:0]        Ib6fec22f8466773bb13224a90a4e3c2d;
reg  [MAX_SUM_WDTH_L-1:0]        Iab6dac1909c1564c3890ffecc13418df;
wire [MAX_SUM_WDTH_L-1:0]        Id30dc8c00fd07e9ad68a8fc3c740557f;
reg  [MAX_SUM_WDTH_L-1:0]        I1b75eeb29167a171d89f6e67039436d5;
wire [MAX_SUM_WDTH_L-1:0]        I85777d4d61b8e6fc99706bbe7fbfad8c;
reg  [MAX_SUM_WDTH_L-1:0]        I3a31adc52a1405555017b2ddf219b407;
wire [MAX_SUM_WDTH_L-1:0]        I707e0745e78aef8c802c0fd5a7b58ae5;
reg  [MAX_SUM_WDTH_L-1:0]        Iaadba89c6a370240fc0758029f7d8db0;
wire [MAX_SUM_WDTH_L-1:0]        I513c23daa981e69789b074975a589954;
reg  [MAX_SUM_WDTH_L-1:0]        I4f4a64fb3ced7d9f7ee4513178e9655a;
wire [MAX_SUM_WDTH_L-1:0]        I3b0ea0ad1bf5f5820e582b0c1f97d949;
reg  [MAX_SUM_WDTH_L-1:0]        I0c76ca58f69c91758e755cd581241284;
wire [MAX_SUM_WDTH_L-1:0]        I857759675a04284a230c6e09e993db26;
reg  [MAX_SUM_WDTH_L-1:0]        I2312bce18958346149c868846e04643b;
wire [MAX_SUM_WDTH_L-1:0]        I943326eaa918c39cb3fe412c77d8b131;
reg  [MAX_SUM_WDTH_L-1:0]        I3e154098cb0a48f1c23234f46613f406;
wire [MAX_SUM_WDTH_L-1:0]        I9dcf55a3343d214ab70cbde50a34da4d;
reg  [MAX_SUM_WDTH_L-1:0]        I1645c1c588bcbf15dd62d47e08b8e139;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I1fe6a30dcbcbdcfc0b3d6bbe38e9c3bc;
reg  [MAX_SUM_WDTH_L-1:0]        I4c25de66590e1745d37112e08d8c8e2c;
wire [MAX_SUM_WDTH_L-1:0]        I39216b818931b9d2fb6a93e5eda743aa;
reg  [MAX_SUM_WDTH_L-1:0]        Ia03092ac621b8dd1c206fea1e8b0215f;
wire [MAX_SUM_WDTH_L-1:0]        I24238e5bba0bf63288ad44c5dd3545f3;
reg  [MAX_SUM_WDTH_L-1:0]        I5c9bdb033436dc9f6069baca31f24c2d;
wire [MAX_SUM_WDTH_L-1:0]        Ic0a34c6b56cc30ddec7e5b755e18a27d;
reg  [MAX_SUM_WDTH_L-1:0]        I8f07cf4865480f18ad6945974ec2231c;
wire [MAX_SUM_WDTH_L-1:0]        I45e63318c784a30395ca1bbc692d1402;
reg  [MAX_SUM_WDTH_L-1:0]        I4a7119e8862fe4a6a4100dd9ac67dd24;
wire [MAX_SUM_WDTH_L-1:0]        Iae0e9a6d88b4fba34944cd2f0dd5c9ed;
reg  [MAX_SUM_WDTH_L-1:0]        Id78fcfc6724a05f46d44d7c3e7d0c756;
wire [MAX_SUM_WDTH_L-1:0]        I91d8bc9088850978c17bfa5f0bf93b26;
reg  [MAX_SUM_WDTH_L-1:0]        I7cbd9d619623cbabf8ed6b1fece8f012;
wire [MAX_SUM_WDTH_L-1:0]        I014cecda30cbc4e25a1265a65ed0f0d4;
reg  [MAX_SUM_WDTH_L-1:0]        I58951165d251e370b0f3b3fb537aed18;
wire [MAX_SUM_WDTH_L-1:0]        I845250d1ee6395d022a0a20698eea330;
reg  [MAX_SUM_WDTH_L-1:0]        I21daac106f526d84cb8fa5239c19499d;
wire [MAX_SUM_WDTH_L-1:0]        I5d36a24496d96371aba3f0407c21e34d;
reg  [MAX_SUM_WDTH_L-1:0]        I178029cec3a5d6141abdfa91b91fdbf4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If2f7a871f45dc098b3ebe056153235c7;
reg  [MAX_SUM_WDTH_L-1:0]        I96dfb2efbb55a644616e3474ed07c364;
wire [MAX_SUM_WDTH_L-1:0]        Ib49df5d97f0ba140b6ec5f80aae719d6;
reg  [MAX_SUM_WDTH_L-1:0]        I7a17d8f0e2d16c441044db68ee037731;
wire [MAX_SUM_WDTH_L-1:0]        Ib25900518732253ccc4800716f3d772d;
reg  [MAX_SUM_WDTH_L-1:0]        I2ced9bb3ae6bdc5b5ef2865fb46abf07;
wire [MAX_SUM_WDTH_L-1:0]        I9d9b410818773fca2bc21ed678683369;
reg  [MAX_SUM_WDTH_L-1:0]        I89a93384020d93cf4d26b3902e06cd9e;
wire [MAX_SUM_WDTH_L-1:0]        Ia003b700205a0b2faf1cefa2c85c4df0;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbb47d29b9a45559c13ffa3b046c66f5;
wire [MAX_SUM_WDTH_L-1:0]        I3b98b4efc159ac3eb3c7ea322459b666;
reg  [MAX_SUM_WDTH_L-1:0]        I0034177eb1049577a3578b371527f34b;
wire [MAX_SUM_WDTH_L-1:0]        Ibfe30b79869ff3125c248f623c494d09;
reg  [MAX_SUM_WDTH_L-1:0]        I22d9ea7bb5a1a3405bcd04b9af40fa62;
wire [MAX_SUM_WDTH_L-1:0]        Ice88c3ab21612bbd46676c650d9f4dbc;
reg  [MAX_SUM_WDTH_L-1:0]        I8a632e7a911bf5726fee587189cb6f16;
wire [MAX_SUM_WDTH_L-1:0]        Ideadf767ef2ab66a1495ead1806ffe47;
reg  [MAX_SUM_WDTH_L-1:0]        I3765afc490b34e8a310998a4ebcff8cb;
wire [MAX_SUM_WDTH_L-1:0]        I28749b0f4f83f99b9082f7004e72aa70;
reg  [MAX_SUM_WDTH_L-1:0]        I7607e800ae46a96e016b303120da4247;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I71ef3d84207d8995c13e88c16a0bacf8;
reg  [MAX_SUM_WDTH_L-1:0]        I29b2f1fddee5e32f217d25410bcfce4f;
wire [MAX_SUM_WDTH_L-1:0]        I630979d7924b3c17fe0aeaa04507ed03;
reg  [MAX_SUM_WDTH_L-1:0]        Iba5f8a31a81f6aa06f5e38c03dc6db54;
wire [MAX_SUM_WDTH_L-1:0]        I50a84fa93d73bfe0287f3297707b1901;
reg  [MAX_SUM_WDTH_L-1:0]        Ifcb5c907ad503331317599e4e0ce7be8;
wire [MAX_SUM_WDTH_L-1:0]        I19d6383f6319e9ed4b4f16fdf7a40cef;
reg  [MAX_SUM_WDTH_L-1:0]        I62d6f2ab4ec8b6ecfa544ad4d90eb30b;
wire [MAX_SUM_WDTH_L-1:0]        I3515fa4f304e4b1537c612ca0212b4bc;
reg  [MAX_SUM_WDTH_L-1:0]        Ide65414c51b3cb182c0f2f238903d60a;
wire [MAX_SUM_WDTH_L-1:0]        Ia154b83a5a01bf0ea74fcc873e45d980;
reg  [MAX_SUM_WDTH_L-1:0]        I03a8dc2288eaeb619e746990e20cc868;
wire [MAX_SUM_WDTH_L-1:0]        If021572d95ea7fcbae1454447dbbe212;
reg  [MAX_SUM_WDTH_L-1:0]        Id81c1b44d16ddbcd466382c60fe84986;
wire [MAX_SUM_WDTH_L-1:0]        Ib6c860f3146839d2c0e925007ac02d67;
reg  [MAX_SUM_WDTH_L-1:0]        I503d72f4a2fd20dbf35aa27321d2ede7;
wire [MAX_SUM_WDTH_L-1:0]        I21ae48e98044dcc69386800f72cc5fb7;
reg  [MAX_SUM_WDTH_L-1:0]        Id6595a4cf33062d1f05cbcee2d0685f1;
wire [MAX_SUM_WDTH_L-1:0]        I4f436764c02c61027d89854865770734;
reg  [MAX_SUM_WDTH_L-1:0]        I83ebdd7331ca8fbcf5250851b346c0b0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If213a0715834eb56c9c8862dcd643f36;
reg  [MAX_SUM_WDTH_L-1:0]        I7f6ea26cdfe5986065e7b5aa6842cc1c;
wire [MAX_SUM_WDTH_L-1:0]        If1eced44ede97a4e0ec55c26df8d6935;
reg  [MAX_SUM_WDTH_L-1:0]        Idab1ec32c20f93c4cc1acb38158f92d5;
wire [MAX_SUM_WDTH_L-1:0]        Ibe579be01c1b2925be397ab7d202c200;
reg  [MAX_SUM_WDTH_L-1:0]        I0738add83419502e73674ded2f1ad6c7;
wire [MAX_SUM_WDTH_L-1:0]        I675731b8fceb36c9a103803dea3700bc;
reg  [MAX_SUM_WDTH_L-1:0]        I6c93e63a8e5a2dbd598f1565c7323b39;
wire [MAX_SUM_WDTH_L-1:0]        I01374171f18d419d149433d7c789f1ef;
reg  [MAX_SUM_WDTH_L-1:0]        I4aa57a9d46371f1680d5f95596f60b5d;
wire [MAX_SUM_WDTH_L-1:0]        I9f66291cd8f80896cf27fa0b8382f465;
reg  [MAX_SUM_WDTH_L-1:0]        I5369a7203b78951a3c006c2d3b22507c;
wire [MAX_SUM_WDTH_L-1:0]        I73341b7d2d30f5fe7ce2d8659331de3b;
reg  [MAX_SUM_WDTH_L-1:0]        Ie72a79a6966cf198687b7c8a8bcdeb13;
wire [MAX_SUM_WDTH_L-1:0]        Ieb9c6cc947f6e0429770118119be79e1;
reg  [MAX_SUM_WDTH_L-1:0]        Ie917ae4c44ab0f9c2f1747ff0d2a754e;
wire [MAX_SUM_WDTH_L-1:0]        I2c58e39ab3b79963fa0eddc7180070dc;
reg  [MAX_SUM_WDTH_L-1:0]        I0b1a31ccb34a742552c11b1945e23dd8;
wire [MAX_SUM_WDTH_L-1:0]        I789b342281d9ed8dbc03af5c0c508062;
reg  [MAX_SUM_WDTH_L-1:0]        I9a65a845cf2eced39050e8481665f557;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I95b62a2fcb0af75048d095dde733ddbc;
reg  [MAX_SUM_WDTH_L-1:0]        I3b402b35d38a9fde312c89b82297c1a5;
wire [MAX_SUM_WDTH_L-1:0]        I1e9d61b53dd7ce47230b341cc1b4e8b4;
reg  [MAX_SUM_WDTH_L-1:0]        I309fa33562370e339c19e2377e6a6a7a;
wire [MAX_SUM_WDTH_L-1:0]        If5d6db7c002ad813677ca165380839b0;
reg  [MAX_SUM_WDTH_L-1:0]        I7d06aed81222a030837cad2074c68e19;
wire [MAX_SUM_WDTH_L-1:0]        I0f7ceff0b6160697dbd097293de15156;
reg  [MAX_SUM_WDTH_L-1:0]        I835cc6af0cd8189035f2441c2e0d3100;
wire [MAX_SUM_WDTH_L-1:0]        I2e142efe8de226e1a283576d1ae9ced9;
reg  [MAX_SUM_WDTH_L-1:0]        If6f768d12f04087246a0d65de1aef99b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I88e4b172c1b5c2733bf050fa442964ce;
reg  [MAX_SUM_WDTH_L-1:0]        Ie4b180e1e2cadb865b0eaf6509f99dbb;
wire [MAX_SUM_WDTH_L-1:0]        Ie1f997dc210ff90c7ff78737d1240c30;
reg  [MAX_SUM_WDTH_L-1:0]        Ie329a11fc3f6f59f6f1790612fde3250;
wire [MAX_SUM_WDTH_L-1:0]        I31307a02f9909905fd672eeaf54422a6;
reg  [MAX_SUM_WDTH_L-1:0]        Idb7ddbee4076f7bf49177e69f5e4d112;
wire [MAX_SUM_WDTH_L-1:0]        I1e2dbb3cd67d96f046b39fd52947ff4e;
reg  [MAX_SUM_WDTH_L-1:0]        I614d66a7dca2d08efdfdc157ca803d5c;
wire [MAX_SUM_WDTH_L-1:0]        Icad3b8650e3c4b3a425e1a1c7da14c1a;
reg  [MAX_SUM_WDTH_L-1:0]        Iea16eb0ab70ebb1bc47ae55e11ced62d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I40acfb6473e56562b5bc1e7bfdeed8a6;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa8db43284d5bbebaed4f72d65cf9f92;
wire [MAX_SUM_WDTH_L-1:0]        I06a6d7c6a5be68cb75d83b2d8a1d3217;
reg  [MAX_SUM_WDTH_L-1:0]        I365d9f3e8b2a9890427f07386deeb093;
wire [MAX_SUM_WDTH_L-1:0]        I3d3ebea1cf84cec93ff60459177fdd18;
reg  [MAX_SUM_WDTH_L-1:0]        I466aaa0b6cde2ade1901797b8c11e32c;
wire [MAX_SUM_WDTH_L-1:0]        I59868ed1411b6439564cc73edf55297d;
reg  [MAX_SUM_WDTH_L-1:0]        I7057e329a65ab240ed6cfa824307af65;
wire [MAX_SUM_WDTH_L-1:0]        I97ae3d6c75edf1fd87347a8fd50fd27d;
reg  [MAX_SUM_WDTH_L-1:0]        I624e50e3457d33d12680eaf8e7c34aa3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If98ad7df6cb49466733052834b458bb1;
reg  [MAX_SUM_WDTH_L-1:0]        I9f356fd6820c33fdb5baff05a781e192;
wire [MAX_SUM_WDTH_L-1:0]        I2ea63dcc06519b46da5b70cf36b68c76;
reg  [MAX_SUM_WDTH_L-1:0]        I39b9c7c664fe7017731877d145d55b44;
wire [MAX_SUM_WDTH_L-1:0]        I979c3adad47ed2b8488aa7beaab7a565;
reg  [MAX_SUM_WDTH_L-1:0]        Ic62ffbb9e58e0d08b0dec24bba1dc6f2;
wire [MAX_SUM_WDTH_L-1:0]        Idc93f47a3946c69fc0c956ec3e4d4c28;
reg  [MAX_SUM_WDTH_L-1:0]        I8da2a532288fb817e7dc0cb7b4e3761c;
wire [MAX_SUM_WDTH_L-1:0]        I3d57c80540bbdb043ce47c688950fd18;
reg  [MAX_SUM_WDTH_L-1:0]        I6a6e559f5c98f846014e8107fea5a5d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Id2083cbcf2aaa813c72071314c13ae6f;
reg  [MAX_SUM_WDTH_L-1:0]        Ibef9219f577b1a62dfdd77296fbfb24d;
wire [MAX_SUM_WDTH_L-1:0]        Iea95f61532bffc857f39331b244188d0;
reg  [MAX_SUM_WDTH_L-1:0]        I52e6688b5bfff75529d18e20b22832ce;
wire [MAX_SUM_WDTH_L-1:0]        I42dd514d52d448707c7dcc5c799ee7f1;
reg  [MAX_SUM_WDTH_L-1:0]        Iff22c49354eefca0ea3c5959c14b782c;
wire [MAX_SUM_WDTH_L-1:0]        Ib6ee76ae9fed974530f73fb401405e27;
reg  [MAX_SUM_WDTH_L-1:0]        Ie5377bbdb4111ed00356d5b7737102f3;
wire [MAX_SUM_WDTH_L-1:0]        I3aea3d7d9965e4cde24ba83120af804e;
reg  [MAX_SUM_WDTH_L-1:0]        I55bf0f3379a8c44634b8f0a3d06c049e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3b1550f5b3e421d44005a01b0075bf33;
reg  [MAX_SUM_WDTH_L-1:0]        I9bc9541607f4f6aedb686cdde297bcda;
wire [MAX_SUM_WDTH_L-1:0]        I00bc9cf3ab66e198dd7bf2cc930aa2c5;
reg  [MAX_SUM_WDTH_L-1:0]        Ia4620554fbb1d81a71a15a846e4be2f5;
wire [MAX_SUM_WDTH_L-1:0]        I79d4eac1731095e588b7003d1c83aba7;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb31b35388ba8ba2ecf98449308ee67d;
wire [MAX_SUM_WDTH_L-1:0]        I6512194d646b949c1f8037e3911a8720;
reg  [MAX_SUM_WDTH_L-1:0]        Ia20410fb3d56587f89a54c00b943b305;
wire [MAX_SUM_WDTH_L-1:0]        Ief2dcb1d14d5065729e66207068d0519;
reg  [MAX_SUM_WDTH_L-1:0]        I9d268f3da12e35b9a4229b7340c0f018;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib343818dd2f04189d56a6fc40c8da197;
reg  [MAX_SUM_WDTH_L-1:0]        I2fce29bd666082eedb2fb3ec8b5ae4dd;
wire [MAX_SUM_WDTH_L-1:0]        Ie38501f8b5cd9e64ed80bed953adbb48;
reg  [MAX_SUM_WDTH_L-1:0]        Ia1e8b61e2579a90f5c88ded11c7322c2;
wire [MAX_SUM_WDTH_L-1:0]        Id50a8c0b1739857f19228131b51f7937;
reg  [MAX_SUM_WDTH_L-1:0]        I8cf3718ba65b7fed72e3955f190e34d1;
wire [MAX_SUM_WDTH_L-1:0]        I8946d670fb58546b8854b34dad0e8430;
reg  [MAX_SUM_WDTH_L-1:0]        I7e802d300af54d394b4ee041798c0513;
wire [MAX_SUM_WDTH_L-1:0]        I122129edde3336f22ba613499bfabfc0;
reg  [MAX_SUM_WDTH_L-1:0]        Id4fd5a4b97cfa1e176a26f3a823c5516;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I2ce23daae62346911511cfea5bed788f;
reg  [MAX_SUM_WDTH_L-1:0]        Icbf8d4e75fc66c05eb49c5075696fb07;
wire [MAX_SUM_WDTH_L-1:0]        I5496ff29bde6957c01c5d7e5f2d8cbac;
reg  [MAX_SUM_WDTH_L-1:0]        I746a7e90adb2f213b75ae12a161aca0d;
wire [MAX_SUM_WDTH_L-1:0]        I66fe45afee3cd240ed3ef77262387f40;
reg  [MAX_SUM_WDTH_L-1:0]        Icb1029aaaaed8c698862ea9c5e22132c;
wire [MAX_SUM_WDTH_L-1:0]        Id08a0b67ee6d6e08628238b1e5ac0dc8;
reg  [MAX_SUM_WDTH_L-1:0]        Ib93ea7028c172373b53cdafecae32a67;
wire [MAX_SUM_WDTH_L-1:0]        I2b94a5c3e2ee6f13fae5ec588be73ba0;
reg  [MAX_SUM_WDTH_L-1:0]        If9628275b000e418f3903daebfdace92;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8b6ce93d2c7b309d4d043e938ef6cb12;
reg  [MAX_SUM_WDTH_L-1:0]        I830202fb6f08f98c7f71893a881bd555;
wire [MAX_SUM_WDTH_L-1:0]        I46d88449ca1db5f462e0442932bc5f53;
reg  [MAX_SUM_WDTH_L-1:0]        I6f38bc9359562f57c1603355e9ee312b;
wire [MAX_SUM_WDTH_L-1:0]        I402417fdf22d1b9e08e905e3206a6edc;
reg  [MAX_SUM_WDTH_L-1:0]        I4701b732d59c26e3790a63c1936f9a24;
wire [MAX_SUM_WDTH_L-1:0]        I287e3042873300b74530542044f57277;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5d28d8f73d17ab6df6a1291e50c04ab;
wire [MAX_SUM_WDTH_L-1:0]        I4c6118afff7012ebdec7b6168f1ba067;
reg  [MAX_SUM_WDTH_L-1:0]        I81259f391db792339824ad5dd1a0057b;
wire [MAX_SUM_WDTH_L-1:0]        I444e2151e66af9ec6c1e984ad706b7a0;
reg  [MAX_SUM_WDTH_L-1:0]        I6f09ac63effe67a86798b9b4e1690664;
wire [MAX_SUM_WDTH_L-1:0]        I3c800d94a189c70fb956298deb686700;
reg  [MAX_SUM_WDTH_L-1:0]        I370b4b3a0048a93ba374a40e170c75a3;
wire [MAX_SUM_WDTH_L-1:0]        I0b3393ffccd4b2a9b42a68f185b074f8;
reg  [MAX_SUM_WDTH_L-1:0]        I3f8476d0aa0ea2439b67ea1a4adf36c5;
wire [MAX_SUM_WDTH_L-1:0]        Ie1996578a600cbb605703974fcd3494a;
reg  [MAX_SUM_WDTH_L-1:0]        I35b52dba10a8a5b22b518388fecac82d;
wire [MAX_SUM_WDTH_L-1:0]        Ib912bf53b3fc6753b228a488d9d25520;
reg  [MAX_SUM_WDTH_L-1:0]        Ic7db274ed18e6fdecf30381a31238777;
wire [MAX_SUM_WDTH_L-1:0]        I77f81eeb736f7ad4abcd88fa9b952bc0;
reg  [MAX_SUM_WDTH_L-1:0]        I2c4e538a8db759e9799541d9178ec61e;
wire [MAX_SUM_WDTH_L-1:0]        Ic09db56c2b021b09e0cf4fe501f2a5ec;
reg  [MAX_SUM_WDTH_L-1:0]        Ief6d4c3f5ef8663e111ef99347b023f5;
wire [MAX_SUM_WDTH_L-1:0]        I576cf92938eb1c168e0f9ee1b6bf0be7;
reg  [MAX_SUM_WDTH_L-1:0]        Id95e964e5faecb52c72669b0d28a4bf5;
wire [MAX_SUM_WDTH_L-1:0]        Ia1d7ca394ee29ff9cc463c525fbf7947;
reg  [MAX_SUM_WDTH_L-1:0]        I0fcef4538102ac6d24aa7090d5405afa;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I7fff588b55c99166b13cd816d6a5c166;
reg  [MAX_SUM_WDTH_L-1:0]        I055019e38eec6badd1739033d43d7d97;
wire [MAX_SUM_WDTH_L-1:0]        I755d06b657ce02dabc6dbb6d44e619e6;
reg  [MAX_SUM_WDTH_L-1:0]        I35c20a6e823da77a870b421eef2e0a95;
wire [MAX_SUM_WDTH_L-1:0]        If86871aa91ead2d985e915f4d58408f3;
reg  [MAX_SUM_WDTH_L-1:0]        I32cc12cdacef1a4ef64577e0fa977f46;
wire [MAX_SUM_WDTH_L-1:0]        Ie53d1075a122b58f8ee4282b91322ccc;
reg  [MAX_SUM_WDTH_L-1:0]        I26b3f2360ca4a8caee61b2f3a3a08267;
wire [MAX_SUM_WDTH_L-1:0]        I54acee9cb56584f9876867492fabe469;
reg  [MAX_SUM_WDTH_L-1:0]        I5ef9b7dc0c63e9ca6a5fb5f7ffa06041;
wire [MAX_SUM_WDTH_L-1:0]        Ia4e992a0d0c4f89e3bbaba81b6be3c41;
reg  [MAX_SUM_WDTH_L-1:0]        If881473b05090f40a027d7eeee7f7ed9;
wire [MAX_SUM_WDTH_L-1:0]        I8c215a65ea37a535fc9230a0141d209f;
reg  [MAX_SUM_WDTH_L-1:0]        I23bd59ab5b038935301396aaf2acefc1;
wire [MAX_SUM_WDTH_L-1:0]        I564374188b8065f6a46972355d27b0a9;
reg  [MAX_SUM_WDTH_L-1:0]        I874386d94dacf84e699d159af1a49836;
wire [MAX_SUM_WDTH_L-1:0]        Ide9ea9ced1a2398876700b19dd25a080;
reg  [MAX_SUM_WDTH_L-1:0]        I95bfe51a759bf4165168e5e3b99d6b34;
wire [MAX_SUM_WDTH_L-1:0]        I999b0d3276b81801b5a6a5af4d98e6fc;
reg  [MAX_SUM_WDTH_L-1:0]        I4ba5b2f9b7ec0937ecd2c9945cf6de87;
wire [MAX_SUM_WDTH_L-1:0]        I94b6767c45b74142ab2d457b5fe3b64e;
reg  [MAX_SUM_WDTH_L-1:0]        I0b08fb8db0e8a1de3d416907c87fe700;
wire [MAX_SUM_WDTH_L-1:0]        I2062510b4d8249d8a9b75377d4513266;
reg  [MAX_SUM_WDTH_L-1:0]        Ie030d12e5acf9ef4975a17c83b2481c1;
wire [MAX_SUM_WDTH_L-1:0]        Iba97ce79b40d24270208680c74b41799;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7a0e852d3dfcef950804ea0ebb0c80a;
wire [MAX_SUM_WDTH_L-1:0]        I35b405f29c891a3ccaf0b64443d114e9;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa4c38d030eab2b7899399aa0d7886d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib44c2f3a3916b3eaa7452f0126f934ab;
reg  [MAX_SUM_WDTH_L-1:0]        Icce7ff1d652d4d9c2be5ecf679059bbe;
wire [MAX_SUM_WDTH_L-1:0]        I2f0d79178e118fb89f9504e5f75fd612;
reg  [MAX_SUM_WDTH_L-1:0]        If816bc5eacaea23443602e575ddf60b8;
wire [MAX_SUM_WDTH_L-1:0]        I1e5f655fd8601930d7c9307aab545391;
reg  [MAX_SUM_WDTH_L-1:0]        I3b224a4ded05446cc5300d430bdd1947;
wire [MAX_SUM_WDTH_L-1:0]        I77691bc302dff581968daeeeaf44e9a9;
reg  [MAX_SUM_WDTH_L-1:0]        Ia5fc5cfb0e52237b407b37a3858fccb5;
wire [MAX_SUM_WDTH_L-1:0]        Ic0f0982cdd813ef3da99d8534e23c9e7;
reg  [MAX_SUM_WDTH_L-1:0]        I92f8ba6e7f8e9b30fb5b6973eb8fd03e;
wire [MAX_SUM_WDTH_L-1:0]        I449f136e29d92eedd2273b58bd34431c;
reg  [MAX_SUM_WDTH_L-1:0]        Icdfa60d2a024dd934f7e6639c6cb2c28;
wire [MAX_SUM_WDTH_L-1:0]        I0906f557008adaf488966d5aa989e6ae;
reg  [MAX_SUM_WDTH_L-1:0]        Ifff70b976513eaa42b6bd4b80c98611e;
wire [MAX_SUM_WDTH_L-1:0]        Ic0b69b2b6f55b4613bac3aad8e864c9f;
reg  [MAX_SUM_WDTH_L-1:0]        Ica12fa8b631b70a6bbe9f6e92bf73ea0;
wire [MAX_SUM_WDTH_L-1:0]        I6ccadd50ca8d59878cf089a35319b6c0;
reg  [MAX_SUM_WDTH_L-1:0]        Ie69c255335760f706c644b115887269b;
wire [MAX_SUM_WDTH_L-1:0]        Ia5aabf0fe6a5d3731b363c80a7238a14;
reg  [MAX_SUM_WDTH_L-1:0]        Idb06676b41de19bc86eae34c292183d9;
wire [MAX_SUM_WDTH_L-1:0]        I217dc03c6c19195b3c2f478b2b8b0bb8;
reg  [MAX_SUM_WDTH_L-1:0]        Ib21d2306d5ded3406fac754e69a10d20;
wire [MAX_SUM_WDTH_L-1:0]        I70c592140d0fd63e2b9b8ab9b619df9a;
reg  [MAX_SUM_WDTH_L-1:0]        Ib41d1aa2dcf81879976fb8964cbf6f79;
wire [MAX_SUM_WDTH_L-1:0]        I4d9ac478c0c0b7191a0ffeb3c6d7c521;
reg  [MAX_SUM_WDTH_L-1:0]        I5f8f5e246f008b8d8c75f72828337bab;
wire [MAX_SUM_WDTH_L-1:0]        I8bb214c6ec5a16858101699241a1b4bb;
reg  [MAX_SUM_WDTH_L-1:0]        Id6625e78da0e14d2eeb19cc8ac6520e0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iff81d398838ac6181e09d95903bf57a9;
reg  [MAX_SUM_WDTH_L-1:0]        I6d9ddc6afa559ac35c042df1a9390ce9;
wire [MAX_SUM_WDTH_L-1:0]        I710eb104c64c7eb72a55cbfc11bff827;
reg  [MAX_SUM_WDTH_L-1:0]        I9334055c7833676469670372d3c5cc31;
wire [MAX_SUM_WDTH_L-1:0]        I9f2d9117540a1d6902b1a7ec3e9d5ab4;
reg  [MAX_SUM_WDTH_L-1:0]        I0c97d772c737c6ff85b584bf69ccaf93;
wire [MAX_SUM_WDTH_L-1:0]        Ie3204e2e502d2c192994f3c74f1ea38f;
reg  [MAX_SUM_WDTH_L-1:0]        Ic6ce97ae85d91dd8a79f3f9d0da375a2;
wire [MAX_SUM_WDTH_L-1:0]        I97f03a2baec02107032233e68c0b146b;
reg  [MAX_SUM_WDTH_L-1:0]        I83ff9a2750b298b0f7c9b6ce13f574af;
wire [MAX_SUM_WDTH_L-1:0]        I860ccc9f56a3376ea0e8137a045fe650;
reg  [MAX_SUM_WDTH_L-1:0]        I85699a2a05c343a6a9e828af6d445e9e;
wire [MAX_SUM_WDTH_L-1:0]        I7b00537ae91be6f2ad8be0776e29da79;
reg  [MAX_SUM_WDTH_L-1:0]        I51f6e39b24b2554884e381be79f47ff2;
wire [MAX_SUM_WDTH_L-1:0]        I68413adceb35fe859824c32bb76d9906;
reg  [MAX_SUM_WDTH_L-1:0]        I9f65fd05c6929300860c8cbbde5607f2;
wire [MAX_SUM_WDTH_L-1:0]        Ib61183063f591e5845ca8ce70f598c79;
reg  [MAX_SUM_WDTH_L-1:0]        If09761d8f06051d4287ee29ac9c9fa19;
wire [MAX_SUM_WDTH_L-1:0]        Ia7a97e75655c4eaa8652f43c27d5ae50;
reg  [MAX_SUM_WDTH_L-1:0]        I33bfbe0bcca6d32c86b9576577e3f265;
wire [MAX_SUM_WDTH_L-1:0]        I0402af748fe9d48a514d23691a2cb6b8;
reg  [MAX_SUM_WDTH_L-1:0]        If2921210b1c05ecbf00af3a2bcb96ef4;
wire [MAX_SUM_WDTH_L-1:0]        I5e9d62da7f6aeaa717f5a394e2531210;
reg  [MAX_SUM_WDTH_L-1:0]        Ib074e38e280474a782da831a3e0028b4;
wire [MAX_SUM_WDTH_L-1:0]        Idb3666a01522d57729513cd3f18c9798;
reg  [MAX_SUM_WDTH_L-1:0]        I507449dde0bc0c8f53a10759436ec731;
wire [MAX_SUM_WDTH_L-1:0]        Ifb6e917336ab665d9bfea6dcfe21bc8c;
reg  [MAX_SUM_WDTH_L-1:0]        Id55a3e3f2d75baeba71a345fad695c69;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0adf84fd4ea2e882b59a42dad6683707;
reg  [MAX_SUM_WDTH_L-1:0]        I20984f43d22671639a7a178ad15aec04;
wire [MAX_SUM_WDTH_L-1:0]        I1d0e0cb3903cece98c3a65f920e5ab21;
reg  [MAX_SUM_WDTH_L-1:0]        I59f88336d6bdd50ded87d353fb5ce3e9;
wire [MAX_SUM_WDTH_L-1:0]        I8b12d3b1f65fad05577cf25e8d7950a5;
reg  [MAX_SUM_WDTH_L-1:0]        I488635e3f7ed77ea88199f5bffd4b1d6;
wire [MAX_SUM_WDTH_L-1:0]        Ifb24658924186dba2d1a85ee28fc0313;
reg  [MAX_SUM_WDTH_L-1:0]        Ie6893017d21c050ba10d206854f4a9f4;
wire [MAX_SUM_WDTH_L-1:0]        I067250d29597d7c71da50f8cf557eb61;
reg  [MAX_SUM_WDTH_L-1:0]        Id3f68b4dc0ab60673208b7d2081f3533;
wire [MAX_SUM_WDTH_L-1:0]        Ic86c9a00eacc20772706da9399aab4ba;
reg  [MAX_SUM_WDTH_L-1:0]        I433756b944e061a824a89bda241e879f;
wire [MAX_SUM_WDTH_L-1:0]        I8271913876a2729269e844dc4809a25f;
reg  [MAX_SUM_WDTH_L-1:0]        I2eb60a922aa4f7482dd92b9351d53a2d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3af8e500702e46e7330796cb23979266;
reg  [MAX_SUM_WDTH_L-1:0]        I0867979e1b159c8ceae548930376f482;
wire [MAX_SUM_WDTH_L-1:0]        Ice852e353c55faedcde1922d0179b30a;
reg  [MAX_SUM_WDTH_L-1:0]        I4accfbeae8a5ee0dbeab23ef3a116145;
wire [MAX_SUM_WDTH_L-1:0]        Ibb9864cd5bcd1ef1fc7bfd822db3150b;
reg  [MAX_SUM_WDTH_L-1:0]        Ic7570b0b7c5bef5758f68562ae4c90f6;
wire [MAX_SUM_WDTH_L-1:0]        I13f58835ab9e6362ffddf06976c97207;
reg  [MAX_SUM_WDTH_L-1:0]        Iceadadc4456881fdeea85934a9bf4d6c;
wire [MAX_SUM_WDTH_L-1:0]        I35bfac2d8d88c61e93a27db564f9ecef;
reg  [MAX_SUM_WDTH_L-1:0]        I7b2b617ae67424f54961eebce42de77e;
wire [MAX_SUM_WDTH_L-1:0]        I7ecdf9f7726df27510f35fe6c1b5b4be;
reg  [MAX_SUM_WDTH_L-1:0]        I953f0f8af76f89b2d9ab4abf19fb411d;
wire [MAX_SUM_WDTH_L-1:0]        I7327385650ea109a8bb07f1c92252d28;
reg  [MAX_SUM_WDTH_L-1:0]        I915b4736dcb20f831d02e48f4e79f008;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib5d66de65bb7bc9e1f7b3f05e4bd703b;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7eec587348ae1ca1f00c0a3ad10ad27;
wire [MAX_SUM_WDTH_L-1:0]        Ifca73a480a501ea2636c47e487987167;
reg  [MAX_SUM_WDTH_L-1:0]        I001a212686304248c8359e5fc01227c0;
wire [MAX_SUM_WDTH_L-1:0]        I75a3f16cb4ddc4b0478fb1c07c10aba8;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb7554e012c0fc1223c29b759c900666;
wire [MAX_SUM_WDTH_L-1:0]        I5603979fb76ebb2bab9a8764c4833b52;
reg  [MAX_SUM_WDTH_L-1:0]        I9aeb9c42b54a05be6bf9b7b88b6860ba;
wire [MAX_SUM_WDTH_L-1:0]        I939430bcba9f8bb28f5782040a4c76e7;
reg  [MAX_SUM_WDTH_L-1:0]        I6a5a5966965b0790b906c6fda71aef80;
wire [MAX_SUM_WDTH_L-1:0]        I71ed74fcff44b1a6ec1ddf7b18cf8a31;
reg  [MAX_SUM_WDTH_L-1:0]        Ic943083ca65ace6c42d73f4234739a06;
wire [MAX_SUM_WDTH_L-1:0]        Icc204071ef0dd850f42840be901a1c8c;
reg  [MAX_SUM_WDTH_L-1:0]        Id0b321686d4c39621024cf0dd99822dc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie8187be889aa7f205231e2e60cb827e3;
reg  [MAX_SUM_WDTH_L-1:0]        I0839dd3787442f1b79b87e02436bfdce;
wire [MAX_SUM_WDTH_L-1:0]        I18c57ba0c68acdec8308c2ba40482668;
reg  [MAX_SUM_WDTH_L-1:0]        I89e6a9fd97d8aa4dd3b832c3be4697b2;
wire [MAX_SUM_WDTH_L-1:0]        If45f0a6203e1a6ef6e0d86ccccab3920;
reg  [MAX_SUM_WDTH_L-1:0]        I93d4157f48b132642752220059861e98;
wire [MAX_SUM_WDTH_L-1:0]        I834626bbcdd99143f36052aa6e77de49;
reg  [MAX_SUM_WDTH_L-1:0]        I8fc4faa2891d7fd3479ac1f788f481dc;
wire [MAX_SUM_WDTH_L-1:0]        I58860aa281debf67db1369b2e22b9f5b;
reg  [MAX_SUM_WDTH_L-1:0]        I440f30e9cb4bc89233b46ea00b4cbeb4;
wire [MAX_SUM_WDTH_L-1:0]        I885d19716778193c3288c8322cfd32ae;
reg  [MAX_SUM_WDTH_L-1:0]        I6568bfd8780c11e0b1b049a01f92abd8;
wire [MAX_SUM_WDTH_L-1:0]        I19a6d51c460b600130966b5be281d23e;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf7dc4da07f9955d5d4c7e1f63f1ad68;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I7a4326b2355162700b8647861c80f43f;
reg  [MAX_SUM_WDTH_L-1:0]        I7ec1a328587b72a39c462083efea0ee0;
wire [MAX_SUM_WDTH_L-1:0]        I40ce63d36b1aa901d29c0ecc3ad20a66;
reg  [MAX_SUM_WDTH_L-1:0]        Iaf028e7ab4dc77a7649f15d603834b5f;
wire [MAX_SUM_WDTH_L-1:0]        I32230b8893dd9fd1da4ce1f2553b5550;
reg  [MAX_SUM_WDTH_L-1:0]        I58db79a8e9f0cd1ded379897ba2f27ae;
wire [MAX_SUM_WDTH_L-1:0]        If7fb4fa70b6803a7e4c64a834669dbfa;
reg  [MAX_SUM_WDTH_L-1:0]        I6d3cb4ccb4e51c7e6603d0abd1a082c4;
wire [MAX_SUM_WDTH_L-1:0]        Iaf1e5c8b7267eca64468227734dcfbdb;
reg  [MAX_SUM_WDTH_L-1:0]        I79f75f49ea8a29d684af396014b2f3ab;
wire [MAX_SUM_WDTH_L-1:0]        I5ab38b4a054c50fced80e9323f4a9ddf;
reg  [MAX_SUM_WDTH_L-1:0]        I9c5ecd86bedb189fada40fae9d751a68;
wire [MAX_SUM_WDTH_L-1:0]        I779f57a085e170d2ab7e7b5f046e42e6;
reg  [MAX_SUM_WDTH_L-1:0]        Iad5f06e1989ead7d306c70a3b02cb8f4;
wire [MAX_SUM_WDTH_L-1:0]        I120e630331e23d75054584a44aafaf63;
reg  [MAX_SUM_WDTH_L-1:0]        If6d1a410df5a4aea6a01337a6074fbd9;
wire [MAX_SUM_WDTH_L-1:0]        I3f690a6c75649328d7cccf08cc6ca81b;
reg  [MAX_SUM_WDTH_L-1:0]        I3bc40a4db14566b5099b14cee5f61135;
wire [MAX_SUM_WDTH_L-1:0]        I2105fce588dc6840254a1eaf02b549c9;
reg  [MAX_SUM_WDTH_L-1:0]        I7e683fd8235d7cfbf4ff407a286f07de;
wire [MAX_SUM_WDTH_L-1:0]        Ic0b28cd43f561513b63ff20e31038f37;
reg  [MAX_SUM_WDTH_L-1:0]        I97afcedf05e588b7976d6005191dc916;
wire [MAX_SUM_WDTH_L-1:0]        Ib4e0926a64eaefff0e36fdde4783e923;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8d8eec0aaa662adf2837c9b705fce7e;
wire [MAX_SUM_WDTH_L-1:0]        Ieb485d7a868decbc901fad618f56412a;
reg  [MAX_SUM_WDTH_L-1:0]        Icbd765be950123705955e2c5d7ace84b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I71853033c5b7e4e98414209075b4d708;
reg  [MAX_SUM_WDTH_L-1:0]        I706e8f5617cfae1e6fc83db18c8b5fe3;
wire [MAX_SUM_WDTH_L-1:0]        I37621b4bc9c88a42a47d3123465fa4d5;
reg  [MAX_SUM_WDTH_L-1:0]        I1dd8f8c7f1b673898096b1f3ae383197;
wire [MAX_SUM_WDTH_L-1:0]        Ied0d483617ee30ac0539009fba84a684;
reg  [MAX_SUM_WDTH_L-1:0]        I10ca8978cf4659265ed25a27d09acc1c;
wire [MAX_SUM_WDTH_L-1:0]        I574d31b300f16225a707bbae0918c445;
reg  [MAX_SUM_WDTH_L-1:0]        Iec4656b32460def4a608b6b0f6486af9;
wire [MAX_SUM_WDTH_L-1:0]        I9fef812393d8a5f87abc46add3371777;
reg  [MAX_SUM_WDTH_L-1:0]        I5f4475897d1d58965da1b35fe0ef8c01;
wire [MAX_SUM_WDTH_L-1:0]        I64a11eacbd9a28d7e65c56c38127876b;
reg  [MAX_SUM_WDTH_L-1:0]        Ife61469306df3cf220666b187f1496a9;
wire [MAX_SUM_WDTH_L-1:0]        Id11f93a74e2de2ea1e27e9d2858a472f;
reg  [MAX_SUM_WDTH_L-1:0]        Ib49319b9dfa4914f92f423ceaf840014;
wire [MAX_SUM_WDTH_L-1:0]        Ibd0708af1cccb49fded84694d6ffd6f7;
reg  [MAX_SUM_WDTH_L-1:0]        I93ff2f879233cac9b9f0dd2f4c082c09;
wire [MAX_SUM_WDTH_L-1:0]        I18edce191243df3a622232f681b7e3f9;
reg  [MAX_SUM_WDTH_L-1:0]        I44597d694e9c5d29280e503d72a27c8d;
wire [MAX_SUM_WDTH_L-1:0]        Ib68ae994fc94acf008e424d8f8c8eb4b;
reg  [MAX_SUM_WDTH_L-1:0]        I04a19448c5e75af8021ad02d1a708bb0;
wire [MAX_SUM_WDTH_L-1:0]        Icb6bc0221ed78051fa10967f5cce4a7f;
reg  [MAX_SUM_WDTH_L-1:0]        I71a3093121c2f19dcd1412b468652fa8;
wire [MAX_SUM_WDTH_L-1:0]        I3abb9a64f85be533ac16eafaf85c5ad1;
reg  [MAX_SUM_WDTH_L-1:0]        I3ae09c82029c617034fe6aacbe9e94e6;
wire [MAX_SUM_WDTH_L-1:0]        If6badde34faca49e04b3dde9b11c0556;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7af6b3b441f910b000a333afad6c76f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I09d6aa4053f5e1280d70556ad1cc89a4;
reg  [MAX_SUM_WDTH_L-1:0]        I4d71dfea8407aa5b5cbb991bc4fea963;
wire [MAX_SUM_WDTH_L-1:0]        I9d1f949ca74fcf76431906a3a95d4866;
reg  [MAX_SUM_WDTH_L-1:0]        I1a082caecc831a90e74674ba35da4183;
wire [MAX_SUM_WDTH_L-1:0]        I10221054a7689d49c97a1e908e2fb44b;
reg  [MAX_SUM_WDTH_L-1:0]        Iec1de44616a2354a56ab1f681059d4c5;
wire [MAX_SUM_WDTH_L-1:0]        I4ec67f577ac5c95d8a93f21935a4fb7f;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3c2318e64d0e218c3db557404c4aac8;
wire [MAX_SUM_WDTH_L-1:0]        I069f6a3e5c61b47031648ed6e7ab0330;
reg  [MAX_SUM_WDTH_L-1:0]        I9a251d50f41e51b1a5cc2475f267e8a0;
wire [MAX_SUM_WDTH_L-1:0]        I4b15910b07c427bfb666057cf4700947;
reg  [MAX_SUM_WDTH_L-1:0]        I9b5767a49f7b9dcb8fdaea924835033c;
wire [MAX_SUM_WDTH_L-1:0]        I5694aa90f55816a9ca217470b70f29a6;
reg  [MAX_SUM_WDTH_L-1:0]        I6ca1e6700a19d03621a193c7240bff54;
wire [MAX_SUM_WDTH_L-1:0]        Ia1d3638756959bfb67f32a37c58fe190;
reg  [MAX_SUM_WDTH_L-1:0]        I931c597ff12bffce581f653346202f83;
wire [MAX_SUM_WDTH_L-1:0]        I3e81666362b0209c98c5337a74dcbfa9;
reg  [MAX_SUM_WDTH_L-1:0]        Ia3a2c5d59f6340917ca3933c05ba4678;
wire [MAX_SUM_WDTH_L-1:0]        Iaa723368e8f531ae9bf99c9b99fdf0f7;
reg  [MAX_SUM_WDTH_L-1:0]        Ie83d0a8ee5ed214bc7577467748aaa04;
wire [MAX_SUM_WDTH_L-1:0]        I3713f644fba6dd9d4bb4dc3b4c91fe77;
reg  [MAX_SUM_WDTH_L-1:0]        Iaac29552e5fc65aaf4f0116f917b707c;
wire [MAX_SUM_WDTH_L-1:0]        I5a3e3131db6fdd74e5c822fde6a8f2c1;
reg  [MAX_SUM_WDTH_L-1:0]        Ie2c8eac7204b98139c03b6fbfff9af36;
wire [MAX_SUM_WDTH_L-1:0]        If18033df3d6ee029fdecf3323ad8d62d;
reg  [MAX_SUM_WDTH_L-1:0]        Ied7fcdaec662cb3c2f89f131986fa102;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I7514cd65da98bd214b4e1da34ac358f1;
reg  [MAX_SUM_WDTH_L-1:0]        Ib16a17d6430570b45a304d847ee2b11c;
wire [MAX_SUM_WDTH_L-1:0]        Id947f3ca55c826ef94d1ac4ad2a227bf;
reg  [MAX_SUM_WDTH_L-1:0]        I42169e454756fe4d1c5f17f2eeb2e091;
wire [MAX_SUM_WDTH_L-1:0]        Ia6f83033bc647143bbf5377056c7072f;
reg  [MAX_SUM_WDTH_L-1:0]        I6fde38a3a92e06fa77123e3279813c41;
wire [MAX_SUM_WDTH_L-1:0]        I21dd15d84c5abe8d2ac53f65236f587c;
reg  [MAX_SUM_WDTH_L-1:0]        Id8ee16437e8d6d6da6d37440e04097b6;
wire [MAX_SUM_WDTH_L-1:0]        Ia88c70253514b080daa27d2df0aef202;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf249d8e5acced9b064132575f40e001;
wire [MAX_SUM_WDTH_L-1:0]        I3cd11d85b17ce4c2181dfd2430ff4595;
reg  [MAX_SUM_WDTH_L-1:0]        I580659084e3d17b48de6b1c66154fcf5;
wire [MAX_SUM_WDTH_L-1:0]        I9817361d029cc98d7407cf3b8b020567;
reg  [MAX_SUM_WDTH_L-1:0]        I7a14e45d43ab77b265501902152c8616;
wire [MAX_SUM_WDTH_L-1:0]        I47a6f2033a2356ac604133d12d7e0c0e;
reg  [MAX_SUM_WDTH_L-1:0]        I81ba868784103e0eb05a44d981d4d666;
wire [MAX_SUM_WDTH_L-1:0]        I3da1998324eb1853e5ec747b112095aa;
reg  [MAX_SUM_WDTH_L-1:0]        Ic6b88783957cbaf253648a30b22f6b1c;
wire [MAX_SUM_WDTH_L-1:0]        Ic729cdba5f8a3933121a0ef35da99f8c;
reg  [MAX_SUM_WDTH_L-1:0]        I4103c218a85a1d08db5c4f4b5686b2e5;
wire [MAX_SUM_WDTH_L-1:0]        Id7542fd1fe3a099d7274f15c008f1cc5;
reg  [MAX_SUM_WDTH_L-1:0]        I0e6c0958af503e4a120a49d02a432863;
wire [MAX_SUM_WDTH_L-1:0]        I1a91347d29cd64af8941a3e042228a52;
reg  [MAX_SUM_WDTH_L-1:0]        I8f76b31e8f15c0e5fe24dcb723418111;
wire [MAX_SUM_WDTH_L-1:0]        Ic6b16867c426103b3e53db94469de2cb;
reg  [MAX_SUM_WDTH_L-1:0]        Id1457221b58344b60070aa026436df2c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I7361a720882c68965c1c28c2d6ba1dff;
reg  [MAX_SUM_WDTH_L-1:0]        Icc31966508e03d8869e81d8aeb243705;
wire [MAX_SUM_WDTH_L-1:0]        I668a239256c66a858129b4788b0001a5;
reg  [MAX_SUM_WDTH_L-1:0]        I9dcccf542ba434b6e0fde6f012f98f92;
wire [MAX_SUM_WDTH_L-1:0]        I73a72fba51f575f80ded2357a6b71af0;
reg  [MAX_SUM_WDTH_L-1:0]        I51ccbb824a5e1e340eefd173c4491728;
wire [MAX_SUM_WDTH_L-1:0]        Ief9131d8e69f733c51e9f9167ad5fa4a;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7ae1730dcd8bc708bbfcc6a9f97ac66;
wire [MAX_SUM_WDTH_L-1:0]        I1e6904544c93f0f4bf403793e50dbf99;
reg  [MAX_SUM_WDTH_L-1:0]        I4714f5c91203fcfa552f0fcf71b87442;
wire [MAX_SUM_WDTH_L-1:0]        I74f9e6de534920d70eda17b59206a4af;
reg  [MAX_SUM_WDTH_L-1:0]        I3b6d1e84fdd1019249886fa5fe65895b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ied74515bab35cad5e94048a9f210b7a5;
reg  [MAX_SUM_WDTH_L-1:0]        Ia8a7d4207dbabc7970bf36f3fe74f72d;
wire [MAX_SUM_WDTH_L-1:0]        If38f871a7b021ceb84cdb3010d08f667;
reg  [MAX_SUM_WDTH_L-1:0]        I84047457b43ef33874f4550c3b773460;
wire [MAX_SUM_WDTH_L-1:0]        I12a578d51082c42fcc5a9e769535ac0a;
reg  [MAX_SUM_WDTH_L-1:0]        I5e51563c3e69beca0b463742e6e5f9ee;
wire [MAX_SUM_WDTH_L-1:0]        I404f31fea404e730a9c4e04bec369c1a;
reg  [MAX_SUM_WDTH_L-1:0]        I6c8d14e31c80811ccab1b6ab09d28089;
wire [MAX_SUM_WDTH_L-1:0]        I915d15cb464b6e78cf9939232618b14c;
reg  [MAX_SUM_WDTH_L-1:0]        I50b3b7490c9b65b6e662cc86b163a2df;
wire [MAX_SUM_WDTH_L-1:0]        Ia8531e691cc60dcc32225eef6d8e8a2b;
reg  [MAX_SUM_WDTH_L-1:0]        I8351a2110a3d73ad8803cf17e3317017;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5f7cd38f8b6c42a3dcc52664ea7c08a5;
reg  [MAX_SUM_WDTH_L-1:0]        I1e6c696951688d581f21ab2302593335;
wire [MAX_SUM_WDTH_L-1:0]        If3f0f6acad563083949c5116ad78ce20;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9840e28133eebdca0be313552195c7b;
wire [MAX_SUM_WDTH_L-1:0]        I2b8c7ab8f53d7fbda984ab8760e05fd3;
reg  [MAX_SUM_WDTH_L-1:0]        I82812258a8032e273cab7139266be1b6;
wire [MAX_SUM_WDTH_L-1:0]        I29d486911dcffddec336f69b981e1e50;
reg  [MAX_SUM_WDTH_L-1:0]        I27ab6fd9927518e29ed36d7a7a241498;
wire [MAX_SUM_WDTH_L-1:0]        I893881a7874f85e519089559ac4604bf;
reg  [MAX_SUM_WDTH_L-1:0]        I05b0f33a3808ac53b29d8d8309447650;
wire [MAX_SUM_WDTH_L-1:0]        I0b730d0a75cf72482ffc5b0d0267fd83;
reg  [MAX_SUM_WDTH_L-1:0]        If150ebf242231f0d22c996a71552f6eb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I9beb581fcdf85cc7302da093363e3b02;
reg  [MAX_SUM_WDTH_L-1:0]        If2d0a2b58510715e74787cb60719cb5b;
wire [MAX_SUM_WDTH_L-1:0]        I0e35fb521572c6f87dbd06a8ce213337;
reg  [MAX_SUM_WDTH_L-1:0]        Ib6745a6d17034a29501e022bd846bf2f;
wire [MAX_SUM_WDTH_L-1:0]        Ia01e93b03cf0ff22e2f002f2e84eb9d2;
reg  [MAX_SUM_WDTH_L-1:0]        Iae09c127dfe86c9f7bdbeff447c777f5;
wire [MAX_SUM_WDTH_L-1:0]        I98a2d427581a73c639cbc9f4bf4c8802;
reg  [MAX_SUM_WDTH_L-1:0]        I742128de6b237ed48e3a7ccd3788f0d7;
wire [MAX_SUM_WDTH_L-1:0]        Ie60ba6ee53f7a01764001bc74fb90d61;
reg  [MAX_SUM_WDTH_L-1:0]        Id5e8fda13ba8f6d95d694d0f30da75bb;
wire [MAX_SUM_WDTH_L-1:0]        I508e632bacf8c083a8376f73cec11bc6;
reg  [MAX_SUM_WDTH_L-1:0]        I1aa5a04e40f9b1685c77e4d101c3ccf4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I47ac3c977bbfad06ee1782b8eac6d9ec;
reg  [MAX_SUM_WDTH_L-1:0]        Ife1adea26d13bc299bb2de241ad4a6ea;
wire [MAX_SUM_WDTH_L-1:0]        If8537bb117e0bebd25ece101a23674c8;
reg  [MAX_SUM_WDTH_L-1:0]        Ifcf6c761f0f253921710af87ab1d2247;
wire [MAX_SUM_WDTH_L-1:0]        Ica8f952cb456e825c608f2e73ec9abd7;
reg  [MAX_SUM_WDTH_L-1:0]        I1478e6a9113c124bdc4361908af6643f;
wire [MAX_SUM_WDTH_L-1:0]        I1a332ceae6f1a640e4577c82b2bf4511;
reg  [MAX_SUM_WDTH_L-1:0]        I0afd42151925883835844cf5deef6156;
wire [MAX_SUM_WDTH_L-1:0]        I82c5b5deaae0b927c14adfa3b477c8df;
reg  [MAX_SUM_WDTH_L-1:0]        I2b4ab0aadffb3a1bb86f45ebc8acf085;
wire [MAX_SUM_WDTH_L-1:0]        I37b08ee3258fb8359ba4c1653101e03c;
reg  [MAX_SUM_WDTH_L-1:0]        Iffa867719ba9c31a8756cc5e6bf81147;
wire [MAX_SUM_WDTH_L-1:0]        I58fa785303fe60b1f1c596420aab4b5e;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb62b6cb003f0d5549c864075f23d19b;
wire [MAX_SUM_WDTH_L-1:0]        I1ceca376c3f4cd24c22cf8672c9343ba;
reg  [MAX_SUM_WDTH_L-1:0]        I3690d101ae99f258cc58b4482cc378c8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ieca948a12a0806b9fd483ace71c8b98e;
reg  [MAX_SUM_WDTH_L-1:0]        Id597e95ce8a168ab67890085a26870d0;
wire [MAX_SUM_WDTH_L-1:0]        Icd2579fee72faaa432876ec8fa124d40;
reg  [MAX_SUM_WDTH_L-1:0]        I98df60eb8f65641f9cccce4023be905c;
wire [MAX_SUM_WDTH_L-1:0]        Iec4164641d5b71630d9d5aefb1ed5676;
reg  [MAX_SUM_WDTH_L-1:0]        Ibcb4fbdee372353b79c460cdeafdfe4e;
wire [MAX_SUM_WDTH_L-1:0]        Ie43841b2ee3b5369c3863417b60e5851;
reg  [MAX_SUM_WDTH_L-1:0]        I74dbf75966d047a4a9e91c1bc793666f;
wire [MAX_SUM_WDTH_L-1:0]        I1e7346a531973e40fb2582a68f96e383;
reg  [MAX_SUM_WDTH_L-1:0]        I79b8d9f9447c4c1b551ec6c1e8903040;
wire [MAX_SUM_WDTH_L-1:0]        I53b62438d1bb777cf10761bf95b22718;
reg  [MAX_SUM_WDTH_L-1:0]        Ib34b66548621fabe0753223712b1369f;
wire [MAX_SUM_WDTH_L-1:0]        I6b8a0d9d8fe6ac6fa08c495b0d0d5264;
reg  [MAX_SUM_WDTH_L-1:0]        Ie5b3eb4c00bedfaecc3215d43ff28362;
wire [MAX_SUM_WDTH_L-1:0]        Ibcec436bb431239047a99c495262bf87;
reg  [MAX_SUM_WDTH_L-1:0]        Icf3a1b0b6dbcf959b44379024f3c4169;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Id9d1f164781aad87bbb332ef7c0b5113;
reg  [MAX_SUM_WDTH_L-1:0]        I918c2bbe7c71f8c6a07b0bad8811f4e7;
wire [MAX_SUM_WDTH_L-1:0]        I76a91ad2a7f0323b5874f857eb914d67;
reg  [MAX_SUM_WDTH_L-1:0]        Iedd960a21b1c08b4a5293cff200218b3;
wire [MAX_SUM_WDTH_L-1:0]        I9aab2781bbd57dbe4381c695f130d5b7;
reg  [MAX_SUM_WDTH_L-1:0]        If9722c28747df3a59b0ecf8200907e98;
wire [MAX_SUM_WDTH_L-1:0]        I11c62ef31300f66f787bb7285596b995;
reg  [MAX_SUM_WDTH_L-1:0]        Ib83df72c8b73a333d0699a8bbbec16be;
wire [MAX_SUM_WDTH_L-1:0]        I7e62705e1f1e7abb04ee4a94753183b4;
reg  [MAX_SUM_WDTH_L-1:0]        Ide3798a77f709a9f694523338b081f70;
wire [MAX_SUM_WDTH_L-1:0]        Ia4d8ab77dd8598d550c4b3c57f02b328;
reg  [MAX_SUM_WDTH_L-1:0]        I0a9722a805604433562f85c62b168b96;
wire [MAX_SUM_WDTH_L-1:0]        I23c2886f2707bae85fe967379c105eb5;
reg  [MAX_SUM_WDTH_L-1:0]        If9480ec13cd538ed03a43e56bd6264a6;
wire [MAX_SUM_WDTH_L-1:0]        Idfb980ae7487145d65bdf83b97751e6f;
reg  [MAX_SUM_WDTH_L-1:0]        I433ecf86b7704c5552e5fb5cafe0d529;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If7916cdab9aa2621009bc0671d985133;
reg  [MAX_SUM_WDTH_L-1:0]        I8326f0b2d25139609e2c5e466724f224;
wire [MAX_SUM_WDTH_L-1:0]        I1969f6d312f67452ec24690813fc07ae;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbe211d9955cdf2810c9003d1fb78074;
wire [MAX_SUM_WDTH_L-1:0]        I6b3c96ebbba2bfe8c549caea4a266656;
reg  [MAX_SUM_WDTH_L-1:0]        If15e950b569a92b590127d0ca6f20a16;
wire [MAX_SUM_WDTH_L-1:0]        I73172f8b4bcb0bdbe27a09cd7ec204e0;
reg  [MAX_SUM_WDTH_L-1:0]        I03e0532841ba39eb1d4ae823c4de2f7d;
wire [MAX_SUM_WDTH_L-1:0]        I96acfb8f7e6c42f616a880b3657f42a9;
reg  [MAX_SUM_WDTH_L-1:0]        I1be81a7b73987ee023e396cec87312d1;
wire [MAX_SUM_WDTH_L-1:0]        I5cdce64ba621df381f9efbb8b0c8e10a;
reg  [MAX_SUM_WDTH_L-1:0]        I4ce1a767a78673590c4074f3f03bad8d;
wire [MAX_SUM_WDTH_L-1:0]        I61389621065261b79f16e6dae7c7cdac;
reg  [MAX_SUM_WDTH_L-1:0]        I57806bb7da625881e68ae315543f70d6;
wire [MAX_SUM_WDTH_L-1:0]        Ide44caca4eb1b6edc9b55c584239ff94;
reg  [MAX_SUM_WDTH_L-1:0]        I8b0ab476b4790150575abb06bcdce2b3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I892e07e7e972dd521f273519694e4ee7;
reg  [MAX_SUM_WDTH_L-1:0]        I8846a8961b7d557df4fc62dada679c33;
wire [MAX_SUM_WDTH_L-1:0]        I43c8950bb200a93cec12c09af4a38dae;
reg  [MAX_SUM_WDTH_L-1:0]        I7909a0f96a92e93f95023cddc742a5eb;
wire [MAX_SUM_WDTH_L-1:0]        I591f0a636f176d5a398cb6ed6d67f627;
reg  [MAX_SUM_WDTH_L-1:0]        I43ac4857544c0fb79d04e850435ef673;
wire [MAX_SUM_WDTH_L-1:0]        I8be467496bf21fa2c46fc5db2442a339;
reg  [MAX_SUM_WDTH_L-1:0]        Ia6dfa47c465325c1d9fb9b9c5ce08f01;
wire [MAX_SUM_WDTH_L-1:0]        Ifa0294e878bf5a4f1c6c7cfa52c46e7d;
reg  [MAX_SUM_WDTH_L-1:0]        I2e9eda5bea0cc3d88359ce8a7a82f21f;
wire [MAX_SUM_WDTH_L-1:0]        I35a8b04ecb2c6d2d7bd52a64010038ff;
reg  [MAX_SUM_WDTH_L-1:0]        I53ec2486418e41b2ccfa8fd82777eaf0;
wire [MAX_SUM_WDTH_L-1:0]        I38629158c9fc8600b05a3e32589cbeda;
reg  [MAX_SUM_WDTH_L-1:0]        I18387c05cef21970ecbc39c20a87aafb;
wire [MAX_SUM_WDTH_L-1:0]        Ie20705331f5fabb4c9f720a5c6592c7d;
reg  [MAX_SUM_WDTH_L-1:0]        I2b23eae78cb925008ad59f45e80e165b;
wire [MAX_SUM_WDTH_L-1:0]        I425d66a6ead3859f364e20a797b0e4e2;
reg  [MAX_SUM_WDTH_L-1:0]        Ic69eb7677638a90b7a54389d47be46de;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I66a2577a791bae1f31c5b99b0c3f324d;
reg  [MAX_SUM_WDTH_L-1:0]        I8cb9a216f4da7c27f678386cb214c59d;
wire [MAX_SUM_WDTH_L-1:0]        I77350e171f060c2d49e50c636fab084f;
reg  [MAX_SUM_WDTH_L-1:0]        I48cb720a6323697084ac3bbd8fcadfcb;
wire [MAX_SUM_WDTH_L-1:0]        I2101d085d5e55ef5b8247de3898a80e7;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8dc3c1885c92cdcce7fcb58d65d03e7;
wire [MAX_SUM_WDTH_L-1:0]        Id38879e0d52fba6818597bd60dfc2b2c;
reg  [MAX_SUM_WDTH_L-1:0]        Ic3aa51a5c758405fa6e2dbed707555b2;
wire [MAX_SUM_WDTH_L-1:0]        I68081efdf01e540fe5e07643a2bc3463;
reg  [MAX_SUM_WDTH_L-1:0]        I4d418179c859feb8bc7d750416bb1004;
wire [MAX_SUM_WDTH_L-1:0]        I2d70e6f392396c2ee505687f5a950a6f;
reg  [MAX_SUM_WDTH_L-1:0]        If207b2adc6f668f85cb76bf54673fe18;
wire [MAX_SUM_WDTH_L-1:0]        I6e6eae8e8a955b80abb7cb722a940e27;
reg  [MAX_SUM_WDTH_L-1:0]        Ib08b8067ea75e210e83526ca4a37217e;
wire [MAX_SUM_WDTH_L-1:0]        I54cfd5f12219687ba48be0c57a979add;
reg  [MAX_SUM_WDTH_L-1:0]        I95b30f641cbf7bec1886643c4468017d;
wire [MAX_SUM_WDTH_L-1:0]        Ifda70e49dbdc4b5511961649914ecc71;
reg  [MAX_SUM_WDTH_L-1:0]        I1978531a6f8d1d25ee6d404025ec4753;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0feba37f523d6c6371bd934796519c59;
reg  [MAX_SUM_WDTH_L-1:0]        I6c9698ba88db16b8d22ccebd58cc541d;
wire [MAX_SUM_WDTH_L-1:0]        Ibaf70dff036e0bc11df75e2a1fe4fb34;
reg  [MAX_SUM_WDTH_L-1:0]        I0d8ac5e09b200a55bf5ba6f834cc9174;
wire [MAX_SUM_WDTH_L-1:0]        Ib00eb8856f044c3af325f0134d16a970;
reg  [MAX_SUM_WDTH_L-1:0]        Ib58b7d3d77a54ff1a180c6fa5f1400e6;
wire [MAX_SUM_WDTH_L-1:0]        I4e89f11e414b55e9574f5c3d79dc4506;
reg  [MAX_SUM_WDTH_L-1:0]        Icf6b990098b7ab91800bfcf1e643153c;
wire [MAX_SUM_WDTH_L-1:0]        If25b7447f1f34072a597f70a4234a16e;
reg  [MAX_SUM_WDTH_L-1:0]        Ie4308b9ac6fb6de9329ba02b1eeb0e8a;
wire [MAX_SUM_WDTH_L-1:0]        I76ae0b929aefad162304529ea04b725f;
reg  [MAX_SUM_WDTH_L-1:0]        I01d4f02a356c51d7e4e1993de0d8eebd;
wire [MAX_SUM_WDTH_L-1:0]        Idffaf5edec0ef7b25c24f3c5e636fb75;
reg  [MAX_SUM_WDTH_L-1:0]        I36c351e3641b01cc43e1dd5de0a649e5;
wire [MAX_SUM_WDTH_L-1:0]        Id041de10db620915a3755358fc2d9a41;
reg  [MAX_SUM_WDTH_L-1:0]        I4fc983e94c5b8f7bafca61fb0d351c08;
wire [MAX_SUM_WDTH_L-1:0]        I92ddd31add3c914ce6b0271e77cb67a0;
reg  [MAX_SUM_WDTH_L-1:0]        I1fcb82fdf96cda14a55fa6358cb62c1e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If80ebbd3419cd9fd63a745412b7233b6;
reg  [MAX_SUM_WDTH_L-1:0]        I665e54ea6bdca483149d3b7f3ee42a2b;
wire [MAX_SUM_WDTH_L-1:0]        I0b67c1f8e03165404e0b76d1a05d88de;
reg  [MAX_SUM_WDTH_L-1:0]        I925df2307b5af6d1b166e5435641d3bd;
wire [MAX_SUM_WDTH_L-1:0]        If78c15d7c2dc19cef26743eccbb52e6c;
reg  [MAX_SUM_WDTH_L-1:0]        I9b14f48aa357d09e460a445da86cdf89;
wire [MAX_SUM_WDTH_L-1:0]        I228c0b3c3919aaf70ea24874f314eaa5;
reg  [MAX_SUM_WDTH_L-1:0]        I78e94ecb6c92fa8ee24edaff33b6f82d;
wire [MAX_SUM_WDTH_L-1:0]        I986ca3b0590709588c3d9d2274a1fd34;
reg  [MAX_SUM_WDTH_L-1:0]        I5ebeb9ce5adee72a7c9527ea6d3a3028;
wire [MAX_SUM_WDTH_L-1:0]        I765867ea6452d51f31e96ec83f68f9df;
reg  [MAX_SUM_WDTH_L-1:0]        I90d7b28ec09142ca8086836fc0c5ea0d;
wire [MAX_SUM_WDTH_L-1:0]        I6e970e7bafbfa1866203483ed18a7db7;
reg  [MAX_SUM_WDTH_L-1:0]        I27d9985415e6d0b117e5a4c2863aa7f8;
wire [MAX_SUM_WDTH_L-1:0]        Ia31bbc3e099eb2180960917330d6b2e1;
reg  [MAX_SUM_WDTH_L-1:0]        Idf9b563e5d10c2bdbcc07e81d74467eb;
wire [MAX_SUM_WDTH_L-1:0]        Ibc94d96e529274004dfed98c98915827;
reg  [MAX_SUM_WDTH_L-1:0]        Ie351922194483938302ff6cafc477e4a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I60eb0a19c8d75780a4dae7d33ba46bd4;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb2da5faf236ca8636677bc1dc35c4db;
wire [MAX_SUM_WDTH_L-1:0]        I701ff10dac46e4482b3bcaa387c9a725;
reg  [MAX_SUM_WDTH_L-1:0]        Ie15825d216685ae241b528fa9c158ff3;
wire [MAX_SUM_WDTH_L-1:0]        Ifd170f2b9fa5df9a7d0817307b5586a2;
reg  [MAX_SUM_WDTH_L-1:0]        Id92c2d8bc61245c0c8e40bec2424c3c8;
wire [MAX_SUM_WDTH_L-1:0]        Ia5feb8ce451f12382cb66853e948047d;
reg  [MAX_SUM_WDTH_L-1:0]        Icd9fd8d7114b6e894dbee493b6797df6;
wire [MAX_SUM_WDTH_L-1:0]        I3a971f30fe10de02e604402b55c181da;
reg  [MAX_SUM_WDTH_L-1:0]        I29ff688c085f2b18e7a3af969f18af76;
wire [MAX_SUM_WDTH_L-1:0]        I3350d782125dfaa1c32d06e6ede68e0f;
reg  [MAX_SUM_WDTH_L-1:0]        I6d56db9fcfe69dfcd747521a1ff62297;
wire [MAX_SUM_WDTH_L-1:0]        Ia07581cdc470c8ba833acbc8a58f7d0e;
reg  [MAX_SUM_WDTH_L-1:0]        I2f17f7c79a0118b39a63894917c6affa;
wire [MAX_SUM_WDTH_L-1:0]        Id91d824405f52636dc30344bf8c088ec;
reg  [MAX_SUM_WDTH_L-1:0]        I7350af5d5ee09ad28c459e3674a829ab;
wire [MAX_SUM_WDTH_L-1:0]        I36beed9320665d5988556ea089ee26f8;
reg  [MAX_SUM_WDTH_L-1:0]        I67b6415c5135e3d6a41d56d98d3f8315;
wire [MAX_SUM_WDTH_L-1:0]        If05d018c797e7d4348fe5bd5423b23cb;
reg  [MAX_SUM_WDTH_L-1:0]        I4a6fffd8bb7244599383f2aa3a1c8916;
wire [MAX_SUM_WDTH_L-1:0]        Ia78ed58e20602b99c01f2208cec79dfd;
reg  [MAX_SUM_WDTH_L-1:0]        I7dbcd21016231546b76aab175cac9f74;
wire [MAX_SUM_WDTH_L-1:0]        I229890d0e3576523fabea29f8594a853;
reg  [MAX_SUM_WDTH_L-1:0]        I9aeff3dc44ed0d0f32518590a900dcc9;
wire [MAX_SUM_WDTH_L-1:0]        I3f0ac12bf9d4014f5418383146bcc1ab;
reg  [MAX_SUM_WDTH_L-1:0]        I988b7d5d56d22d2c77c5c8c125129a50;
wire [MAX_SUM_WDTH_L-1:0]        I38e35040b0a7e5476f308d265b7fbf67;
reg  [MAX_SUM_WDTH_L-1:0]        Iff35cd97f2a6d37a7861b9cc1a655ef5;
wire [MAX_SUM_WDTH_L-1:0]        I90c35b33579355f50d23995dc25cc2af;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb3f2a1bedfe41c73d198046a2a3f177;
wire [MAX_SUM_WDTH_L-1:0]        I19a71e86490479795328e31521b6b842;
reg  [MAX_SUM_WDTH_L-1:0]        I37ddc6ccbc188a3eb8c33a501de820be;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5505d84d5ef89111fd375ce986e33c52;
reg  [MAX_SUM_WDTH_L-1:0]        Ica608f1136da397e2ab61bd4a5d83201;
wire [MAX_SUM_WDTH_L-1:0]        Ie47404148e49f0bfa2775b3573dee999;
reg  [MAX_SUM_WDTH_L-1:0]        I80636a3df4541bf29780bcb4d0ee48f9;
wire [MAX_SUM_WDTH_L-1:0]        Ibae1afc3891aaf6fa2751a693cbf5e1c;
reg  [MAX_SUM_WDTH_L-1:0]        I9ad99d544187db3cc7090b92c9933a31;
wire [MAX_SUM_WDTH_L-1:0]        Icbc45a900f0692fde798caa8c1b9b223;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa8a2b6fcd469869efcf0b75ca38e68f;
wire [MAX_SUM_WDTH_L-1:0]        Ib8aaa1d409ba2d09187c3cf4ad4a1fec;
reg  [MAX_SUM_WDTH_L-1:0]        I9a171d2d8eee362a0073ab7b139d3037;
wire [MAX_SUM_WDTH_L-1:0]        I6a97c95991e02e0e36ec0a1f7c006626;
reg  [MAX_SUM_WDTH_L-1:0]        I84cdcba86bc5991feb391003cd7be40b;
wire [MAX_SUM_WDTH_L-1:0]        I30c34fb37caafa3e5870ae3ee43693c1;
reg  [MAX_SUM_WDTH_L-1:0]        If9e5c3a848acce5daf570458f78f6aad;
wire [MAX_SUM_WDTH_L-1:0]        I8f23d2c62e919062678a00aa98eff7ea;
reg  [MAX_SUM_WDTH_L-1:0]        I73247d4348333f67a491fc607b15af0e;
wire [MAX_SUM_WDTH_L-1:0]        Iaddc9a87ebf5cfb7bbabe07260c592b1;
reg  [MAX_SUM_WDTH_L-1:0]        I021c745eee4b85a2cd91d9d8d2b18b2c;
wire [MAX_SUM_WDTH_L-1:0]        I24abea8ce306ff137aabea504932da94;
reg  [MAX_SUM_WDTH_L-1:0]        I1381c0a0bd28b1c5542992084635b355;
wire [MAX_SUM_WDTH_L-1:0]        Ibee212f9caef9ff8a725aa08e2e955bf;
reg  [MAX_SUM_WDTH_L-1:0]        Ie74eeddc21428254a8fc4c3e293b5eb7;
wire [MAX_SUM_WDTH_L-1:0]        Ie62effeaea232e1a8a50ac3f744f3f3b;
reg  [MAX_SUM_WDTH_L-1:0]        Ib1d0f94258b45de4bfe610086d8990c5;
wire [MAX_SUM_WDTH_L-1:0]        I6712564d12398f5407fade724db8792c;
reg  [MAX_SUM_WDTH_L-1:0]        I138d6d5d60df37870cdbb1d9c51a94af;
wire [MAX_SUM_WDTH_L-1:0]        I5a699ad31ee84bb49eff73572bcaf84a;
reg  [MAX_SUM_WDTH_L-1:0]        I706378735e63e15c8d5395446ea41db8;
wire [MAX_SUM_WDTH_L-1:0]        I63f0b04113e2c8b0cf0474f8aa4fc1cb;
reg  [MAX_SUM_WDTH_L-1:0]        If8680a7fc4f5532a660006bf4ca6a66e;
wire [MAX_SUM_WDTH_L-1:0]        I0dd55598c5774df690bb002eefd62dae;
reg  [MAX_SUM_WDTH_L-1:0]        Ic59d1ff3051a95166c3c2d5a2881221b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I361cee04efb7ccdb28fbf44a7f9c3467;
reg  [MAX_SUM_WDTH_L-1:0]        I54a551af28c505601cdfaf8faaa94afb;
wire [MAX_SUM_WDTH_L-1:0]        I26225a10fd6209094b91ed34531ca2b4;
reg  [MAX_SUM_WDTH_L-1:0]        I6a3124c03eb83d41c16704133bd1cfde;
wire [MAX_SUM_WDTH_L-1:0]        Ib269184699c52eafef7d54ca1fda31d7;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9ee27b9761af611ab96f0010abd47a3;
wire [MAX_SUM_WDTH_L-1:0]        I586e24737da989e9591444e6d260cc9c;
reg  [MAX_SUM_WDTH_L-1:0]        I305436919f84066a22ab1417ebabd737;
wire [MAX_SUM_WDTH_L-1:0]        I01fe0c5ce70d18bdced623e1bfeb55c4;
reg  [MAX_SUM_WDTH_L-1:0]        I78e63717f436493b756efa32d66cdefd;
wire [MAX_SUM_WDTH_L-1:0]        I31e6b870600dcb417653fd673d0c1a55;
reg  [MAX_SUM_WDTH_L-1:0]        Ic965ba971642db19ca773eb68dc0b9bf;
wire [MAX_SUM_WDTH_L-1:0]        Id79c1fa529c3b719ef4534d1c3abc975;
reg  [MAX_SUM_WDTH_L-1:0]        I579480a66a5f6331fb46de13090ce888;
wire [MAX_SUM_WDTH_L-1:0]        I496765810959107754d8f764be715da4;
reg  [MAX_SUM_WDTH_L-1:0]        I38d78b447217271a63f30f78b424e2ae;
wire [MAX_SUM_WDTH_L-1:0]        If1b62fde8c7b6aa858dff5eba22d51a8;
reg  [MAX_SUM_WDTH_L-1:0]        I4c8d7e5474b19a7c63444d0cb6143728;
wire [MAX_SUM_WDTH_L-1:0]        I5a86b5c97d7b531c201169167a720d2b;
reg  [MAX_SUM_WDTH_L-1:0]        Ia4bc4b7414bf31305ec8f63e7eda61e7;
wire [MAX_SUM_WDTH_L-1:0]        I8e0d580b0f875a9373a3d8fb5523183d;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbebe287d56c7d627f3ffcf706575e77;
wire [MAX_SUM_WDTH_L-1:0]        I0a35c9a4f7596b64d8a6e39878fbc83a;
reg  [MAX_SUM_WDTH_L-1:0]        I83867e6ee369fff7e39ef5c8d5398fef;
wire [MAX_SUM_WDTH_L-1:0]        I9eed09a7c7b86123ee154b783cb7e720;
reg  [MAX_SUM_WDTH_L-1:0]        I1d40df7dbf99674f987bd06db714a702;
wire [MAX_SUM_WDTH_L-1:0]        I45efcc842b324efcbf828c6d68f19e84;
reg  [MAX_SUM_WDTH_L-1:0]        I92f42789cb81760ff2973e3a5fe915c3;
wire [MAX_SUM_WDTH_L-1:0]        I4922b2f4381eb54d365a270b32c944c0;
reg  [MAX_SUM_WDTH_L-1:0]        Idbd5f2a25ab05808721cf9c403017565;
wire [MAX_SUM_WDTH_L-1:0]        Ica29fa9ccbb761ae142e6ae7186aa830;
reg  [MAX_SUM_WDTH_L-1:0]        I7ca5f07d6d3c2a045dfd55ae5214dd65;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie1e5ff68116424c122e4763955e243ac;
reg  [MAX_SUM_WDTH_L-1:0]        I7f4e1445c68abbadce23944b99d206f9;
wire [MAX_SUM_WDTH_L-1:0]        I1c817dbc1d0d04ab8d417d31ef477daf;
reg  [MAX_SUM_WDTH_L-1:0]        Id9f28016678e5e2127d9f0aa93e0b534;
wire [MAX_SUM_WDTH_L-1:0]        Id4bf2c50adae02e36a8c7a862a470efb;
reg  [MAX_SUM_WDTH_L-1:0]        I6b939c57a8b7c7c51ab43e1b1df12f6a;
wire [MAX_SUM_WDTH_L-1:0]        I11f3867bc6c57b2f58b19c0ffbbc0827;
reg  [MAX_SUM_WDTH_L-1:0]        Ic5d0df586d56bf4cb322d4c3ad677385;
wire [MAX_SUM_WDTH_L-1:0]        I630f6f37116aab84814e74017b6d3c4c;
reg  [MAX_SUM_WDTH_L-1:0]        I2e287724873cf6761799eaf464ed6302;
wire [MAX_SUM_WDTH_L-1:0]        I3b0edd5d01b89026be06cf00b6eca7c0;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7a10cffe31a53aafa1104b97543280b;
wire [MAX_SUM_WDTH_L-1:0]        Ifad4e44440835f78f56065a3aa29ad3f;
reg  [MAX_SUM_WDTH_L-1:0]        Ieeb089c6a18791a2227c8571913d689a;
wire [MAX_SUM_WDTH_L-1:0]        I93a1ba64d41cef26b742ba06755d77a1;
reg  [MAX_SUM_WDTH_L-1:0]        Ib29b00328971c3cd67209a5ea5b63b0a;
wire [MAX_SUM_WDTH_L-1:0]        Ib2531654b83ce43d8f11a08c36cca4f7;
reg  [MAX_SUM_WDTH_L-1:0]        I517e0868f2bb9a22c287a1f3eeaad2f3;
wire [MAX_SUM_WDTH_L-1:0]        I984fc2e5cd03bcf452fd7eb62be1b5b6;
reg  [MAX_SUM_WDTH_L-1:0]        I2bc9f76469e2a3f9846560ad1975cf54;
wire [MAX_SUM_WDTH_L-1:0]        Ide09ff97f4d7b3049872064c78fd2b14;
reg  [MAX_SUM_WDTH_L-1:0]        I9f089315e435cd69d2929fdd936a8a77;
wire [MAX_SUM_WDTH_L-1:0]        I99c143788bcb9dfcb14e29b1f9117770;
reg  [MAX_SUM_WDTH_L-1:0]        I9b54c9fb4179423c731217286e329930;
wire [MAX_SUM_WDTH_L-1:0]        I4c4a40069ce9f6b40b8a1ec7787cade1;
reg  [MAX_SUM_WDTH_L-1:0]        I82fb41ab743146badfd2e82258afb310;
wire [MAX_SUM_WDTH_L-1:0]        I5a345140c4181b5307ea3c5b79e62b11;
reg  [MAX_SUM_WDTH_L-1:0]        I5619b91de99eead78befdcba1c62411e;
wire [MAX_SUM_WDTH_L-1:0]        Ib9e2a08275b9e2571238c39945aba5d2;
reg  [MAX_SUM_WDTH_L-1:0]        I83dd2047dece99cd841b2e7955819d57;
wire [MAX_SUM_WDTH_L-1:0]        I203718fd22ec9e6e4ac7a9c1973d6837;
reg  [MAX_SUM_WDTH_L-1:0]        I8c927e66ccbf4d19f07af5ef9fbfe3fb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8fa60b209a1ac0d2738e58662612206f;
reg  [MAX_SUM_WDTH_L-1:0]        I0793fa8938acdf65486e5582d01b9e5a;
wire [MAX_SUM_WDTH_L-1:0]        I579c31eb0b51668db2b1edb1f10a372f;
reg  [MAX_SUM_WDTH_L-1:0]        Ied68d7ba0ee9974eb33767e737760b4d;
wire [MAX_SUM_WDTH_L-1:0]        I425545d21b0a9447b41481b5874c6a26;
reg  [MAX_SUM_WDTH_L-1:0]        I95ba37056659b29fd4318a68d85445e8;
wire [MAX_SUM_WDTH_L-1:0]        I2d1670c45bd1cc15172a12175f7fb906;
reg  [MAX_SUM_WDTH_L-1:0]        I08d7051a18f358d08728f1c401c15c47;
wire [MAX_SUM_WDTH_L-1:0]        Ia4c9bac1a64e1a17f7964491d880660e;
reg  [MAX_SUM_WDTH_L-1:0]        I768b6f55827ac49eb6ac2655e9397be1;
wire [MAX_SUM_WDTH_L-1:0]        Ibff15c9092ff0ab60ccfd9528d5477bf;
reg  [MAX_SUM_WDTH_L-1:0]        Ic66f737fe60c55d4c10e5d72b307a061;
wire [MAX_SUM_WDTH_L-1:0]        Iac2e396e7f63a651c52c6aa372419808;
reg  [MAX_SUM_WDTH_L-1:0]        I5653779f15c6c9b0f3b26927c48d6234;
wire [MAX_SUM_WDTH_L-1:0]        Ice856d92219493a98683a6e36f6a81f6;
reg  [MAX_SUM_WDTH_L-1:0]        Iac550729fc437fd67151fab57134ec88;
wire [MAX_SUM_WDTH_L-1:0]        I5e784ab32ea84026fa63ce432c6f604f;
reg  [MAX_SUM_WDTH_L-1:0]        I853b03c5826eedc3c67a2fae7a640212;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I32251a5b768526c3599f145a3eed1949;
reg  [MAX_SUM_WDTH_L-1:0]        If46a6b47c1c52243cc0bc92d1edb594f;
wire [MAX_SUM_WDTH_L-1:0]        I6357b0d86d75dc1018fa50248f3e2deb;
reg  [MAX_SUM_WDTH_L-1:0]        I75b36a9b429cd657afc8151b9613aca6;
wire [MAX_SUM_WDTH_L-1:0]        I8a50948f1b1f5589972c137e91e4eee0;
reg  [MAX_SUM_WDTH_L-1:0]        Ife682dd9f677da4d27294fb61b141948;
wire [MAX_SUM_WDTH_L-1:0]        Icce2cc29f7ad95af1a9605954033fce0;
reg  [MAX_SUM_WDTH_L-1:0]        Ic2b6177a9c586b274b68b25584e6df2c;
wire [MAX_SUM_WDTH_L-1:0]        I276997085c2cbcdac1c886e74bc2e530;
reg  [MAX_SUM_WDTH_L-1:0]        I0d23011c4381496a19cced7bf7960546;
wire [MAX_SUM_WDTH_L-1:0]        I7299d046eb7c80908def7e3ec9665c88;
reg  [MAX_SUM_WDTH_L-1:0]        Ic5992d5eaeafd5dded641a7d9801e763;
wire [MAX_SUM_WDTH_L-1:0]        I8f993e6b8e7313dfb4323ebf4ccdb640;
reg  [MAX_SUM_WDTH_L-1:0]        Ic9e7fe68b9045c6c9eb86185b5f5872e;
wire [MAX_SUM_WDTH_L-1:0]        I2b75fcd754488677526db195256ddc06;
reg  [MAX_SUM_WDTH_L-1:0]        I51ad746720b5e6e09ab50f0283552f1a;
wire [MAX_SUM_WDTH_L-1:0]        Ide04235316ff1098fd97e125d76797c2;
reg  [MAX_SUM_WDTH_L-1:0]        I0c8964888a1315507f5d71959dd24cf0;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I39755c95fddbe19ae343164be78b0fff;
reg  [MAX_SUM_WDTH_L-1:0]        Id4d4f814a0bb3418cbf70c306acf048f;
wire [MAX_SUM_WDTH_L-1:0]        I37d4177c1ea3ac376d3906e49a4a3224;
reg  [MAX_SUM_WDTH_L-1:0]        Ic91bd7b4bd148e526ca21d4a5ba87be9;
wire [MAX_SUM_WDTH_L-1:0]        Ifd04130d9f32af7f7debe20de6b6fa57;
reg  [MAX_SUM_WDTH_L-1:0]        I7959dddc32f0f181b3ba39149afe1016;
wire [MAX_SUM_WDTH_L-1:0]        I7ee40f0225ba9aad10df1dec7a0f25fd;
reg  [MAX_SUM_WDTH_L-1:0]        I087263600b5f38be072a4f1db787aea7;
wire [MAX_SUM_WDTH_L-1:0]        Ic780d894a72f9111937594d50a9ce311;
reg  [MAX_SUM_WDTH_L-1:0]        I78d17a56de5cbe08191ef23b9731c485;
wire [MAX_SUM_WDTH_L-1:0]        I36feeea802ed7e4122a43a71d976b7d2;
reg  [MAX_SUM_WDTH_L-1:0]        I82f713a43596df3b935d6da6f8041dc2;
wire [MAX_SUM_WDTH_L-1:0]        I698319d790c8eb982fb1b113437d93be;
reg  [MAX_SUM_WDTH_L-1:0]        I422987396853a6a39dabb6e7ddbf91fb;
wire [MAX_SUM_WDTH_L-1:0]        I69c4cabd4c61dd816fbc44ae02f3d8ab;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb6556671e104141dd33188ea5fc024d;
wire [MAX_SUM_WDTH_L-1:0]        Id504dcc780b333a51585556c4b58c610;
reg  [MAX_SUM_WDTH_L-1:0]        Ie42ce76076a2a5e887e0112086012da6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0c8aff3de7ee8ede0d8755cb4aebe427;
reg  [MAX_SUM_WDTH_L-1:0]        I4aea430599b9c0702b3bebd5960b5c91;
wire [MAX_SUM_WDTH_L-1:0]        I1898ec6433c0e994bf697eb3b7ae5eb3;
reg  [MAX_SUM_WDTH_L-1:0]        Icbe11a3970136e485eee1bc5053e7273;
wire [MAX_SUM_WDTH_L-1:0]        I41b391dce086564a0de53aa3f82b510a;
reg  [MAX_SUM_WDTH_L-1:0]        I0a7f1ea1719c1f5ff104445a4130a5a8;
wire [MAX_SUM_WDTH_L-1:0]        I90c35450751e2a9607e95ebe3115c51c;
reg  [MAX_SUM_WDTH_L-1:0]        I1802d759f26dd919bc315bfd4156238d;
wire [MAX_SUM_WDTH_L-1:0]        I02be13e15f91f4957ba7086ee96c1ca7;
reg  [MAX_SUM_WDTH_L-1:0]        I2148493e253783fad70f4f2807b83008;
wire [MAX_SUM_WDTH_L-1:0]        I02cc4624a6245c0c54b079dfe50420d4;
reg  [MAX_SUM_WDTH_L-1:0]        I39e7f78d33aa7f50264908d2efe23634;
wire [MAX_SUM_WDTH_L-1:0]        Ib0942c283a523d31d5d11a51f01fa016;
reg  [MAX_SUM_WDTH_L-1:0]        I844be5874def16af98de935019f35fe8;
wire [MAX_SUM_WDTH_L-1:0]        I93ad63d6294ac100b7027b8190f15387;
reg  [MAX_SUM_WDTH_L-1:0]        Iee5172ba70a6e368b4903f9ff1d93471;
wire [MAX_SUM_WDTH_L-1:0]        I8b92187b5833150d05b4b09f74441a20;
reg  [MAX_SUM_WDTH_L-1:0]        I1f34b473283291e0970879465c005e2f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I02846f27754a2fbc493cc1d0848b9090;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1e0b5120737a7f4bf845618ccd22239;
wire [MAX_SUM_WDTH_L-1:0]        Iea2573c99c098c5fe2ee97a9c1aae44d;
reg  [MAX_SUM_WDTH_L-1:0]        I8abec3020ee5358f8768e5595e9992b4;
wire [MAX_SUM_WDTH_L-1:0]        I8c250d6e46e2d8a7f2f77035526c1f8e;
reg  [MAX_SUM_WDTH_L-1:0]        I6fe683073211a484cb6e3c416b365d9f;
wire [MAX_SUM_WDTH_L-1:0]        Ic968e5570985a076b609845c9968110c;
reg  [MAX_SUM_WDTH_L-1:0]        Id7d764da58ade36853e8a45b5ee19dc3;
wire [MAX_SUM_WDTH_L-1:0]        Iccd14e61a9147bf5aefe4a196485ef03;
reg  [MAX_SUM_WDTH_L-1:0]        I3cee2fdf353643deac7d6bca20c8fb52;
wire [MAX_SUM_WDTH_L-1:0]        I4e09b4d678ce7239bad645b57535df20;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9b8f8f0434fe3783c3d8f68fef30e50;
wire [MAX_SUM_WDTH_L-1:0]        I6bdb1743d21a19cf2ce13b056271d1b0;
reg  [MAX_SUM_WDTH_L-1:0]        I68cba8ad7742cbb34d0b1fb16be4a58a;
wire [MAX_SUM_WDTH_L-1:0]        I6259bbd85d21c216632a71648eddae35;
reg  [MAX_SUM_WDTH_L-1:0]        Idcea56657d40e0fdf9a1c2d920938fd6;
wire [MAX_SUM_WDTH_L-1:0]        I8a654b2420f09bd4b14bc5f5faa7d40d;
reg  [MAX_SUM_WDTH_L-1:0]        Ic549ffab8f0ce161a177faa2ffd1326d;
wire [MAX_SUM_WDTH_L-1:0]        I50d163f8fe5bbb86e3843bea768f049e;
reg  [MAX_SUM_WDTH_L-1:0]        I4d463d500f93f74b2724972ec1d62439;
wire [MAX_SUM_WDTH_L-1:0]        Ic3e2b4869f7ac3d189713dcc40a1fb30;
reg  [MAX_SUM_WDTH_L-1:0]        Iba2f362e263953331649c726afa9c481;
wire [MAX_SUM_WDTH_L-1:0]        I3d8f79c5f5af5112dc5f7fdfaf0a2434;
reg  [MAX_SUM_WDTH_L-1:0]        I6a053d931fb030e03d4882856d3bda75;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0544d6bafecefee496a6227c698a4d1a;
reg  [MAX_SUM_WDTH_L-1:0]        I27ede93004e0c240efaa56cc8c570910;
wire [MAX_SUM_WDTH_L-1:0]        I6672e8613ad03882a4b7f4141a56d535;
reg  [MAX_SUM_WDTH_L-1:0]        I61a11c1711ca10eefea3438722b40bff;
wire [MAX_SUM_WDTH_L-1:0]        I1542f0db2447a8b733077daebe1d2321;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7924c88692cfddf24fb1eff66eacb7e;
wire [MAX_SUM_WDTH_L-1:0]        I3038115e5ee2b90df4a7ad7e25d5337d;
reg  [MAX_SUM_WDTH_L-1:0]        Ibcfd01e622f7f5a5156dd9b335b4e5e0;
wire [MAX_SUM_WDTH_L-1:0]        I758ce2910b56968ca8ebc74c19f2cb47;
reg  [MAX_SUM_WDTH_L-1:0]        I7f6f418ea51b4298da8758bda3f6a21b;
wire [MAX_SUM_WDTH_L-1:0]        Ifd3191045c45b2f46fbbb63b1766e9fb;
reg  [MAX_SUM_WDTH_L-1:0]        I7185da8937449e23abdd0f39a4b3ed7d;
wire [MAX_SUM_WDTH_L-1:0]        I5a15f4c8b810f7234d421967f4d926c6;
reg  [MAX_SUM_WDTH_L-1:0]        Idc3e3ffa31d9b76c7cf9358a5b2e65d7;
wire [MAX_SUM_WDTH_L-1:0]        I6f82614fc25bf322e359b929caa86025;
reg  [MAX_SUM_WDTH_L-1:0]        I31fe8c887c4aff7c69336676cd31aaa1;
wire [MAX_SUM_WDTH_L-1:0]        I4dcffaa8c903a955a4c4b5197cd2d728;
reg  [MAX_SUM_WDTH_L-1:0]        I59684d5fe6bbb4b54ac097bd25fceef5;
wire [MAX_SUM_WDTH_L-1:0]        I71dbc37567c4c703f28c39b97c44d1dc;
reg  [MAX_SUM_WDTH_L-1:0]        I86a7cd69148f9590ce91d0aa270d6c54;
wire [MAX_SUM_WDTH_L-1:0]        I224678d6b3b2a1ed8f2368d7035134d4;
reg  [MAX_SUM_WDTH_L-1:0]        Iabce1ccdd968980f622f0e137b159d11;
wire [MAX_SUM_WDTH_L-1:0]        I6942bdfb9c73af7b24e91f3cc2c40443;
reg  [MAX_SUM_WDTH_L-1:0]        Iff02977d7b4c733cca1794246f630931;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8eae50dae3f5eadae891e7875180bd47;
reg  [MAX_SUM_WDTH_L-1:0]        I9026c904e5ead7ff2994c4f781d61466;
wire [MAX_SUM_WDTH_L-1:0]        I5ab8c899cb9e33273d3e5758757dbdfd;
reg  [MAX_SUM_WDTH_L-1:0]        I99d7489ba87c629c6dd9702a9bbfd3c8;
wire [MAX_SUM_WDTH_L-1:0]        I23890d77a1b1c3fea977146599cee178;
reg  [MAX_SUM_WDTH_L-1:0]        Ifaf191e0d00ba6da7019c2efcf08e1d9;
wire [MAX_SUM_WDTH_L-1:0]        Ib311a6a7fc40711d6920e3c43b31c5c2;
reg  [MAX_SUM_WDTH_L-1:0]        I4c295991fb08c90862a2f3ba6489000a;
wire [MAX_SUM_WDTH_L-1:0]        Ifc3cc051690f3d687caa05e26dde6d93;
reg  [MAX_SUM_WDTH_L-1:0]        Iee61d179da125934298400256788cbb8;
wire [MAX_SUM_WDTH_L-1:0]        Ida60773a931859ee7e5e2db24b9bb72c;
reg  [MAX_SUM_WDTH_L-1:0]        If87c84440426fb24070372dc1d4bf315;
wire [MAX_SUM_WDTH_L-1:0]        Id5e39679bbe2407407a53366e77aed13;
reg  [MAX_SUM_WDTH_L-1:0]        Ib9259a807b31c1b7a528d336bfc403ee;
wire [MAX_SUM_WDTH_L-1:0]        Ie3eab29a9004627e296a198708459545;
reg  [MAX_SUM_WDTH_L-1:0]        I411c4d909b2a571e685cd703245516d7;
wire [MAX_SUM_WDTH_L-1:0]        I86c0872f8ce743bb3fa7b3fca2dea33b;
reg  [MAX_SUM_WDTH_L-1:0]        If8425453cca8fc8623cb85375c4b8a1d;
wire [MAX_SUM_WDTH_L-1:0]        Id1aa022173e0fa45a3f26b4d31e113a3;
reg  [MAX_SUM_WDTH_L-1:0]        I654b497f62df75fa283127b5de29b1ad;
wire [MAX_SUM_WDTH_L-1:0]        I0bfd4314a81f9f0930e549a09ef4c68f;
reg  [MAX_SUM_WDTH_L-1:0]        I2768519342f7b8a1ee40c1d5ac502b66;
wire [MAX_SUM_WDTH_L-1:0]        I2e90a66f2eedee35927bcb8c5ff26fbe;
reg  [MAX_SUM_WDTH_L-1:0]        I8e354c1c5ba44fe5430887248ce0c43b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I9d6828434155b5672b44a1172ae9b6eb;
reg  [MAX_SUM_WDTH_L-1:0]        I8970d8a8aea29913e8696c14c153d16e;
wire [MAX_SUM_WDTH_L-1:0]        I0483abcf888b35d85e8a62c901b6021b;
reg  [MAX_SUM_WDTH_L-1:0]        I3555c6e2fd480a6be11549bf95a9b0b1;
wire [MAX_SUM_WDTH_L-1:0]        I8f6514c2e33675cd94350a1e1b0b5f80;
reg  [MAX_SUM_WDTH_L-1:0]        I8d5600a352e8ba4756f917f912fda6dd;
wire [MAX_SUM_WDTH_L-1:0]        I23d3830f616b3be90cd63e45b606fc2e;
reg  [MAX_SUM_WDTH_L-1:0]        I7e99d73c95e7ae5c3fe07a3c60ef52eb;
wire [MAX_SUM_WDTH_L-1:0]        I106ef13f4b977bc5b978b5977cc06eb7;
reg  [MAX_SUM_WDTH_L-1:0]        I831633aebe5c6a52b98d630205376f3a;
wire [MAX_SUM_WDTH_L-1:0]        I3fdcbddec1b193cc85d20d4796aef72b;
reg  [MAX_SUM_WDTH_L-1:0]        I82e35482de74223be0d2558334ac2dfb;
wire [MAX_SUM_WDTH_L-1:0]        I3956ec3a4f9d8ea94a760b5c6388f2b0;
reg  [MAX_SUM_WDTH_L-1:0]        Iae2a6f9649ef1bb193e4f0ab5ecbc3e3;
wire [MAX_SUM_WDTH_L-1:0]        I5541cea9c0da962da2b7d9154c66de98;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8eca65d791ad2f6e8f4ed244f22ae3d;
wire [MAX_SUM_WDTH_L-1:0]        I0c1edbaa3c2f47d66034fccd799b5387;
reg  [MAX_SUM_WDTH_L-1:0]        Ic24146b01094df9b9ccd455a791f239d;
wire [MAX_SUM_WDTH_L-1:0]        Ia6eb0c9c2e6c3a440defef2c3879de88;
reg  [MAX_SUM_WDTH_L-1:0]        I1c9031fd54ff9417d44c9fb17dc1fc63;
wire [MAX_SUM_WDTH_L-1:0]        Ifcef7363a6ecbb3b3248cb65bb6b0d17;
reg  [MAX_SUM_WDTH_L-1:0]        Idefa20487bc5ba6daff03e6b327d76c6;
wire [MAX_SUM_WDTH_L-1:0]        I5e36ed7643bf47aef14bd47a835e1a01;
reg  [MAX_SUM_WDTH_L-1:0]        I6f984fd9ea27b40ab3afeac8afd29ade;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Idc662c9332f4a6cafe820ad2bc0d16e1;
reg  [MAX_SUM_WDTH_L-1:0]        I0be92debced4961df5f461fe81e80bf1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Id51e465dc2adba5eedf6ad37d0a25aa3;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7bdaba4c6601b7146498aea6c9a3e07;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If0d4550f2f3884c49d1cf5a40251cd58;
reg  [MAX_SUM_WDTH_L-1:0]        Id450c0a1cabe087be051fbf4158e6016;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3af1a3cc1733db0dc42ab6214351aa99;
reg  [MAX_SUM_WDTH_L-1:0]        I656d0d69f6e243746b87ad67764dbc3d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I022b7b4693a7e7b654b8bd85a94f0d9c;
reg  [MAX_SUM_WDTH_L-1:0]        Iab9d870dc1ad159bbaecb20a9b72f005;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5bd1d6563b4acb8dc10d348ec0a2346a;
reg  [MAX_SUM_WDTH_L-1:0]        Id53b60854f19e095c38f2c255dc57f29;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I17bbbddc2ace71bcd660f93fdf5e32a4;
reg  [MAX_SUM_WDTH_L-1:0]        If9ba44a2e4a8f0b61692fc69ebeb82bd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I4eb0952c6dd9719774c57b76d3cbe87a;
reg  [MAX_SUM_WDTH_L-1:0]        Ief95e8620a1c8ddfd6df673a3a223bd8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I6fb63afabfeb4cc43c164e04d35a6c76;
reg  [MAX_SUM_WDTH_L-1:0]        I61519bc0aa02ed461dbb91851d0ae19e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I91ba6681ef5a1092784cd98b48dc420e;
reg  [MAX_SUM_WDTH_L-1:0]        Ie0c11d584811174a66ca221baf87c36b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I6eda15abfd6c1f377d25d70e35373596;
reg  [MAX_SUM_WDTH_L-1:0]        If10f4f45ff0fd17541735934ad20f187;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Idf9a54c3bd991a031e09982424a8054b;
reg  [MAX_SUM_WDTH_L-1:0]        I445919f07a6fa8654211301a9a6126bd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5d7b50b4839c16d1c7010ef2c8c535c2;
reg  [MAX_SUM_WDTH_L-1:0]        I64102b82893352549abd2e2132b19476;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I821836ca9d1bcb5e0d12c348bb323c9a;
reg  [MAX_SUM_WDTH_L-1:0]        I1fc1933fe891ac26f35a42a1b242d919;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I31f94bb809811efebb378517c2138b7f;
reg  [MAX_SUM_WDTH_L-1:0]        I84dfba8bcf8ad3b85f9472fd60d607b5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3f203b62c645fd01c54ed43399b390e5;
reg  [MAX_SUM_WDTH_L-1:0]        I4302fccefe5ee13161f9ad49f9ddf43c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic01c569fbe524a2fe3626e4d22414e62;
reg  [MAX_SUM_WDTH_L-1:0]        I59d7153724d3b3805af799692fbe245a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5a30e151cf8a2259d8cde3fa76389e78;
reg  [MAX_SUM_WDTH_L-1:0]        Id1650d0e39be078027493f58e9bbcbdd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic5340f7fa98175b85f475a03156a04a6;
reg  [MAX_SUM_WDTH_L-1:0]        If40ad4aca8dbb3bf7dde8c2ff2e5b8f2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0b25b22531e117125c9dc82b1fb69166;
reg  [MAX_SUM_WDTH_L-1:0]        Ie49f173549396caeab1d13da36e37c65;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic0c22023bce6b4e011b52acb0ac89944;
reg  [MAX_SUM_WDTH_L-1:0]        I3002a0e0cdf8e79bc7186a876410d106;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I7f474f465227aa0e2aaa3986574ed756;
reg  [MAX_SUM_WDTH_L-1:0]        I2b50fa03f584d10e9af3be085a02a12c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8869bb7415e726932972a16630d4090a;
reg  [MAX_SUM_WDTH_L-1:0]        If473d172a7bff5aeae99245bbb72978d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic1afbad56abd1a486de1d72dc835ea03;
reg  [MAX_SUM_WDTH_L-1:0]        Ib89f7b5625995290a64bcfb143d978ca;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0cc174ebcf049214088dd4a7dad9ebf0;
reg  [MAX_SUM_WDTH_L-1:0]        Iebe0c9b4a87d58a1c55e2ee6b01603c4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If9a4389e51bb56f222cf06e66dcefbbb;
reg  [MAX_SUM_WDTH_L-1:0]        I104411bb641d2445c7e1385a809bb682;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iff6098f0561da4ad6ee64dbcbf7a8b94;
reg  [MAX_SUM_WDTH_L-1:0]        I47dd28b4ae4f7151aff5bb271e35b716;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I26a679e345a21470331cd4fb2512dea0;
reg  [MAX_SUM_WDTH_L-1:0]        I3a27d5573b748df459b90a5a347f9d09;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iec11498f4ab0492570a3454760ed5679;
reg  [MAX_SUM_WDTH_L-1:0]        I2dbef85d2b2b95af39c3a98c4e143253;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I78154c0ca0236b79bb58bc2942b0f51b;
reg  [MAX_SUM_WDTH_L-1:0]        I510d39830ae7b0a857ac11baa7c144d3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3a2c3112d5ba223b037baab170e9da79;
reg  [MAX_SUM_WDTH_L-1:0]        I2751a94a66ea4cb44c512df4c509937f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ia56b6d58ede63ec2b56533f0804b16df;
reg  [MAX_SUM_WDTH_L-1:0]        Ic9a003bfb70ac2da6c229fcad09246d4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If8bafc8e64df4d25c725f8c577e6db43;
reg  [MAX_SUM_WDTH_L-1:0]        I34ed986182a3311a8cb005b3dccc224b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie7452b79bbda04bebf83147d7f2ddcec;
reg  [MAX_SUM_WDTH_L-1:0]        Ic79281755397f6099ff30c5d07d7e6de;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I29a84f35944a4e286c267c60d9899c62;
reg  [MAX_SUM_WDTH_L-1:0]        I8d6559ccc33cbc663584923a55b928b5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iae0a8cc0afb8366a7c9df146c0d08eb0;
reg  [MAX_SUM_WDTH_L-1:0]        I4f0a4c241844e390318f11899a0f2c5a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I39d0497d0550115c6a2c08676c451845;
reg  [MAX_SUM_WDTH_L-1:0]        I45fffa266ce3838f82d755b59216a4d6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ia96a79462a86a7ed9e337df66d99bf92;
reg  [MAX_SUM_WDTH_L-1:0]        I8f0e65f5db47d5460d4ec2172807a3e1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8ef19b31ec6d7e52e78b0c673f23ce12;
reg  [MAX_SUM_WDTH_L-1:0]        I34127c0d1af2438e13b6f4709ece80ba;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8081b1486e6def0f6ae514513c7ef4de;
reg  [MAX_SUM_WDTH_L-1:0]        I3a67de0e76bbf29d8c77c21865abda2f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iee5a68c2d52ef1cdd3f19b0a912603cf;
reg  [MAX_SUM_WDTH_L-1:0]        Ic64e64aeb754249b868e14311ea19759;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I4b5525780a9259b57497235bd0bc69a4;
reg  [MAX_SUM_WDTH_L-1:0]        Ic4aa0dc9014c8445f8d9a7723d7263f5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ibd65f08dbbf43d438c3a985c7b17f2e3;
reg  [MAX_SUM_WDTH_L-1:0]        I47b988d017580bdfe8f443904b1f3aac;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ifaa5785a3e04cd1e3be505042347fe26;
reg  [MAX_SUM_WDTH_L-1:0]        Ica9ff13e8c3850be6c70b0b06c1d9fbf;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If0cb8cd465ff1f65de99688abd92aef2;
reg  [MAX_SUM_WDTH_L-1:0]        If2efeb489911f295dd7722cb22ea521d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I10ff180c115b9372f9b4b12df313372f;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa16dffcc01e41e6ff17e92bdefe3df5;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I64f177202fe847d13a8a12bd80a45946;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8857b9841fbd795a4192976ef7ecc25;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5df97e26d5887da447669b8d932fbdd9;
reg  [MAX_SUM_WDTH_L-1:0]        If12aef69eea28052aa3bdb6ac31af205;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ibdc07eb6a0a66e1393cb2dbd9ac77c72;
reg  [MAX_SUM_WDTH_L-1:0]        I0b3c6162ae2b9221738a18a29489887f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3d353247a021629a4dd38a784eba5c1e;
reg  [MAX_SUM_WDTH_L-1:0]        I08211bba29e87faf4079152bcc973e7d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I20d77ee5328ef46daa4a54c0ae98d31a;
reg  [MAX_SUM_WDTH_L-1:0]        Ibff3da265f1c3f21548f5b019e1a9dc1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8284c3a4664f99934170474b8e0e73bd;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9fa1762d7844b0d781afdfb0771cea9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iaeb44f2b4b78055f103df8070110b5b3;
reg  [MAX_SUM_WDTH_L-1:0]        Ia677d504b9f7fc2698c0345f236428ba;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic8242c1f7d2f582c63c3cea63d929945;
reg  [MAX_SUM_WDTH_L-1:0]        Idebce29121c0481df83d755b60ff632c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib9dfa491b9914f9ac567ae8681a2cd6c;
reg  [MAX_SUM_WDTH_L-1:0]        Iad2c780a6386674d50cca54d8c4ebd86;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I029b75f94f58485022bf37590df82900;
reg  [MAX_SUM_WDTH_L-1:0]        If1d7944e7c4828ddb91ffea28609cbc7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I1cc49a7f6f5c1ecd775d2734c3321364;
reg  [MAX_SUM_WDTH_L-1:0]        I843a68ceb0adab829091f31d0de56eb6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I596867e7be52dbcabd95cdd2600396a0;
reg  [MAX_SUM_WDTH_L-1:0]        I59701b9eb54dda2744a79cebe7d73f3b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iec0928bbbc2730b835fb20d75a988a7a;
reg  [MAX_SUM_WDTH_L-1:0]        If63cf5e8f47e4e51176401f0d954ea23;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iabaf04fabdf2dc5fe29d1eae22b23f7e;
reg  [MAX_SUM_WDTH_L-1:0]        Id09454844b525697de3e3727d89551e4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I678858a018330bbc4ddb8fe46ff09f49;
reg  [MAX_SUM_WDTH_L-1:0]        I6d1b2ce4368945b56eee7814638471cc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I453a3e7067a9421392ad43b673f203e1;
reg  [MAX_SUM_WDTH_L-1:0]        I6079945faa57335b1c902ccf7f960a70;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I1a3dcf633defa34860b0db5fed0d710d;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7752906ac55cf51f3e96e8c0046f1aa;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Id4ba510039040276d71a221b3468977e;
reg  [MAX_SUM_WDTH_L-1:0]        I2d7d4135a94f5df949283c043228791f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I7b9204a45b89e3800944d49a811a930f;
reg  [MAX_SUM_WDTH_L-1:0]        I99c75e3d26c5d01f6ae9abcd05407d8c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ia9d671775a9c5d0c1c0886abc70c5100;
reg  [MAX_SUM_WDTH_L-1:0]        I81e6f97621dbfb2fed6fc236005a2b19;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ief6f4ea0ada586ed46ce19d0761edf66;
reg  [MAX_SUM_WDTH_L-1:0]        Ieac60532dcfc916a65054e35cf31d6d2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I02e35fcbb30d8951f129525146af7f9d;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7eb83ba73e0dc17f69c357b6ca555bf;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ia55f4e6ae1e56d5aee09414ba7617fc5;
reg  [MAX_SUM_WDTH_L-1:0]        I5139d8a7a099e3c619c60647c15b7420;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I4f077fadda92556acba301e0990a8d47;
reg  [MAX_SUM_WDTH_L-1:0]        I6ccd2e11ebd5b2de80b120e20650a602;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8fc930fd14a7605288eea0d3f7561930;
reg  [MAX_SUM_WDTH_L-1:0]        Ie669cebe5fe39e1a841f8dd3c1f6bc57;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I29eceabd1f5dfb4cc3028ec248645616;
reg  [MAX_SUM_WDTH_L-1:0]        If32acb9fc212c4af34099acf6df2bc5a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If55674824a5a3574ffb2f7da75e2f2d3;
reg  [MAX_SUM_WDTH_L-1:0]        I075ce236a181bf925c8ccce91d9bc8cd;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I12b13bd78932e54099144478a82ae60d;
reg  [MAX_SUM_WDTH_L-1:0]        I541d4e422b999a0dfca44d275178e1d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I09a98ded5754d5439ec3a384635d63c8;
reg  [MAX_SUM_WDTH_L-1:0]        I3e02657f3d9f79338cd083ed024bf96c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I802fd7e7eb9c1b2fd917b1eb657e71b9;
reg  [MAX_SUM_WDTH_L-1:0]        Ia5e5537405ab8edcc7cd43c86837d43d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I264cc4045cfc24b211d08488ad2eb105;
reg  [MAX_SUM_WDTH_L-1:0]        I07ff388e3b6c7288f0f6c35a345023fe;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iaa96c298cadeb650acccbd3e548cf281;
reg  [MAX_SUM_WDTH_L-1:0]        I56cb3b3e193ca5068734417fd0ec4e02;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I463f424b1cc557868a77721849b635a3;
reg  [MAX_SUM_WDTH_L-1:0]        I5bbf1765d8f81581d0cf31c0bc755fb3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5fe371b91ca52980957e017a6dbd2308;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa1643095e518846cdede4d5a90dff84;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ia301618cac1f678b17595d3e87a85068;
reg  [MAX_SUM_WDTH_L-1:0]        Iee6e12f4717a3279dd31b874eabae69e;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0ce7b89ce37757be43c464793608e6da;
reg  [MAX_SUM_WDTH_L-1:0]        Ic52a9edbbc5283844d2514ea142ca6e2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8abcaf2ec878673e81c94be11046e97e;
reg  [MAX_SUM_WDTH_L-1:0]        Ice3e978c8da2a7de5b28542a5589f0a2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie394af0713a3eb30d9d5c0cb38414b90;
reg  [MAX_SUM_WDTH_L-1:0]        I336a425aed221c85ca80b9a97d21d6b1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Idc8ef4846c1f33c0510b0d4c1b027c81;
reg  [MAX_SUM_WDTH_L-1:0]        Ie477c0f3b77bb299ba8b1a410d211ef7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib0e1198c7bb8c8bd611fd9afed1bf0ac;
reg  [MAX_SUM_WDTH_L-1:0]        Ie62920d089ae762603cd33fbf97d92bb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib2224de3f3f6f644c9e2278ca159eb90;
reg  [MAX_SUM_WDTH_L-1:0]        I2ca952e4e676537fd5a8fc71ecfa10e9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iad987f88aaf1b32bee71e96904d0c51f;
reg  [MAX_SUM_WDTH_L-1:0]        Iefd31e7ff3c829c88f60bc89d70afcf7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0831e757dd5e5868bb023dd9004fb68a;
reg  [MAX_SUM_WDTH_L-1:0]        Iafa987a413fd8fcacfe872bc0f5bc2d6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I64b4330df88134dffb32e0dfd8d4ab36;
reg  [MAX_SUM_WDTH_L-1:0]        I305c1ea420d666f258e38c5a65847367;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5066c1fb5193c037de084c7463947151;
reg  [MAX_SUM_WDTH_L-1:0]        I9f040c4088bfab72d74e5332e9710d1a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I76c57762b38b9546bc862bccfde73a81;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2f41f9778324a06daeb185c736516a4;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I4720972ec687864e66b86780a4a03e47;
reg  [MAX_SUM_WDTH_L-1:0]        Id9778ba5fbdbed4d33a092da6b68c414;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib0da91fdb282ea40f13881671d9736b3;
reg  [MAX_SUM_WDTH_L-1:0]        I27c2c79d0d719c71c8e28218d1174a13;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ifac345df39972bcecf0cf454e30c0cea;
reg  [MAX_SUM_WDTH_L-1:0]        I2a9d6a774769b12ae20bc0cee0c36f5c;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I47ee2c7239716a56029d9d7dd2efeec2;
reg  [MAX_SUM_WDTH_L-1:0]        I2c567b75f1399c069b95284f4c36b6d1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I02398b40df5e80a6818d7f7c20896897;
reg  [MAX_SUM_WDTH_L-1:0]        If3d3eb609abfd6e315eec803d2e94490;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5943d30c92a0938ea3933ba61819ce91;
reg  [MAX_SUM_WDTH_L-1:0]        I9c58aea7ce986b1d28f5808b347c015d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iab0a2d1699d14959918590a17d221dac;
reg  [MAX_SUM_WDTH_L-1:0]        Id139c7a783196941100003b6cb0cd1e7;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        If30544b94b0d43b30a8e4a1a6f67e461;
reg  [MAX_SUM_WDTH_L-1:0]        I524d7614b01460778da3ce98f6aaa3d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I4d6cdcb3b63c51d9dd8b915eb0645255;
reg  [MAX_SUM_WDTH_L-1:0]        I8acda65f116d5c91cbe2662ac282aa31;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Id147fa768121368db44934717c87f635;
reg  [MAX_SUM_WDTH_L-1:0]        If67dbe22f8d22b3430215fb0deae8204;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I7f67e05ed60a537f26feebbbe643a67c;
reg  [MAX_SUM_WDTH_L-1:0]        I9a35cd7512787263abedd6d9913cf507;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I376c401480a2d8e6131123a91e6fa1cc;
reg  [MAX_SUM_WDTH_L-1:0]        If9cca23469c5e6001650f1f8b1360ae8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic33856f32df0ab980accff5678cceebb;
reg  [MAX_SUM_WDTH_L-1:0]        Icc2606ae8f9a3b425225ae7339112b9d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I97e41b86305179e201cce4d69c2ffa21;
reg  [MAX_SUM_WDTH_L-1:0]        I34aa1802d24e074ae54563898929abfa;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iecaf532a526a0f689b65a6dd749d66cf;
reg  [MAX_SUM_WDTH_L-1:0]        Icb85b3464dc40e8504c53c377e889c45;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ia54ab64aa44544f38180c57e0864e071;
reg  [MAX_SUM_WDTH_L-1:0]        Ie595a7d10b5ac84c0301fb55bebd3680;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8ed5770ee3c9a504d934506743f6b427;
reg  [MAX_SUM_WDTH_L-1:0]        I9c217a672cabc05efbdff218637123ba;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I7541c0e729546e0e13e98f4658b95a1d;
reg  [MAX_SUM_WDTH_L-1:0]        If20f3780b4af857ffe8083056085517a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Id861f8b6cc578cfb1d83d065ae78dedb;
reg  [MAX_SUM_WDTH_L-1:0]        Ic2e275bfa8ab3d2002d2aa374ac9bfe2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I6fd4a37bc3b6eb96e6b7e814b203ed21;
reg  [MAX_SUM_WDTH_L-1:0]        Iac5798fd9915b6778700da6a14f6a381;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie31fceaf1518af42616d21bd8247577a;
reg  [MAX_SUM_WDTH_L-1:0]        Ide3204bf317fdfb993410d338085b174;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I89ecfbed8d99ec79402dd5f3f1e64100;
reg  [MAX_SUM_WDTH_L-1:0]        Ic3a95140fc1029efa17a6557bc977719;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iddde66a99ea9a0caa45b06e168194488;
reg  [MAX_SUM_WDTH_L-1:0]        I647d3a46bb2c7ed0f1ec08760b3858be;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib645c9e05a543ca3e8ce0994e56aac70;
reg  [MAX_SUM_WDTH_L-1:0]        I4816747af9d9fc8dc85fd831336ec710;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I29fedc646a3ba823d0dcbb3ecb9b9ad6;
reg  [MAX_SUM_WDTH_L-1:0]        I1f66c026a5437320bd1f4df2ff71663d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie89f6128d6d68c146ffcecb551618321;
reg  [MAX_SUM_WDTH_L-1:0]        If347c58c328193f420286ea27a4afa20;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3388d6fa5159183888944f2951de9361;
reg  [MAX_SUM_WDTH_L-1:0]        I7a126c8304be920f2a920315dc61ba7f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3575e2d60ee8b0b71c67d53b496e2775;
reg  [MAX_SUM_WDTH_L-1:0]        I237327d6a74df1fb05537dc3691ebf11;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I52cf4fceee16d75ea59dbb574ea7c7b0;
reg  [MAX_SUM_WDTH_L-1:0]        I64a3e8bb4c87b066806d33a5306a2c53;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I59cfcae849791453127d60b213ff7355;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbca6ec39234473fb517447a8beacafc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic218ffc97e5e89851d44554326aa5bae;
reg  [MAX_SUM_WDTH_L-1:0]        I78327356176a16fc996188b83b058cbc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I6886b93a81c52c7f93b506404b6a4252;
reg  [MAX_SUM_WDTH_L-1:0]        Ifec496c87a7a2474855067305ac8cba3;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Id9c9ac52a48ef3207581bd31c0593b22;
reg  [MAX_SUM_WDTH_L-1:0]        I41584165a62caaa37ddebbf79bb8b617;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ib3c08e618350ef723607b4ee58bb4dd1;
reg  [MAX_SUM_WDTH_L-1:0]        Idf0916d6b025aad6eccb98ada5ba3aca;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I2481f5b76264c857df96942bdaa941ca;
reg  [MAX_SUM_WDTH_L-1:0]        I00ef133d5a53f8f99f35b50327e5272b;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I3a5aa34be4c3adccf4aad2772c38e972;
reg  [MAX_SUM_WDTH_L-1:0]        I6f0e302d38d75982d0761e306ce9f146;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I95b6796cf442383290a32bad614664e8;
reg  [MAX_SUM_WDTH_L-1:0]        I127eed5de00e10a020717e796de76c7d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie45ac55c4add6c3390924c54d2e8d65e;
reg  [MAX_SUM_WDTH_L-1:0]        If9aad73aefb1b225f35e8c813b85fe87;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I0935498f4dd90c1fed52d2246ebe326b;
reg  [MAX_SUM_WDTH_L-1:0]        I00a89ac37676521a081a21b1ec1a0798;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Iac314ba0cecbd52f3992323dbce81856;
reg  [MAX_SUM_WDTH_L-1:0]        I06f3a34f2b1770ef82ddc2a732b3d4fb;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I2f8a71c2c9078e2581087c7662c961f4;
reg  [MAX_SUM_WDTH_L-1:0]        I4744d64a746f16004e3bedaaa41465f1;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I38c53b94ea9a59a52cdcfe6681491da8;
reg  [MAX_SUM_WDTH_L-1:0]        Ifae0cc6cc1c65d24bbe84c4ba938e2ea;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I5c2c6a0ca07e820e699062299b7064e3;
reg  [MAX_SUM_WDTH_L-1:0]        I1223c21129382d41e4f38ef4bbe60c2f;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ia962052eea10222a1c16ce5800e1c063;
reg  [MAX_SUM_WDTH_L-1:0]        I14e36e16df00adcd7dc1973d3852d2d9;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I33ecd2de3fc7f48821e40313b5dc2093;
reg  [MAX_SUM_WDTH_L-1:0]        I0d05ae27b53fb6939e4c2f862a8d20b2;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie4d5fc4a5bf560bf75561f7f6baa761e;
reg  [MAX_SUM_WDTH_L-1:0]        I97a6fcc08929c3b7d15e36d7706ed13d;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I57de351c4dcc2f9c6bacdf1f39961723;
reg  [MAX_SUM_WDTH_L-1:0]        I1f04e86bf27596718836d0a09adbe120;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ibf1a5a90d4a7922c4bd6273c9a3f1701;
reg  [MAX_SUM_WDTH_L-1:0]        Ie40873cfd6d10a61a94a761becf588a8;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I8a9e51ef30c6434e44fe23412d20425a;
reg  [MAX_SUM_WDTH_L-1:0]        I61960ed74fee948cc12bd1fd8384559a;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I796d4045b29e6c1100dfed4a78dbb912;
reg  [MAX_SUM_WDTH_L-1:0]        I8533a3ec4be4c49166184c94761eaebc;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I32551e388a1ee2ecc7d7da3a4646177e;
reg  [MAX_SUM_WDTH_L-1:0]        I00be319b5bdb85ffaf3bb0eca0b348b6;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I6c266cffd4d2836af16d4d81bbd11250;
reg  [MAX_SUM_WDTH_L-1:0]        Ie889c916b5af185b52ff5e2e3cc23045;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I9feff48bffd8e1f9eee0a587b4b026d5;
reg  [MAX_SUM_WDTH_L-1:0]        I89697be6dcb2e7f972db498c1b1dea71;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I6c540a2cc92ae1fc269a3a395504a08d;
reg  [MAX_SUM_WDTH_L-1:0]        If13dfbfff7cd8e197bb44006a3db73bf;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I683c93eb9205a2272d286e4ad0e998fe;
reg  [MAX_SUM_WDTH_L-1:0]        I87ed6c3e172c7a06bf6aefe7bf718d70;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ic92cbaba339661a83c8bbd3f8377c105;
reg  [MAX_SUM_WDTH_L-1:0]        I0db87adc849839fab3a4c9884d5a4882;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I81850f6963cf07be478907b167cf9206;
reg  [MAX_SUM_WDTH_L-1:0]        I535e01a6c35fd7b455e4b79b1d4bb414;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I6d94790ac6714bb8c62a82bb06960fbf;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2d1c752cc4b405adb97a815e90a7b96;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        Ie19542cb6dc9324368b1ea75a5d5c274;
reg  [MAX_SUM_WDTH_L-1:0]        I9ac12eb3878f6fc7dc428fe5e7f35d97;
/// Ie86b28b55eaf8feb03e24730be892314 I31c6b3fdfaaa80dba2dbf92a4600524c bit
wire [MAX_SUM_WDTH_L-1:0]        I6c96e6686c458cee66b9d93d6d71f350;
reg  [MAX_SUM_WDTH_L-1:0]        If46fa11dfadb0691eaaa0a40836e08d8;


reg  [MAX_SUM_WDTH_L_P1-1: 0]    I748f85f6680918a2e992df339b4b6558;
wire                             I204375b1fcd1f62621b32a06a9dd0bb6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ib0f57837099e3fdf1b908d78bcda4a43;
wire                             Ic0ae28dd2fa2d9e0b2a9edaaffd88aff;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If75e99660e3997f53f7b903bc366f47f;
wire                             I63323f8807804f4534429d8aeafc7d23;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I3253481bee7dbfc0f3eac94c3252ee4e;
wire                             Ie8554592e62dd20a36ef79e06af24a22;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia80693da8182ee2c3708b6ec21d397d2;
wire                             I67458f3b57d906d3626d4e7656049538;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I7fa3f2648baacebf9e4b59c179601fa6;
wire                             I523d96cce3a523da8ca8e065aa5d8f64;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id7699f8f89380c315303644fdebacb32;
wire                             I3fad2338742a91d05694c9bbe0584126;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ibf3e1ead3776901898d4b154aeb61267;
wire                             Id30ee39232f016f983f45208ed802126;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ie486617fc1d6354c7f347692cdbd894d;
wire                             I149dbd0f3f68786fc3a842bb0064f0d4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I7ba403c6745e7d026282ad704e065702;
wire                             Ib383a8f851cd16df009c975ec7efb305;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I93cb3974b8594665b2e7ce5593fde69b;
wire                             Ia2227bb2140f18af451ea4c397262178;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id6a9ab06d58c3a01e1fe04fcf61406fd;
wire                             Idf0b6d7bfa5a9a38e1362c4b3b0d5b99;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I261bd53528b82128acabd405389c8d60;
wire                             Iaa15139339207505f231f71669ce022a;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If7fa833bf1b1438e7a5bc783ee745252;
wire                             Idc30dece6bd74ad2ff6c0822347a800d;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ibb103853fc21f8f3d466ca16557ccd3e;
wire                             I7492572ef50294af38fc778e173a60fc;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I37446eb66ccfd268cb418655b8160fe1;
wire                             I4c6718b74573391494789da2e33c1e2d;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id17f6250f8c7f1d7f75fd27f92698da3;
wire                             I03659b77af3e47129d9206af314ec521;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I9957b02e8d0d888e6950eb553d9084d7;
wire                             If0fbb2a55965bb66cfaad70fd9241456;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic71258b745437bc8463fb4f847c55e27;
wire                             I4f8bea1f3f8cb9ff1b6d1388c6377861;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I24bb5c315eacf0f4e8c86f6582389e39;
wire                             I765559024522a12448e338401c10f800;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I607f203694ff76930cfee4103cb73c30;
wire                             I815daf68a1ed9f91b02ede68298cc5f3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ica8e4c56ebb37e189ca8e6b3daafdb80;
wire                             If0e526189886cb9e8af7be4797d8a637;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I7089386c94261e0febf3b4f7dc1aec30;
wire                             Ic8dfeb5746649e88e59887cda08fb62a;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia1e4f20f32f7371cb0078d6e80fe8b7e;
wire                             I0bd3e1beb510558b20c2b4f0f8f20e76;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I790cbca796af58b1726d0a4680cc164f;
wire                             I647c8a9b1fd2281c8e129d2cebdd597e;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I0a93f095f9efb1542116a295c0db9c8b;
wire                             I6a803347e6d25dbd012caf725e35c256;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I989ba39f188a44475a83e65a4960d2af;
wire                             Icf6deff8d81d69b92659b257bbdb53c7;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I9bcc1d9b3dd258fa7b6042f0185d48cb;
wire                             If282e264f908747340e4e4d2022a66fc;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I9ba14715d9f33ef45681ad52f5be9593;
wire                             Ib5ca6dc87c214c3d73b265fa0e242452;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I396a897f79b519f4fa02af39d0274f64;
wire                             I3b8dd3a8e7b21202977c976ba687cb7c;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I197c0cd576e16ee2197a28c86397f801;
wire                             I4e1743e1634bdb7ad6e8d072e19f0abd;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I094a178e55425f27ac1ff6195217396b;
wire                             I4ccbbd7d8e03a7c7410acaf35ef87608;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I3177408f7d08b431be99297fb10586e6;
wire                             I1848d733a31c474bcb2d3e4b9b736e94;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id4948c876d48bdbf317d32f135e645b4;
wire                             I6fb841a6fe0ad7d433f1a182706d6ad6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ice5ff01d4fb4583898498651a0ac0171;
wire                             Iddb16107d5ce4ef65024a1cd5387dcd1;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I0fb33a5ced3d15622c9aefa188052e24;
wire                             I8eb4596c73d1cb6ae5a783a6582cbffe;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I0074e1c3ca0ff903a9201ac5fe7ca841;
wire                             I014c1931d012f79e954a12e10178f1d9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If65f587e987a51c093e8dd4df532e26c;
wire                             I8ad79c41a8896712d7c26d29c0b1e7cf;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I33d7e77d08590f0dfb1867e741dd8b6b;
wire                             I1b16bbdd1e23bbe571bc7769731a03d8;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I678c22563e0273403b046df4261f21cf;
wire                             Ib0cea939898e64f9ec4ee41aa3f062fb;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Icca700c12ae2e8155ca6b41e692e8a8c;
wire                             Ief16fc889b2326a53224b3b60ecc8955;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I5ed74e81d2497681af5a0ca13fe23088;
wire                             I774b99eb9e3c3c98ce6dd3c60df7eff5;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f;
wire                             Ide90044338620a38b90b5877ce0eb52b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I26010e26e22d8a2ea831e86fae34a24e;
wire                             I2271e9b3a663941eed3b939bf80ed2a1;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I578efe5c2c504f12c8f2466a7f734215;
wire                             Ifc1b458539905b3557d79c94954747c0;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ida86d05f907d23ff9fed06927c2ec9d9;
wire                             Ibe27dea48dd30331b9723a1aec226f0f;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I9d9f8c7a23d9750ec44e706bf763df76;
wire                             Ic214eae29f89949c797816779332aef2;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I0b41b002a32b8e9e2fe68e819f228fb7;
wire                             Icd48fe364089e0250b4fee636590fe28;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I0e872d4c07169cac84549178fa144274;
wire                             I15d7c9e33bce9e3ee1059f73832bb9ad;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I6f4ef0f404ae046519b8436171d51e09;
wire                             I9514bd70ebe24af7d8bf346ae09219f7;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I4d04e66ad9103a685fbe088b74517452;
wire                             If987109479436b8d51629513310a948d;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I988e525020c1e43d238fad41dab4e6ea;
wire                             I6a91c509b367469511d65174ad4e3b44;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I90d92887cb2526a2956d5e8c9fad760c;
wire                             Ib0fc75acbd769930a34393612c6f4fca;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I00fe3792cde1eeab36e576fd6634c4fa;
wire                             Ie9ac51d5e0f07e135eb10651d94829d4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I6e586c5ac59a28b30c377e51287bf04d;
wire                             I6faf08de30d6ba38e76cbf7c868a6f73;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ib5dc74106d8841d25a793010fdac599a;
wire                             I6a5a58a73d0557e080e6327ee386020b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I3eaf142d2734d2d0decef084dc037b50;
wire                             I3704ac8ccceb7a319344229dc2db6693;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I2d171ad83e27a3745d204849a6f46954;
wire                             Iebedd8e3b4af888431e0a294d56c5c9f;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I977f1083f5e4f6f8ac38e2c5aecf1b79;
wire                             I7bc366f56c020144390350e85747a6f6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I9bcd673a4293e14fd20b48fa20492df7;
wire                             Ia3252e7c4f3897ef6637bd063b00d3c6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Icb7422ea46b22b9330c123b40fe343fe;
wire                             Id135567b50e17e28d140be2906bfe185;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic414cdba230d7ea73972b0eda1ec6b1b;
wire                             I3e5c9230c5b091b31ec13fddaea37a8f;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ie4e1e00503dba189b0f871c3c0810d76;
wire                             I1c3a83518d660eb2549b1b8d2a2f6186;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I721c43ab62b42a18c3f5228fc0a73262;
wire                             I86e509fc0160543f825aefa4dea4eaf4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I1f7cb03cf806b247be1cace4d75de942;
wire                             I6cb732a94dbf7bed4e70f4b6a1c393f1;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I775cc766b069022bc00220050feee4e4;
wire                             I0d3ce639167582d0b25085ff5b98f7c4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I08b78f774ed494fa7f119977bd92679e;
wire                             I7f786778e022e1cba9aa7032c0d43db9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic7dc7f94af108ca7c8003a2d07e1e168;
wire                             I4722e6750746bbe43018b591688ac3e9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ibe1327961152cc2d26b3f19476a6e2c9;
wire                             Ie320d1535571a2af4ec61057258a60b6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I5ba97de444af4e8c9744c3b707502edc;
wire                             I69c88d14b5244f55911e23f7685f37d0;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I3e4f1314042010b5d7384693b580da7b;
wire                             Icbb724c2e16e099c0820935ac4fe21e7;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I4a47ce6e21c1a274578397e480c184c9;
wire                             I01b9e488ff0277a2e1e8b52004e4cbd3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id184731beb200ad6a53ce273b963bb3e;
wire                             If329f0c1b6d206280da518bedeb1b5c3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I3317f2f6eef9a8ef1fe1ff68b47c5d03;
wire                             I47e322cc161d674131f11ca70479c538;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia6b9fa10c79e6f3847f89b35afb4cc59;
wire                             Ib343e5b8ebe704ab55692f487b06c156;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I91e98b804ef82eea53c5e8eccfec827f;
wire                             I1a6bc8e0684efd6ea5f73651688f9cc6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I5f1e0d0c6b50f70a6f5584124e095501;
wire                             Ief7890423e793f41bf2b9f27ff47b4a3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id61fcc605b4b581f5d42024c2610c8b7;
wire                             I145a313064c4d2c5c30fd9458bd32d56;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id64738b7668931553151dbadd5605b71;
wire                             I2dfaa00d2d1869026f6c8651ad8cfde9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I3bdfb451eb96d256da542864d39024df;
wire                             Ief703cb630f99bc2d59ae0e27bfb3572;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia740d8ccd8230b28d078b2ea3e58d6ba;
wire                             I3c5c01afc7096f90c8c6f875dd9686b0;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I574050722f82569d34bc2cfae1eedaa9;
wire                             I5ec91f70ba0346f55caacb7e78f714d4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic8f7ec6ee09fb9ee2467e3cea30a44a3;
wire                             Iccf8ad1402095a65a32897af9d8ce23b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I2b77d922a74fdcef0d57debc789bd539;
wire                             I18950ce49f50b9fd4aa6b1d69b162fe6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia1d8127af4944b23475bd7deac91d60e;
wire                             I6ad8cf59d777a2e6832471a2cb713eb3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I247abcede9914633c0a33fc402bf58ae;
wire                             I8d24e40d6e2c96260bb58024eb57765d;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I1f413d3e081c6aea012b122fc94f73d5;
wire                             I7ebb24e284f0aeb792723e15024fdd7b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I1b812fb764d3b48511c0d15a7efaea29;
wire                             I717cc8e9bb50878c67c3cef72088f279;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I88882bd8a9f8718411564221ad85b223;
wire                             I9140c28397eaeffd7a3446096bbb8419;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I232f24e2798488ee66003f3b8cc294c0;
wire                             I1563ae311393b429f4fe42180f1c61a4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I856284e951773518eb6c4232ea7f3d40;
wire                             I068dc4e9969e691dec22979b38ee588e;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I82cbeaf5b3e4796b2aaf33dcbd119f4f;
wire                             I9820fcf4305469c0390cf04be00ddf1b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Iaa7791bbc193412e5fe25000ceec23d6;
wire                             I24a3a82a62c3c1348663e84e1d80de10;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I44bdc0baed3d51ef54ce2728618ad339;
wire                             I10b2505a209c84c3468bf8c5564ff7b2;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ib6bc7e75ce750a26113cbb8895c2f024;
wire                             Iac33806e51f5fcf8e571bfa02272151e;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ib4188380f7e96d5afb99f5045674193d;
wire                             Ib0f7718835e96a6b3ce6e7eacc5ae37b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I5bba219c5024301e420e9a5acbdc5845;
wire                             I68bcde39ac1f26fa5c8daa7e616b7924;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I1bb52988c9ba03e16b1b69335d3d7e7c;
wire                             Ia320bdbc669ece554e4dcac16a650551;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I1b9990aaeae716f66b0f89fb02be0a74;
wire                             Ic31b8782fe7655bf0dbbbc034acaf00c;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Iceec2cf6aba9138648a3340390f39fe9;
wire                             I7f1175afac88a045954988d97e6c014a;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Iad7842f3d4672f42c1064c28d4c8ec4e;
wire                             I2aec42e2d6c3389d51b99855f4b31413;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ie5a53cf9343fdcdb5788667c45fadc83;
wire                             If6053e257420db5a04d9864730adcb98;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I30e06d190906bc9eb6f1c3156c47f9f1;
wire                             I107da1e40d1217df6353e403066bacc2;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ieaaaced47e22029ad2945eac9cc45e6c;
wire                             Idb29269890e208fbac5a370a883f180d;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I08dc6f8e837b1f6b80bd3fc742290dab;
wire                             I5ca6297084710e3fc6d343511e4c8e42;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I8eb6a9c907c5909dad6cda98022d70b8;
wire                             I586b30878699ef8f0d09e922262a19d4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia5067b1b458af82c3c2cd50653099854;
wire                             I2a833dfb485a2a420a799ef5854b1dee;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I198c6753cf12d423c709d1512e66fa9b;
wire                             I598ba40aca3b048d684323016e46c777;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ib600dd8a39fda48d28e1289d44d49a84;
wire                             Idfe3a41188b5115db103d16bf7b4417b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Iabf09191227584c76d7fbc634b706d12;
wire                             I7679c765ab544db47fae6a7867974d61;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I4869ba08cab90a6dcbc454b0001a7a20;
wire                             I30afde55f450fcb898f5854004d618e9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If97974406672507f8c9a1c507c4b6951;
wire                             Ic216abe8348824570dce569f4ff9d186;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I4210341f99ac7cb08245137999739114;
wire                             Ieb0dc034a1be9a5d3f2919b4d00d0960;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic24f4dbd99c8f4d88c8450d4fef762b8;
wire                             Ia4a51f9d6b4d72bc7edc29acc1938b67;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I68dffa1a13eb6ab54615347729c1d6af;
wire                             I83757c2cdf0e4516bdafb5f6b4760aa3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I10153d5548b184b9ac2cecdba4ec4b1a;
wire                             I949a414f7676d024a216b21e3d1a9cac;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I104b7f0512440cffc0fcce25e477f537;
wire                             Ifa3590aff64fc8ef90046c547e6e6f88;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I18b6758319272eebbe76e1eee5ae55b2;
wire                             I133c6136e389a5bee5a3006d939a0a6c;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I780263b10b98f9bb0eaf66c045d8d37c;
wire                             I4b615d38e855bc21d809e3e5b24732b7;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I37b772442e55cbcd44ba892a0608d662;
wire                             Ib8e420738c31144696b4cf90eb99e270;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I0ac256a6659ff5c6673fd110a8bf578f;
wire                             I09a993ba748562fb5ca4df9f36f683e6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If134e1d27e736005e5a390e7a2ea1f4b;
wire                             Ida3263e09545600a85caf500b5cba32d;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I7b37b8f908cd82683832536e02faab0d;
wire                             I55f6d7a4bbd8422555543abe0171d576;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I08b4bf60c9c7e7229bd1952cc88bc7b3;
wire                             I9fa0e35a8ecacfa315845aeb73ccbab3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I267d637eb63fef9f4723f7978fad88f0;
wire                             Ifdcee23865377289dc0e9986c92325be;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I4fb56a70e5ffa71f58f715da36368e04;
wire                             Ic8ccb35ab31c6d17b98e5f63c022d187;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I5e9e2acb258baf96ac4b525bba54a462;
wire                             Ibfaf924a5a317dbcc967127e153d56ba;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic40f61443a4d8f87769067fc39381cb3;
wire                             Iedabfd30e25648ea4e62808e1922f016;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ieb36710c9a3726f33407436d62639c8d;
wire                             I437ac9b58f5e248aebec968c948c4125;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic804af393da2e4b9c8ef25d4a3b4e8d5;
wire                             I0cef2090a761574041a230f80dfce8f9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I52e4c446693c29a42bb3b665f72d382d;
wire                             Ie25a0d7f0c4b7b25ecffa8af65866f60;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Idbf02cf10add496d30fa44bbb18458c6;
wire                             Id33e269cf9da206ef2c24e1eb4a1184a;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ida095585ad26e215f1c1bf989912da89;
wire                             I9d21b9384524b55c2eb70826c045052f;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I19f1ffa05c7c9a0df5e7014044024c7b;
wire                             I1332e87f7d43cae554ff461d3957edb9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I4d68a2fe778fa93faac38b138138291f;
wire                             Ie11bc6b5b26c889cf8d2236c17f9ca98;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I54393ada6f76ac82c31f2668e228e29d;
wire                             If1cf7892a4b06f5e88f3831ba6bcecc8;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If5b9ef84f09680f3593250b13a852c1c;
wire                             I76a07c1dc9d6d51fe3a31ea3a58ef916;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ibb759bc4179e5b7aa759d850c7cfa467;
wire                             Ia51886b7fca8fc0eda0b93c40d8ccc64;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I05e8b5f8b83f07b609b5ebf272bb2229;
wire                             I48c3c239dfc925169c61fae6fcd16eba;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If6ac15373ec1146d38e7aeb71c3ece64;
wire                             I87a5898180c3b4934fa6d4832b6507d5;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I2ab3675e1eede757af80716ba980a4e6;
wire                             I18279e41940f794e7bfcca8062c42ee1;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I388c271687ab31b57421ad57192273ed;
wire                             I04cc6e9d889d548aed3e517b1c7a98a4;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I6121679cec8caa51dc5ff0d1a61f9821;
wire                             I5b319b9f50e43a7c850594b015d24ef8;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia0649b990bf5716cfab230127cd5d47f;
wire                             Idad08f7167bd930530e12f9180bd576a;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I867a0626ca22108b16267d95c0aadf4f;
wire                             I044b9326d592e52c74056c2385d9a07b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I1af54bcb73d7c6b93e55450871207976;
wire                             I838a7c657b5ddc47cce2b9fcbd433548;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I91883553543d0425e9c6dd726dce3d27;
wire                             Icf019d30479d47cec2a9508e6ac4882e;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ie95405659701278e3f87bf1f823a037b;
wire                             I344dd9d785b1ec8f6c3a0d8fc1f400f5;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia42392e2104b50c0908aad82738a5ee7;
wire                             I380dd5278a22dbf0fd4b86985f91dd6b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I68ad63230a51b9b9e3daffb307ea970d;
wire                             I5feb2a46a916f5ed44638712d5ecc3a6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I7a052d63944ccf42e598efe3a95b88f8;
wire                             Ib184353aaeae5ef036ff36d0bd35a27f;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I2b3c6d69f79c8d51e4d1614c62c44fcc;
wire                             I53729ddbc242ad9a8724d93648868db6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ifcef0e92f50e3920bf1208af5d64c632;
wire                             I6429512833e3251e949ad734bfb1dbfa;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I111340a19625901a3c1b95fd0bd1570e;
wire                             I96babc82431ae1d3713786eb68c2e372;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I11aec4fa85c30f6fe1fd9fa72542ef6c;
wire                             Id76e3859fce7aab300a173587243b0a9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I80cc333c181c16a96b7bd6501c27c2b3;
wire                             Ie607dd51fbd545d298488a6e9c9430c6;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Idc6354325a6280ae9890da33c06c33ec;
wire                             I00e222e2e16487cfbac6206d913ebc21;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ibb04cf82acc4ac16599ad3ddb0c2ada2;
wire                             I400dac72f25c87765a07e72c3d04240e;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I3ed096dfd8a14f4acb4d53a70cf8aceb;
wire                             Ib0b26ab3c5d3109999c55b41e8399c4e;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I0fa07f95e96326cb0599c0c3f76e2b48;
wire                             Ibd55c6f55d6481b76591e2c565217e4c;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I87d98fbc97d9a78c2e7d6a6280e7a49a;
wire                             Ie5764d99afa00cd108404de18693c4c9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ib7ddc4dca877f7cf5697a02c3d1915ba;
wire                             I5234341950ae6353868b35e84b0d837b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I3612ef280891f6017fad205d0484bde7;
wire                             Ice8048703f0f8018353d8666516e2b7d;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I561547649aeb5b4c3f10d9506db1f3cf;
wire                             If4ab153a2932d079ae16480dd788d298;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I84cc76c0079b86da7b994844c3ccb875;
wire                             Iffdd32b08a1072206b9b83981560b341;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Iec013c508d0c6401d7eb856e7eb60446;
wire                             Id328a2bf60eddb0da7bc9fe44eb81163;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ifd8979aac6b6b24aa560b46b18240e92;
wire                             If39c82e97c07c30522a1b489ec896577;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If12394e78dc913b01890b56650856a44;
wire                             Id78ace2bd65545c4add80a2720338443;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I94d18aa10695f3f22b23246884b72822;
wire                             I26cd0e322d30abad73493e57d4157954;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic90b38835dd7e760dd54067b196f8470;
wire                             I6d27a778e8595666903f4d20d47dc053;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    If3691ea51f6efe9b165a31964854d2fe;
wire                             Ic220ac5d53b5c26985e5c7de2d95d896;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic2ce582555add38a14f5006d3c87eb15;
wire                             I9793ca0ff4f0324792cbb1da51d60904;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I58cc950ee2cbe56b7c5a619be3792511;
wire                             I76b19931a9589b4658dda1384f13f30f;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I0d8e329ec5873db96df1ec309445a096;
wire                             I0726346b2914d4aeb149e512d31af95f;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I106325488e2ecfdba1cf9e5201e6bc8c;
wire                             I399c5a08f19fda00d218b1fe4376eb5b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Iff73a0085541a511d3912b64686a82c5;
wire                             I7c3e36e47bc35c16a8420d88b356e9e1;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Icdab59de68f2870504598c9ea18f1d2c;
wire                             Ia0bc5e9d76d19f62b221c666f533d959;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I75604d727e82c977741f90113719183a;
wire                             I366301d215cb0f4bc390aa6a5726d86b;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I6f50c4d0d2639857b2dcca300c2d7b04;
wire                             Id039bdeb594da7428838b1dc4d6af8c2;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I5cd013a2be2e761c10c6a957632517de;
wire                             I2df05059b08aa3babba9542b51367c83;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Iafeedddd02428bd2610c576e68d4ae25;
wire                             Ia0a811eaed4d73f4012e1fb6217cbda2;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I912d6325e34180e0f668f0f024e63581;
wire                             I43333dfaf1cd037fd6bc16d290e0ea86;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id1e05294dfd02df499ad0c08bb5c191b;
wire                             I4a7337b53c190d757d250223ede3daf3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Id3bb9b100ee4302473b49ac14615e9b0;
wire                             I49d3d7a17c12933457f26c5232277395;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ief32db1cfc443119b6202b0cc7bf70a2;
wire                             Ife2b1721d683a43be53c43e49d96e0f5;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Iad7dbe9909b5eed3261adf92d3813acc;
wire                             Iecf2a3bbabca3f1ee3c9bbc3ea3d2083;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ie7daf0789c35caaadbba06cafabd2b70;
wire                             I388f3758e343ea6ee2ca6c14a6a8afac;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I2bd1f9b75d9ab94af9ddceb7528935e8;
wire                             I70754064855cd8d49164f5a24c2087e7;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic3d9f5c6677758810e4865779ec303e3;
wire                             I9443c16fdec0687f97a3fe287787e4b9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I00af04882a25e2832d913a67d4d86d7b;
wire                             I5d871bf470d68cb1651c695f14a2dcb7;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ic9db631df0a1a9108c10c3e0eca7bf15;
wire                             I30a21066d0f7ad97b21dfdcc42fe3aee;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I749f9ed1fb2dddd40ebc28f638e02935;
wire                             If0cb066c4e37fd6772da2ee943543829;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ia45b2a24df24bd5e3c95885c8928686c;
wire                             Idf3132bae12e52ed9560eac88e2ead65;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I7427464fde340780aba7f9847b4ad564;
wire                             If092511da36f3f493f7e3f34a35cb9eb;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I33fd1ae225e2b881b2b41e0358675e22;
wire                             Ice07207e1867f71dbb58dc0b3d28f5d1;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I2e21a35d1cf560936fd19b944a208b6b;
wire                             Id1c6ccb54bf2d0d03f296cbd502fac6a;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I249522a3d42cc75d7a6b9ede1222ee76;
wire                             I7a2b0491133ed6a2daafb889ff46d271;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I68b4c43d9f40ae4bfd70d2983594392c;
wire                             I4fabd40b7afb192a9c2a255512fd0852;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I63145e0fec15c7e7c0de105f348bfd31;
wire                             I7b39e709a6939751b11bb3ba6fc42bde;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I8af625de86c04016c3424d116fddab5b;
wire                             I3a7a76b3ca144951bb6edeba1650c35a;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I54c9c10527f83b4ee4e1e22f1e4044ed;
wire                             I3c023a3a1a2ce2fb54b2292401df0019;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I972559e47c7f83bd9000ca1cfc14d8e0;
wire                             I804cf7b8b79a124cbee51fe473e664a3;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Ib97a7f941eb7ce2a867503a04ff86a67;
wire                             I33be2a0d4c64f50472091a4503281558;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I5979b55f607c71017537f2b48b40cbea;
wire                             Ie5f94955ed10ae50d92d3dd0e43c8088;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I6a56760b621f238843b091279c69897f;
wire                             Ide6f35e8581e1bec17ec974448b6beed;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    Icec45bf76c241d37c9a50a5cd092da9d;
wire                             I57b47b934005413e4c400a33e7ddc20c;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I2f6d3f61f2890e584d3063a09587e99b;
wire                             Id4e7f9a0c100dfc591e7693d76a496d9;
reg  [MAX_SUM_WDTH_L_P1-1: 0]    I7c396ea2e959d84fd9a6964617cb29c6;
wire                             Ieda30691eb70678f7535eed71e9ee031;

reg  [ 0:0]                      Ib0973b6e90e7678addcb064fded7ce0f;
reg  [MAX_SUM_WDTH_L-1:0]        I5033323484d90d6bfbe03749019fc6dd;
wire  [MAX_SUM_WDTH_L-1:0]       I97afe24956b7f87cd431f048202bab67;
wire  [MAX_SUM_WDTH_L-1:0]       I117235e3ac8e68e4c1ab34db1612aba0;
wire  [MAX_SUM_WDTH_L-1:0]       Ifd700cc9d18f99b63f1947f3ae631976;
wire  [MAX_SUM_WDTH_L-1:0]       Ifffbe3d1007fb07a20d3b37902b3ec95;
wire  [MAX_SUM_WDTH_L-1:0]       If5443777169422ea6e1e3f709b970e05;
wire  [MAX_SUM_WDTH_L-1:0]       Ifaf9fc93e4609d818aa46751754c17f1;
wire  [MAX_SUM_WDTH_L-1:0]       I419caf964986c655df84d043badc37c9;
wire  [MAX_SUM_WDTH_L-1:0]       I3095214ac0e6c1323e75ee4ec85e6821;
reg  [ 0:0]                      Iee06707670e19a82d911c1750bcfc811;
reg  [MAX_SUM_WDTH_L-1:0]        If5dad13ac41b3034bdb034bc86c9b348;
wire  [MAX_SUM_WDTH_L-1:0]       Ided9739bf63937933250a6d0c37535f9;
wire  [MAX_SUM_WDTH_L-1:0]       Id0f139b9f3848b45554ac8429230eea2;
wire  [MAX_SUM_WDTH_L-1:0]       Id9feed58cf9565255abfd0bf7e3ec068;
wire  [MAX_SUM_WDTH_L-1:0]       I30a3be3b5f6ad1880a917eb35659a1bf;
wire  [MAX_SUM_WDTH_L-1:0]       Ie8148d9aa962a733eb65877b902a187d;
wire  [MAX_SUM_WDTH_L-1:0]       I69e98cf3e679183aef6005bb582b18dc;
wire  [MAX_SUM_WDTH_L-1:0]       I7f42a504fc61c9548acebdd8b1858eaa;
wire  [MAX_SUM_WDTH_L-1:0]       I08b1b4639b5a9ca509b943b977f6d4bb;
reg  [ 0:0]                      Id8d5df9e869aaeb107a41a6bca3b89bd;
reg  [MAX_SUM_WDTH_L-1:0]        Iac428f9f798618e1ef495c626c41892b;
wire  [MAX_SUM_WDTH_L-1:0]       I8d7296627d886566783e79c01b9fa423;
wire  [MAX_SUM_WDTH_L-1:0]       I4fc4c97229a8b1f631a3b505941159e4;
wire  [MAX_SUM_WDTH_L-1:0]       Ib9b16bf51891c328dba2699eb9bcef95;
wire  [MAX_SUM_WDTH_L-1:0]       I6c30501ec81fce286817788d614a7824;
wire  [MAX_SUM_WDTH_L-1:0]       Ia4d4f37baec48121a88808075dd655ef;
wire  [MAX_SUM_WDTH_L-1:0]       I385495ea2bf6442a95ab7561456254ac;
wire  [MAX_SUM_WDTH_L-1:0]       I5128e03d383c226befa6f7422f3a6f04;
wire  [MAX_SUM_WDTH_L-1:0]       Ib208908bab4c20713cd17e20139c8db3;
reg  [ 0:0]                      I507f8602a99a1096e4c293ba3c235bbb;
reg  [MAX_SUM_WDTH_L-1:0]        I5a6427c8f18b36d2ea18fe60a0831ef1;
wire  [MAX_SUM_WDTH_L-1:0]       Id939992b99a11c09f4688c10ca1a34d1;
wire  [MAX_SUM_WDTH_L-1:0]       I823453ccb90d5b2b2d9dfc6e8358224d;
wire  [MAX_SUM_WDTH_L-1:0]       I279c5c00b92eb1b872b5afa168b0306e;
wire  [MAX_SUM_WDTH_L-1:0]       I66f25b1c3c0eb226295179adcca2c3d2;
wire  [MAX_SUM_WDTH_L-1:0]       I3068627e91b667d14cd3e55a9371931a;
wire  [MAX_SUM_WDTH_L-1:0]       I44c4e0a2d8a7289f8660b81a9ecfa19b;
wire  [MAX_SUM_WDTH_L-1:0]       Ibe868e258dc87f0dd1460ba6b8354671;
wire  [MAX_SUM_WDTH_L-1:0]       Idc3083c3021200345e3edd35a9d4725a;
reg  [ 0:0]                      Ibdf2178bd18783c4797c21e642388d16;
reg  [MAX_SUM_WDTH_L-1:0]        Icc29441eac6ca7a138d45743d37505e3;
wire  [MAX_SUM_WDTH_L-1:0]       I320d4f19a5b18c23ff407508d47caa77;
wire  [MAX_SUM_WDTH_L-1:0]       I16becf3c92615d98d5ec51ee9641cc0a;
wire  [MAX_SUM_WDTH_L-1:0]       Ifbfacc3b3a0128119943bcbf80176612;
wire  [MAX_SUM_WDTH_L-1:0]       I6b4f670c9e8e25984e8891f2440322ab;
wire  [MAX_SUM_WDTH_L-1:0]       I19bf0990a30c72421f231772b8627e8e;
wire  [MAX_SUM_WDTH_L-1:0]       I3ec3eb096ebe3ee8a47e1cba6487b997;
wire  [MAX_SUM_WDTH_L-1:0]       I7379ef16405c461ac44b66c4315df831;
wire  [MAX_SUM_WDTH_L-1:0]       I79db45b23d21d533a1f9a6e8f94d403d;
wire  [MAX_SUM_WDTH_L-1:0]       I0979534730cc2b53547d413dbb6b75f4;
wire  [MAX_SUM_WDTH_L-1:0]       I5aa2f9c0667d1a6e871efbd4d2bad3a8;
reg  [ 0:0]                      I2c690809d9b9e3482fe5a133b5c00afa;
reg  [MAX_SUM_WDTH_L-1:0]        I0e7754dcbc04a4850e052ae4a2fbe328;
wire  [MAX_SUM_WDTH_L-1:0]       Iadb28dc990ccf2dd3099544de16b8f16;
wire  [MAX_SUM_WDTH_L-1:0]       I1f71aebf698788d6ada66891e9ea756f;
wire  [MAX_SUM_WDTH_L-1:0]       Ib234e9cf7e7616a1ebc6ab99df2a7ccb;
wire  [MAX_SUM_WDTH_L-1:0]       I297d1edcc583ea4d69da780150f0620c;
wire  [MAX_SUM_WDTH_L-1:0]       Ib0a717cbb4fe38a3fc85520ca0826fd9;
wire  [MAX_SUM_WDTH_L-1:0]       I037ecd5945b1f1280b4469d73fe1c7ff;
wire  [MAX_SUM_WDTH_L-1:0]       I367ff6b11b884e02a3065fc7fe811e15;
wire  [MAX_SUM_WDTH_L-1:0]       I6fab19692b512166fe9c74b5e987788d;
wire  [MAX_SUM_WDTH_L-1:0]       I04dd73af505f618ccdb209b3cf97ceec;
wire  [MAX_SUM_WDTH_L-1:0]       If8c559905d4120488d431719c4e8ce24;
reg  [ 0:0]                      I369ffa98995ba0834f8029ecce705c56;
reg  [MAX_SUM_WDTH_L-1:0]        Ia30c019ed8ce395556494a92e7b42a92;
wire  [MAX_SUM_WDTH_L-1:0]       I20ed4f6f14e20ce3f0e106d1b7782fcd;
wire  [MAX_SUM_WDTH_L-1:0]       Ib10626ffa126188c5bf1fc8399107b26;
wire  [MAX_SUM_WDTH_L-1:0]       I29007c52357ac7afbda39d72a5bb60af;
wire  [MAX_SUM_WDTH_L-1:0]       I66d367c046611f145e607a90911cf499;
wire  [MAX_SUM_WDTH_L-1:0]       I9c4c2556f6170a8df61d909855a846ed;
wire  [MAX_SUM_WDTH_L-1:0]       I6fadc3e8d995bb4317bf7b4377c3c2c5;
wire  [MAX_SUM_WDTH_L-1:0]       I99b20e911c189e0616f02376ab736e91;
wire  [MAX_SUM_WDTH_L-1:0]       I5793c12f5dbdd8245dbb202d550ca960;
wire  [MAX_SUM_WDTH_L-1:0]       Id0660e9637cad1ce1a73d37188060154;
wire  [MAX_SUM_WDTH_L-1:0]       If5a7af7ca023e1393526e888f4220a44;
reg  [ 0:0]                      I9ccef4c47ae7cfab43584de0f2e193d3;
reg  [MAX_SUM_WDTH_L-1:0]        I9799695ea8244992a6694eaf5c8ae64d;
wire  [MAX_SUM_WDTH_L-1:0]       Id043eb50634e803e53adc1168379a5d0;
wire  [MAX_SUM_WDTH_L-1:0]       I1f866dd0b129267550aea1a267d9c91e;
wire  [MAX_SUM_WDTH_L-1:0]       I8c4da05c08210fe33139c3d3e5d75d58;
wire  [MAX_SUM_WDTH_L-1:0]       Ib41f7b823681fdd084b6d8436a407aa8;
wire  [MAX_SUM_WDTH_L-1:0]       Ic5b50a785b7acac7e3be4095aa92e50a;
wire  [MAX_SUM_WDTH_L-1:0]       I3ffbe03796b66d00d47fd918be60ab89;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc92a916da938ef6164db250be635f88;
wire  [MAX_SUM_WDTH_L-1:0]       I8ccd42508ce7d5bd897c2cf0c54caeb3;
wire  [MAX_SUM_WDTH_L-1:0]       I4920e7e82749cc036b58a7cd0a03e327;
wire  [MAX_SUM_WDTH_L-1:0]       Ie1040b2aa91f272e4449c4b5f9f8f575;
reg  [ 0:0]                      Ief31fe169c1b360d5933558208dbb602;
reg  [MAX_SUM_WDTH_L-1:0]        I4524cd664b4cb41f642c675fa484c84b;
wire  [MAX_SUM_WDTH_L-1:0]       I65968fb0f63d52ad96cd8fa270126a1b;
wire  [MAX_SUM_WDTH_L-1:0]       I839ac8ee59f51d4c3de92ba5cb26e788;
wire  [MAX_SUM_WDTH_L-1:0]       I33cd95f1919318a0f3df5df7310d64c6;
wire  [MAX_SUM_WDTH_L-1:0]       I4933e8d16fba26cd797b25a9ac2a2de8;
wire  [MAX_SUM_WDTH_L-1:0]       I218f7578eb748e31d0002052f30c5842;
wire  [MAX_SUM_WDTH_L-1:0]       I2a808d1c42ad758ae3baaaee8129dfb2;
wire  [MAX_SUM_WDTH_L-1:0]       I4e851fd3c114af87f5e8c68c02594e3a;
wire  [MAX_SUM_WDTH_L-1:0]       I0da40f88adc46e90f616acdcdb8e0e2c;
reg  [ 0:0]                      Ib8c0317dafcfb91b3da5eb5afae1f2e2;
reg  [MAX_SUM_WDTH_L-1:0]        I64e959d80af111ed2fcd54a5407d21bf;
wire  [MAX_SUM_WDTH_L-1:0]       I0dee7767e472a5fd71250ae6c57cc8b5;
wire  [MAX_SUM_WDTH_L-1:0]       I9f40be7552b3dd625e5bce0befc5a548;
wire  [MAX_SUM_WDTH_L-1:0]       I8fdf98ffd757c8845ed6ffa4ddd1a16b;
wire  [MAX_SUM_WDTH_L-1:0]       I8103b777314a4fa471e0898fde9cde08;
wire  [MAX_SUM_WDTH_L-1:0]       If6c3ee8e0d7dea58043d5be0f4630873;
wire  [MAX_SUM_WDTH_L-1:0]       I711a5171f591f472cdbfc9a0f5e1aa17;
wire  [MAX_SUM_WDTH_L-1:0]       Ic30bc38184dfbbd694af52640692709d;
wire  [MAX_SUM_WDTH_L-1:0]       I422f6fd1d273a3834d04b04ab8e2812d;
reg  [ 0:0]                      I54e3f08f6f4cf784da57ac39f246b8fd;
reg  [MAX_SUM_WDTH_L-1:0]        I3e0da4bcbab4804b5397fb3aa2c94f51;
wire  [MAX_SUM_WDTH_L-1:0]       Ia0fdc60b90ad18b6585ec1ad4e89e80b;
wire  [MAX_SUM_WDTH_L-1:0]       I7809fe7a30d041a7e569ffe890242df8;
wire  [MAX_SUM_WDTH_L-1:0]       I672b14ec1b3c4797545f266727505a85;
wire  [MAX_SUM_WDTH_L-1:0]       If9620d20ebaae6245a2c386d9bf5fdb1;
wire  [MAX_SUM_WDTH_L-1:0]       Ic74e22bffd88f32eefe499cde0fafa8a;
wire  [MAX_SUM_WDTH_L-1:0]       I76d38ce67387bd76ab45c9cba7d18b31;
wire  [MAX_SUM_WDTH_L-1:0]       I44413c6f6f6493f8a86abf6eb32604f6;
wire  [MAX_SUM_WDTH_L-1:0]       I67f632fca617fe06565ddcaaee8fa8b8;
reg  [ 0:0]                      I16c7f1b874b0d05c6d120bbede254416;
reg  [MAX_SUM_WDTH_L-1:0]        I3740b30d31f3c61d93a14a46e3199c4d;
wire  [MAX_SUM_WDTH_L-1:0]       I3fd38a71ce6aa3db1d7a5a9f8a991e12;
wire  [MAX_SUM_WDTH_L-1:0]       I63e5718bf7d8771ef90b91be73d73264;
wire  [MAX_SUM_WDTH_L-1:0]       Ie385e1aeb2b0dcf6d2454be3d7708b27;
wire  [MAX_SUM_WDTH_L-1:0]       Ib2d1b7e105b25b492b45da72536d7578;
wire  [MAX_SUM_WDTH_L-1:0]       I588abf5ef4c583f0fec422736a0ce6a0;
wire  [MAX_SUM_WDTH_L-1:0]       I58bb95c56c7be17c263a2161210d7d8d;
wire  [MAX_SUM_WDTH_L-1:0]       Ifaf0e1f21b3bd7393c475b5126540a72;
wire  [MAX_SUM_WDTH_L-1:0]       I7027db9e0450724a6d417d708f1043f2;
reg  [ 0:0]                      I0c3cb2de514ecab0dd311e86a4dc3cdb;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf0a30abfec9031737eada436ac1a0d4;
wire  [MAX_SUM_WDTH_L-1:0]       Iebcb7206d8860b5094459c5d10b4efed;
wire  [MAX_SUM_WDTH_L-1:0]       I6bbf2b47a7dc50e66a3d8d258d6e31fb;
wire  [MAX_SUM_WDTH_L-1:0]       I8459abaa907f5afcd11884b1ec8c06c5;
wire  [MAX_SUM_WDTH_L-1:0]       Ia16ae2f6ef5000d47b6b84ed058252aa;
wire  [MAX_SUM_WDTH_L-1:0]       Ica32690dbc9ea110fefdce92260b125c;
wire  [MAX_SUM_WDTH_L-1:0]       Ic431d9383cce30b1889c92e2be4cb9d0;
wire  [MAX_SUM_WDTH_L-1:0]       Ib9cca4c0e58373c26d5fd9f51f793898;
wire  [MAX_SUM_WDTH_L-1:0]       I99bf0bc8ac20832b3724b2753f6ca449;
wire  [MAX_SUM_WDTH_L-1:0]       Ie701008f3c60c51ed72c5f964a8fc36e;
wire  [MAX_SUM_WDTH_L-1:0]       I3e2d78f8307a1787f8b2eccba94c7557;
reg  [ 0:0]                      Icc5ba4554d7a44bc3b43377efbe3b5f8;
reg  [MAX_SUM_WDTH_L-1:0]        Id36e8953a02400a5ab1f4dfdb0422e6d;
wire  [MAX_SUM_WDTH_L-1:0]       Ic1b4444ab0df9745d29bf893d9b83168;
wire  [MAX_SUM_WDTH_L-1:0]       I5f52dbf600656a8f5dc6b6b8a45ccebe;
wire  [MAX_SUM_WDTH_L-1:0]       I7f307af79f45ad4b9511e3961c917078;
wire  [MAX_SUM_WDTH_L-1:0]       Ie17a5be2a16d2efb98c976d7ee882535;
wire  [MAX_SUM_WDTH_L-1:0]       I5f19d2adff2f34a4bebe03f929a09c49;
wire  [MAX_SUM_WDTH_L-1:0]       I3cd69aeed9e869a2096d6dced5c209a0;
wire  [MAX_SUM_WDTH_L-1:0]       I359b6a22c9568a13b81670c741281393;
wire  [MAX_SUM_WDTH_L-1:0]       I24ba99614df383c38bbac50ae8b4487e;
wire  [MAX_SUM_WDTH_L-1:0]       I7498bee46de6b1c946ce95fdcc89f6e5;
wire  [MAX_SUM_WDTH_L-1:0]       I0f644f42cabf871b71e5a82871bc7b5d;
reg  [ 0:0]                      I5e51f49adb6dce65a9f19ff736526c4b;
reg  [MAX_SUM_WDTH_L-1:0]        Ica71108a53bfcfd1892b4d03ef68110c;
wire  [MAX_SUM_WDTH_L-1:0]       I71f9e059726a6cac8bdf0efcc0eadd2b;
wire  [MAX_SUM_WDTH_L-1:0]       I0c9b2c1da30bfab514bbb556ae7bd4c4;
wire  [MAX_SUM_WDTH_L-1:0]       I7918b2e37e96aee94fbccca7e0f75fc4;
wire  [MAX_SUM_WDTH_L-1:0]       I76eebd77eb77e0abcbc727d2c511370a;
wire  [MAX_SUM_WDTH_L-1:0]       Ibb2288e62110bae5b2d3fe901974e5c7;
wire  [MAX_SUM_WDTH_L-1:0]       I080f931dfef9d8adfb1dc1ee073eb64c;
wire  [MAX_SUM_WDTH_L-1:0]       Ide1106431e3565158bd81ccd6b18f3a1;
wire  [MAX_SUM_WDTH_L-1:0]       I63df19931e8d28666cccd79922cbd418;
wire  [MAX_SUM_WDTH_L-1:0]       I9a7e4a59447048de90446f877eb06627;
wire  [MAX_SUM_WDTH_L-1:0]       I0917e92ed84363ca92fd2074acd74eba;
reg  [ 0:0]                      Id57092394c7cda397f42374df4aa3fec;
reg  [MAX_SUM_WDTH_L-1:0]        I7c97629ec6e594f9b2160815ddd133cc;
wire  [MAX_SUM_WDTH_L-1:0]       Ie3eefdf7b5561a90a6ddd9e6aa432509;
wire  [MAX_SUM_WDTH_L-1:0]       I56eeb10d11e886cff629457a640a1c76;
wire  [MAX_SUM_WDTH_L-1:0]       I7a9eea89c4e76d856df44b6bdc332840;
wire  [MAX_SUM_WDTH_L-1:0]       If8d8f4333e893788fcb9ec54256e5b7a;
wire  [MAX_SUM_WDTH_L-1:0]       Ie4af0e7e04778d85f5dee73da33376a8;
wire  [MAX_SUM_WDTH_L-1:0]       I019a4e997adf54f5f5ca651f80b7901b;
wire  [MAX_SUM_WDTH_L-1:0]       I10294667f09abbfd4e2f757c414072fc;
wire  [MAX_SUM_WDTH_L-1:0]       Id4e8ab8f15b36bd27d1e4ebc5cbe1495;
wire  [MAX_SUM_WDTH_L-1:0]       I6c93588ca9e7c623d75314da39e89a91;
wire  [MAX_SUM_WDTH_L-1:0]       I1020412efc78d12a9ebcbaeb83e5dcea;
reg  [ 0:0]                      Idd6a4f8ae94c431f2fa3312b4fd287ba;
reg  [MAX_SUM_WDTH_L-1:0]        I4823c8239ace86dc399e906c1b5a0d74;
wire  [MAX_SUM_WDTH_L-1:0]       Id0b574f35a83dcfd4481a10043cd1884;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc577e5c2c7288373a8c5e3969ac1589;
wire  [MAX_SUM_WDTH_L-1:0]       Id18a1a17c1cf6e8a2492aa73b62898f2;
wire  [MAX_SUM_WDTH_L-1:0]       Id8ce8f636723b9f119bb86c25017e6b3;
reg  [ 0:0]                      I9f1f8590dcf596097bc81001d51684b9;
reg  [MAX_SUM_WDTH_L-1:0]        I10ad572ca72c2ea991487c39f7eabd7b;
wire  [MAX_SUM_WDTH_L-1:0]       Ic29a18d8d504a2d5280c1d7771346518;
wire  [MAX_SUM_WDTH_L-1:0]       I96a79193aa2956b8f901d5fcc9cf65cf;
wire  [MAX_SUM_WDTH_L-1:0]       I8c97a246c749fbef029f8b1671c772bd;
wire  [MAX_SUM_WDTH_L-1:0]       If9ba9d221909ce7499725f6fd7d519f8;
reg  [ 0:0]                      Icecd765baa87877675b0f3972d78c02f;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9f3fd3a6d16316e55addbe0e336519f;
wire  [MAX_SUM_WDTH_L-1:0]       I53a7878f44253f0f1a82d9d27b1a44c3;
wire  [MAX_SUM_WDTH_L-1:0]       Ie0e928125f9d3d17d123d97e00f1fc34;
wire  [MAX_SUM_WDTH_L-1:0]       I2bd0f77efeca09eebe82ea234e9fe638;
wire  [MAX_SUM_WDTH_L-1:0]       I94f2e7ef9b3463bd598dc9049f6fb0ef;
reg  [ 0:0]                      I401a38ea1d71dcc71d17a4694ceb0988;
reg  [MAX_SUM_WDTH_L-1:0]        I07965bca84276dd56da1af98e64b0adc;
wire  [MAX_SUM_WDTH_L-1:0]       I6dc16510af6b61b79b339d0fce77ac24;
wire  [MAX_SUM_WDTH_L-1:0]       Ic655e213ab81f5d61a018d3ed7016b12;
wire  [MAX_SUM_WDTH_L-1:0]       I2ffc4a604025a2f5c4e273c1d070a725;
wire  [MAX_SUM_WDTH_L-1:0]       I1c76818a9a3b688ca897aa479f7d807f;
reg  [ 0:0]                      I3db9b61e28a51e974e2d5e323ad53c1e;
reg  [MAX_SUM_WDTH_L-1:0]        Ic2ade31b8bcf68c4dcc1a371ff14074b;
wire  [MAX_SUM_WDTH_L-1:0]       I3bfee9d3d88f0569010a4e0101200c19;
wire  [MAX_SUM_WDTH_L-1:0]       I5d4738755a26beb6d0f61dd3dec0f804;
wire  [MAX_SUM_WDTH_L-1:0]       I2f3c800091275bcb72d1a2a38fba53f3;
wire  [MAX_SUM_WDTH_L-1:0]       I378e67cca7c4ff6325683f8346963210;
wire  [MAX_SUM_WDTH_L-1:0]       I04c8915a7f4bbde003f7facc84435c1a;
wire  [MAX_SUM_WDTH_L-1:0]       I3f50b10072f38b6addee6845e6df9118;
reg  [ 0:0]                      I96d0a4387f9b959bc779ac13351182cc;
reg  [MAX_SUM_WDTH_L-1:0]        Ic0edcf240048fbfde4e938c3e4c5e281;
wire  [MAX_SUM_WDTH_L-1:0]       Icc60eb18ba740036d2a17f98f15cfb98;
wire  [MAX_SUM_WDTH_L-1:0]       I1677daa18aa8b226753b1a887b9420d1;
wire  [MAX_SUM_WDTH_L-1:0]       I36bc2d4c9a4480daa9b0944c08b50738;
wire  [MAX_SUM_WDTH_L-1:0]       I38419a6905f50135a6783aacca0384dd;
wire  [MAX_SUM_WDTH_L-1:0]       Ib48892dcb0715987289662a14672611e;
wire  [MAX_SUM_WDTH_L-1:0]       Icd9c94f929dbc71c9b836fda3019630b;
reg  [ 0:0]                      I64082bc75fdbeb69a52a4361ed2d5883;
reg  [MAX_SUM_WDTH_L-1:0]        I8b42e89ff5f780d4ef8cd1cd5c99ef61;
wire  [MAX_SUM_WDTH_L-1:0]       I5d0249d9a772805b3fba3f3c7f5d35bd;
wire  [MAX_SUM_WDTH_L-1:0]       Ie97341deb6fb24d49eb8b96bd0fd3f35;
wire  [MAX_SUM_WDTH_L-1:0]       I17dd788f9d8e91307b6b1ab7488f9ce2;
wire  [MAX_SUM_WDTH_L-1:0]       I92ae370022ed107b152b10fd0aa3d2b7;
wire  [MAX_SUM_WDTH_L-1:0]       Iebb39f0d19ec1208bbfba6cf67a3bfc7;
wire  [MAX_SUM_WDTH_L-1:0]       I81861f6bb8bbbab6e93407cfb4a852b8;
reg  [ 0:0]                      I62929057b7c214bd38fd532e20ba5623;
reg  [MAX_SUM_WDTH_L-1:0]        I70b1b8521b36920707e95fc9418eb8a9;
wire  [MAX_SUM_WDTH_L-1:0]       I217b2e3ca0a534fc5b1910adf3c1b57d;
wire  [MAX_SUM_WDTH_L-1:0]       I8429b08891dc56af24c72ce1b7725457;
wire  [MAX_SUM_WDTH_L-1:0]       If96747262303f6c5c6b129e39224bd23;
wire  [MAX_SUM_WDTH_L-1:0]       If7012457af15c405baeaa1710319b541;
wire  [MAX_SUM_WDTH_L-1:0]       Ia0a0229ef71b85195352bb664ea4e4e3;
wire  [MAX_SUM_WDTH_L-1:0]       I42aeb7c23accc2ca874c7f8221c3af93;
reg  [ 0:0]                      I641179f37fef63e7deec603b3291381c;
reg  [MAX_SUM_WDTH_L-1:0]        I4fb1c32a62cbbaeb585c6564a3c938f9;
wire  [MAX_SUM_WDTH_L-1:0]       I7df6a95bf51f40693c439c6df36510d4;
wire  [MAX_SUM_WDTH_L-1:0]       I8fe65f9c344d7ec8657f192abefc3fb6;
wire  [MAX_SUM_WDTH_L-1:0]       I4d75c95d34d8d8aeeb528456bbe136e1;
wire  [MAX_SUM_WDTH_L-1:0]       I43746054a38c9521f8da9db9d0e91f99;
wire  [MAX_SUM_WDTH_L-1:0]       I0430ac2a4b2b2e2fc7f8154bf946553c;
wire  [MAX_SUM_WDTH_L-1:0]       I25dc807fd55b81c9f24fd0d1edcaa758;
reg  [ 0:0]                      Iff04b7ec87148f5bd408b4ec4b0590a5;
reg  [MAX_SUM_WDTH_L-1:0]        Iefc37daeec14e14ef2fe0716f73109dc;
wire  [MAX_SUM_WDTH_L-1:0]       I7881184f1779b9fd4fdf329c5f7664da;
wire  [MAX_SUM_WDTH_L-1:0]       I8e6de2d692a307ee8a5a4b2a9265a633;
wire  [MAX_SUM_WDTH_L-1:0]       I54b2b18ab051b468808a3d0fc4bc893f;
wire  [MAX_SUM_WDTH_L-1:0]       I37ee86e2ca32832862cb57efe76bbedf;
wire  [MAX_SUM_WDTH_L-1:0]       Ic95f2fc697574803c0f7fa35c2609f0c;
wire  [MAX_SUM_WDTH_L-1:0]       I933a30c52c9bec5172530b2d739a3b63;
reg  [ 0:0]                      I198bfb18d6f91c8f62777e6f592a88fa;
reg  [MAX_SUM_WDTH_L-1:0]        Ibd15f164f6d2ac9e5721a21464bc2c5c;
wire  [MAX_SUM_WDTH_L-1:0]       I7bbd7df18f85197c22fe8cfe37312af6;
wire  [MAX_SUM_WDTH_L-1:0]       I50d5ada7c91c7af16492c6b41151b68f;
wire  [MAX_SUM_WDTH_L-1:0]       I32c8e7996b3473d4906c40018799a16b;
wire  [MAX_SUM_WDTH_L-1:0]       Ic0eacd5a4812ad7ae3fa251ab2db4694;
wire  [MAX_SUM_WDTH_L-1:0]       Ideecf8ab87d28a840cd93851169ab05b;
wire  [MAX_SUM_WDTH_L-1:0]       I1ac6775eb38457b7962241d2e7336b0d;
reg  [ 0:0]                      Ia1562c88b4f56d8935c3a5d6ead0f816;
reg  [MAX_SUM_WDTH_L-1:0]        I951dfff9507bb70214d48e03a0ebb3a7;
wire  [MAX_SUM_WDTH_L-1:0]       I2ecaa89698604fddd863d7e28d643a57;
wire  [MAX_SUM_WDTH_L-1:0]       I273e0fe9c51c8549c8dfff393ca2e4e1;
wire  [MAX_SUM_WDTH_L-1:0]       Ifb1fc76002f6920a1f44c7b1bbcd0020;
wire  [MAX_SUM_WDTH_L-1:0]       Idf6d4e3aa753aa396a9bffb27732f851;
wire  [MAX_SUM_WDTH_L-1:0]       If14ca1f5d1c2977f9da79eaebaad1bf9;
wire  [MAX_SUM_WDTH_L-1:0]       If8f1505d9f10e30bd3320f500d34932f;
reg  [ 0:0]                      Iaccba3030d9d9f8a56f86d6e34ed6325;
reg  [MAX_SUM_WDTH_L-1:0]        Ie78e30b2a2eda75d0df7d10fd67b5e36;
wire  [MAX_SUM_WDTH_L-1:0]       Id32aa77c6406b35a00168bb5452b12fb;
wire  [MAX_SUM_WDTH_L-1:0]       I9a73686acefeb361337511f6943b036b;
wire  [MAX_SUM_WDTH_L-1:0]       Ib6eb7ce5a070f3a87bcf0e18be8c855d;
wire  [MAX_SUM_WDTH_L-1:0]       If69b0b717c35d33fc8c0e59b07eb9edc;
wire  [MAX_SUM_WDTH_L-1:0]       Ibb0d73078b779585e6b0e228391ecb96;
wire  [MAX_SUM_WDTH_L-1:0]       I2894546e399fe3e33d7579772a1310df;
reg  [ 0:0]                      I953dfeeacee8c44c08d0a425fa549e49;
reg  [MAX_SUM_WDTH_L-1:0]        Ia0b83a372dd4115dc4d61eb8ff0811b9;
wire  [MAX_SUM_WDTH_L-1:0]       I97f99a266267859aed199b278a430417;
wire  [MAX_SUM_WDTH_L-1:0]       Ie18cc792329941a3654322376a937d8d;
wire  [MAX_SUM_WDTH_L-1:0]       Ie914a99f08d60b74c3c36a632a4ca9b0;
wire  [MAX_SUM_WDTH_L-1:0]       I82916e9dc3894ad88e12de01a68d6aa5;
wire  [MAX_SUM_WDTH_L-1:0]       I6cbf576b3d652e34c0221f8316b5a392;
wire  [MAX_SUM_WDTH_L-1:0]       I9141b2516d7f855cd186472780af7b67;
reg  [ 0:0]                      I214a50bf9f879fe747904f4679fdd1f6;
reg  [MAX_SUM_WDTH_L-1:0]        If5c5bcbbea01aa22f242b913f0d01929;
wire  [MAX_SUM_WDTH_L-1:0]       I07bf32ed72de9c02abf700c64853af61;
wire  [MAX_SUM_WDTH_L-1:0]       I52663a2999fb9571834d517538691b6f;
wire  [MAX_SUM_WDTH_L-1:0]       I8dcb88c94506367aabe8d7ed62cc56c2;
wire  [MAX_SUM_WDTH_L-1:0]       Ie676a4bee61154145391d9cc473fe91d;
wire  [MAX_SUM_WDTH_L-1:0]       I9502c8fbf6b48749bf9f84a89a937dfe;
wire  [MAX_SUM_WDTH_L-1:0]       I0c91e540e7106f32ae59491d8ed1853e;
reg  [ 0:0]                      Ic88f2c344a8ad254fc7d7034cb594f6d;
reg  [MAX_SUM_WDTH_L-1:0]        Iccba58cd3519fb4cc75a61b50da1d562;
wire  [MAX_SUM_WDTH_L-1:0]       Iddfb8a8e261389eb4a2a10880c19446a;
wire  [MAX_SUM_WDTH_L-1:0]       If0d55f861d4b3f0970c529024ca142d5;
wire  [MAX_SUM_WDTH_L-1:0]       Ib054f5d3f5cbb29a053d0e50c23cb3a8;
wire  [MAX_SUM_WDTH_L-1:0]       I1d65e9f97e93de8cc2a5dd532f8e482a;
wire  [MAX_SUM_WDTH_L-1:0]       I3bdeab8c87325d46e45d9e2d44756934;
wire  [MAX_SUM_WDTH_L-1:0]       If9228f7ecf19c41f4bbd8dabd0d5816c;
reg  [ 0:0]                      If299d1a4e044acbc70bc3b7bce9f86e9;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc0999e4d0b3cc2650f9348b8c204b14;
wire  [MAX_SUM_WDTH_L-1:0]       I9e3edee214c4937d2aa462d3cffa624b;
wire  [MAX_SUM_WDTH_L-1:0]       I9fcbbd2e81b006b50e2d35ed2627bf83;
wire  [MAX_SUM_WDTH_L-1:0]       Ie16f3d50ad5e5581ca099549db7232d2;
wire  [MAX_SUM_WDTH_L-1:0]       I6345e93f3fa7f5eb2008dd41742afc2d;
reg  [ 0:0]                      Idb373d2cf788f6a93a0e5df7f9179292;
reg  [MAX_SUM_WDTH_L-1:0]        I2aeff1fb4b839a581acaf26f90f9113c;
wire  [MAX_SUM_WDTH_L-1:0]       I698b93e10073b5d29357cde4bcac9dbe;
wire  [MAX_SUM_WDTH_L-1:0]       Ie7ced910d84655790823e6173a5a314a;
wire  [MAX_SUM_WDTH_L-1:0]       If6e3b6fd1810f6964e9024329d7cb3e3;
wire  [MAX_SUM_WDTH_L-1:0]       If1045908c6d7476bd5507e57d08c406c;
reg  [ 0:0]                      Ic73b8c8f76a985330d4ac1fa0cc28e7f;
reg  [MAX_SUM_WDTH_L-1:0]        I7d60d53f883f8187700c4e78b4c22f1c;
wire  [MAX_SUM_WDTH_L-1:0]       I4d4f6705ed77a16ff31b34bae0d8b6d9;
wire  [MAX_SUM_WDTH_L-1:0]       I70a492396580ac1143d8a2f4b181e873;
wire  [MAX_SUM_WDTH_L-1:0]       I2fade32b5bdf245fa15289620dae2670;
wire  [MAX_SUM_WDTH_L-1:0]       Ie0dc166f57fea074496241a32cdb6015;
reg  [ 0:0]                      I134dfb2c57d8cdffd2789e2f442c3247;
reg  [MAX_SUM_WDTH_L-1:0]        Id6fcf4b7af4a37c854a12e2ae80851fa;
wire  [MAX_SUM_WDTH_L-1:0]       If6a2518891412caa6d6d507082501f1e;
wire  [MAX_SUM_WDTH_L-1:0]       Ic9912e5a838a377b26a19d22148a64df;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc0fca22d16444bc17877106ca772c31;
wire  [MAX_SUM_WDTH_L-1:0]       Ie4291d233597d5d676a80fd62d9bd208;
reg  [ 0:0]                      I0c735e43be8030078ec10bdb6882e79c;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa5e5f7d753964f14f0f16dbe552fd85;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc13b798d76aa70ec1877c275fb31d36;
wire  [MAX_SUM_WDTH_L-1:0]       I57d6637f0bdab578a790e4a12ccaa16b;
wire  [MAX_SUM_WDTH_L-1:0]       If8ea04fe685b4f20cdaf9a84984d56fe;
wire  [MAX_SUM_WDTH_L-1:0]       Ie0c86f20c28bcbe410b191b90d29bf76;
wire  [MAX_SUM_WDTH_L-1:0]       I3dc5d3f66726e15968a70cbf3d3b656a;
reg  [ 0:0]                      Ie9951415c1d599570af1787767caa2dc;
reg  [MAX_SUM_WDTH_L-1:0]        I900d471b087cf5a436c2ad66a84d8280;
wire  [MAX_SUM_WDTH_L-1:0]       Id674686e7ac37fd6f63846f9a9cede19;
wire  [MAX_SUM_WDTH_L-1:0]       Ie2ed9668d13d219c60f2e0614488cd42;
wire  [MAX_SUM_WDTH_L-1:0]       I98abc995ff89934534543be93c6e3ffa;
wire  [MAX_SUM_WDTH_L-1:0]       I579cf9386ab7b08efa204d735335e462;
wire  [MAX_SUM_WDTH_L-1:0]       I9efa4d729d10a6b7cc335fb765ed032c;
reg  [ 0:0]                      I2630f187d63ba9b0af52c77093e6b760;
reg  [MAX_SUM_WDTH_L-1:0]        I6d1434907f0292ea2ee47cbc5b52bfb9;
wire  [MAX_SUM_WDTH_L-1:0]       If9191ebc8e88d4e75f0f35897ebb1421;
wire  [MAX_SUM_WDTH_L-1:0]       I3511287cfe69d5cedc5a8fbcad708437;
wire  [MAX_SUM_WDTH_L-1:0]       I91812179d44cb675b90d477f33ec48ad;
wire  [MAX_SUM_WDTH_L-1:0]       Idb04a1aae91fdc477ca38ed66789ee88;
wire  [MAX_SUM_WDTH_L-1:0]       I566054aece562960590ee28b157e4a3e;
reg  [ 0:0]                      I83db667ace2f04ef4950e2c186e0e6a4;
reg  [MAX_SUM_WDTH_L-1:0]        I938bef7ba7ae1739d8e6a6a7c117a1b1;
wire  [MAX_SUM_WDTH_L-1:0]       I7b2ffb762cd9ef7aa8ba224efb75c46c;
wire  [MAX_SUM_WDTH_L-1:0]       Id90bbb642b0f4434d8a148a28b6b2f65;
wire  [MAX_SUM_WDTH_L-1:0]       Ia4e297e35d484b15adce7e1d67f582b0;
wire  [MAX_SUM_WDTH_L-1:0]       I84996b1d03b692f6f736fb04c7f91e83;
wire  [MAX_SUM_WDTH_L-1:0]       I83078cc7857fc17b30f640854a4d6be5;
reg  [ 0:0]                      Ie818c5ea3f3b879fded32e6cb06ca546;
reg  [MAX_SUM_WDTH_L-1:0]        I6384a9416b2d1da01df1b2d7b16c5390;
wire  [MAX_SUM_WDTH_L-1:0]       I94bb467129904032736fb13dd636c600;
wire  [MAX_SUM_WDTH_L-1:0]       Ifa76758b50f439170ecd6d86ff898bc4;
wire  [MAX_SUM_WDTH_L-1:0]       I9d831dd976e8cd5d8f6a6818601e6424;
wire  [MAX_SUM_WDTH_L-1:0]       I474774ae149804412ed4aaf1cdcaba88;
wire  [MAX_SUM_WDTH_L-1:0]       I964cdcb4e6b49a62d30c2a2540851317;
reg  [ 0:0]                      I3a67a175863091a52844aae6ad277da0;
reg  [MAX_SUM_WDTH_L-1:0]        I5097a79e7cf7a30d38ba198d1407119c;
wire  [MAX_SUM_WDTH_L-1:0]       I6df268bc9f85ce88674a9165664ea84a;
wire  [MAX_SUM_WDTH_L-1:0]       I74fdcbe9f49f7bce1f5e31d956c5883c;
wire  [MAX_SUM_WDTH_L-1:0]       I4a1b8453cb7a21745d5f74ad05653ed2;
wire  [MAX_SUM_WDTH_L-1:0]       I9c53b478b2011fac0615a152fe60d5b6;
wire  [MAX_SUM_WDTH_L-1:0]       Id75dbed8f1a5befda32c60b994681013;
reg  [ 0:0]                      Ia3aba80aead67feab12e4800fef82322;
reg  [MAX_SUM_WDTH_L-1:0]        Ib113c26c8dcf49c972c41a938059a787;
wire  [MAX_SUM_WDTH_L-1:0]       I378a59323b74623c5524f854d6e11226;
wire  [MAX_SUM_WDTH_L-1:0]       I080bf885464a0cc948a4450e9f7d1d26;
wire  [MAX_SUM_WDTH_L-1:0]       If769e73adea227de1fd85c2e89d0ba08;
wire  [MAX_SUM_WDTH_L-1:0]       Ifa6a34b83225e9d9b28b14874c4444e3;
wire  [MAX_SUM_WDTH_L-1:0]       I584b1d4d6fb7ee4f20ad9c96715cdf90;
reg  [ 0:0]                      I1181d42b560fca7bb5c924a81a5db1fc;
reg  [MAX_SUM_WDTH_L-1:0]        I970c4a25a8bce82a9d2846679029fcab;
wire  [MAX_SUM_WDTH_L-1:0]       I265f9b91fbb62164e589dcf96818c4f5;
wire  [MAX_SUM_WDTH_L-1:0]       I3d59a47c88227734cf6fc0d6fd30db11;
wire  [MAX_SUM_WDTH_L-1:0]       I6144b6df2c87ea0948d730343b42129f;
wire  [MAX_SUM_WDTH_L-1:0]       Ia7ca7400e36ea572fba8e19bcc81ecbd;
wire  [MAX_SUM_WDTH_L-1:0]       I302e61b49accf5db556b87517f2341f5;
reg  [ 0:0]                      Ie4e5f3d7c5d2df30653f5666d14567bf;
reg  [MAX_SUM_WDTH_L-1:0]        Ibe2af096ad2db26e54d8b4b3bb05175c;
wire  [MAX_SUM_WDTH_L-1:0]       I5d9af1abff6efe3a55c6568d936b6ec7;
wire  [MAX_SUM_WDTH_L-1:0]       I8cde0aa611c476b5112edeb8f17f15bf;
wire  [MAX_SUM_WDTH_L-1:0]       Icaa40ec40d6d26cdf70bb5ae7d492e47;
wire  [MAX_SUM_WDTH_L-1:0]       I8346f15d822cacfeecbe5d75412cb53f;
wire  [MAX_SUM_WDTH_L-1:0]       I5ee364aab320ab40c0f65feda6f53b18;
reg  [ 0:0]                      Ifd9345cf219c58291c0b437aac093d78;
reg  [MAX_SUM_WDTH_L-1:0]        Ie48569c467fba0c1291f71d6080ebedc;
wire  [MAX_SUM_WDTH_L-1:0]       I1f0ecba054900f96cd7100741191c5f4;
wire  [MAX_SUM_WDTH_L-1:0]       I4faf2caf62966416118a54015908c889;
wire  [MAX_SUM_WDTH_L-1:0]       Idd0329980a36f87859150530ab44b52d;
wire  [MAX_SUM_WDTH_L-1:0]       Ie66bc10dde27f08813d4d347fd7cf6ce;
wire  [MAX_SUM_WDTH_L-1:0]       Ie1d8b3ea7c6603cebf2f9adb776910b7;
reg  [ 0:0]                      I4f2d7bb48918ce51efe6b3b12f9f8e65;
reg  [MAX_SUM_WDTH_L-1:0]        I90e7ded06617b49cdb8b5301fe9c6a20;
wire  [MAX_SUM_WDTH_L-1:0]       Ia37488e9a50cf5cc08de74ade676db96;
wire  [MAX_SUM_WDTH_L-1:0]       I08aa45211cab01d567cd5eb172fd2f0c;
wire  [MAX_SUM_WDTH_L-1:0]       If4ff0c63ec1deb46412858e496451a01;
wire  [MAX_SUM_WDTH_L-1:0]       Ife7bfd15fc4c392b5d2288d9a4e879b3;
wire  [MAX_SUM_WDTH_L-1:0]       I24ac26debafd03c7333d174e8725afd6;
reg  [ 0:0]                      Ifa612e6208151c616c3a0319182a96f1;
reg  [MAX_SUM_WDTH_L-1:0]        I4920014f5d017f4e840dc3b88526955f;
wire  [MAX_SUM_WDTH_L-1:0]       I99d80ad68e2563d0f78a0e3bb82c5328;
wire  [MAX_SUM_WDTH_L-1:0]       I9943733ef305983c629565c881054bbf;
wire  [MAX_SUM_WDTH_L-1:0]       I7cb4420bc55c03a6500f5228d31fe43c;
wire  [MAX_SUM_WDTH_L-1:0]       Ic4d19dec464359c0a9fa75148fe90c73;
wire  [MAX_SUM_WDTH_L-1:0]       I44993416e1d22613dbd78402c37a934d;
reg  [ 0:0]                      I9cb28a0cc6358610854c8f8d1dd3c707;
reg  [MAX_SUM_WDTH_L-1:0]        I03b70553f1c501609400574ae7cd73f5;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc9b94a9dea471805cb442ac6904bc97;
wire  [MAX_SUM_WDTH_L-1:0]       I917d9f9b144d3bffafc77bddae7fba6b;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc91c6c3d56bb8a14e22909c43ffec51;
wire  [MAX_SUM_WDTH_L-1:0]       If7c2d3eddd96b47b6c2aea8b27c8c7f4;
reg  [ 0:0]                      I40bcc924f5cf1f7d587aa35267022261;
reg  [MAX_SUM_WDTH_L-1:0]        I63c9bf68b43ed66c51b0f4c0ed92e9ab;
wire  [MAX_SUM_WDTH_L-1:0]       I4df093ed94d26b058e97db550e347e3c;
wire  [MAX_SUM_WDTH_L-1:0]       Ie90303b0326bee4ab203a8cf1e643da9;
wire  [MAX_SUM_WDTH_L-1:0]       I19030d352fd059156ee42c66f9270beb;
wire  [MAX_SUM_WDTH_L-1:0]       I36767a902c53a384128ae1443cf88963;
reg  [ 0:0]                      I5238f7273b05b8b9f376314acdc6cc42;
reg  [MAX_SUM_WDTH_L-1:0]        If408dfead07757878cc878131bc7d6a3;
wire  [MAX_SUM_WDTH_L-1:0]       I868dffa3f07407f7996bb5bc596939b7;
wire  [MAX_SUM_WDTH_L-1:0]       I7d928be164d0dce8b1322ff230c053e9;
wire  [MAX_SUM_WDTH_L-1:0]       I98be4971a8a9a08abb3ebe474d7f0c6d;
wire  [MAX_SUM_WDTH_L-1:0]       I779e70dea33201e9237f29681ffd5e27;
reg  [ 0:0]                      I7137f56eeb4c4ae08bbc238db4cd3441;
reg  [MAX_SUM_WDTH_L-1:0]        Ia0857d63d309807789b6ff4f6028f1b3;
wire  [MAX_SUM_WDTH_L-1:0]       Ie2262914042172ab7e08599278f36af5;
wire  [MAX_SUM_WDTH_L-1:0]       I4001323da8f7956cdd480ac2d56df929;
wire  [MAX_SUM_WDTH_L-1:0]       Ib1cd6731034887a0a55e405c9db3e8de;
wire  [MAX_SUM_WDTH_L-1:0]       I51aa496e8c03944c28a908102514e6f8;
reg  [ 0:0]                      I02335be013799e2560a98b6a82a0c528;
reg  [MAX_SUM_WDTH_L-1:0]        I53921b825c5e434b63bee0e1ecb7a517;
wire  [MAX_SUM_WDTH_L-1:0]       I6415f3996318472532e161510ccc8ca3;
wire  [MAX_SUM_WDTH_L-1:0]       Ia11b671b59240988737979328c472812;
wire  [MAX_SUM_WDTH_L-1:0]       Id4fabe0165a117a402dc14f2f3ec626a;
wire  [MAX_SUM_WDTH_L-1:0]       I57238f501ab7278b308d76211ced8cf7;
wire  [MAX_SUM_WDTH_L-1:0]       I9b257f8556ca4e5402637f01081b78e1;
reg  [ 0:0]                      Id327bb65156c8307901dfcb4184bb65f;
reg  [MAX_SUM_WDTH_L-1:0]        I5e68f84e123c37f19a03c13892c77e19;
wire  [MAX_SUM_WDTH_L-1:0]       I2e093412a9fa3972cea01664389d8c27;
wire  [MAX_SUM_WDTH_L-1:0]       I17907fd8c6975c8c642535ff929221a6;
wire  [MAX_SUM_WDTH_L-1:0]       I3c6577b04ad56d864bbaa2c048323c11;
wire  [MAX_SUM_WDTH_L-1:0]       I6f0c341c05eaa8f35bbce4521f6e8f94;
wire  [MAX_SUM_WDTH_L-1:0]       Ib72ba950ecf9ae2668374f6633a67ca7;
reg  [ 0:0]                      I56331cb7b310613016958553732cdf40;
reg  [MAX_SUM_WDTH_L-1:0]        Id5270b57c6fb4b18db3bbd0a523e467e;
wire  [MAX_SUM_WDTH_L-1:0]       I3d7c72d725f4563bb562e2992093cb02;
wire  [MAX_SUM_WDTH_L-1:0]       I813c881ac61a59041be3be78f6a466c8;
wire  [MAX_SUM_WDTH_L-1:0]       I866510e7dc721fa5aac312bc5ab5ba0a;
wire  [MAX_SUM_WDTH_L-1:0]       Ib4432359f97849dff6ad3e0f044157bd;
wire  [MAX_SUM_WDTH_L-1:0]       Ic86aa6eb1b4dcc2520309089b43292e6;
reg  [ 0:0]                      Ie3b00960f8af88a5aba7a2104dfca9a7;
reg  [MAX_SUM_WDTH_L-1:0]        I3c18a84617eb21472d53e598700d7f4c;
wire  [MAX_SUM_WDTH_L-1:0]       I0731115afe5c15bcf131f7ef4f05802b;
wire  [MAX_SUM_WDTH_L-1:0]       Ib080b8fd34385aa7986dace4afd95267;
wire  [MAX_SUM_WDTH_L-1:0]       I134890b77451d0b78afc7402a6a28048;
wire  [MAX_SUM_WDTH_L-1:0]       I956da75f13433c1dd7a3cbd3b78922c1;
wire  [MAX_SUM_WDTH_L-1:0]       I440b26c9f1b9ccf70f97c9d5f732d38e;
reg  [ 0:0]                      I7d1ef47f35b7a4c3ea2e4383732de398;
reg  [MAX_SUM_WDTH_L-1:0]        Id36663e7a01fff3170833ecfecac1321;
wire  [MAX_SUM_WDTH_L-1:0]       I5e3a441faca44bffc4368d96d8fb0bfd;
wire  [MAX_SUM_WDTH_L-1:0]       I21d7ba25247a87a1a9c245d0d1f553b0;
wire  [MAX_SUM_WDTH_L-1:0]       I55aafa8162cfc4fccfae68cf78cd1c2b;
wire  [MAX_SUM_WDTH_L-1:0]       Ib99c25f0d8d6493cac4d5c816884c704;
wire  [MAX_SUM_WDTH_L-1:0]       Iee7c9f0a0e8ca127efee008b4874edbd;
reg  [ 0:0]                      Ibb013f036fc42687a04bdcbe2d0bbd8a;
reg  [MAX_SUM_WDTH_L-1:0]        I8d3be15109c7007a79fecaac0d891626;
wire  [MAX_SUM_WDTH_L-1:0]       I17b4a3baae65161387f472037ffc6fc4;
wire  [MAX_SUM_WDTH_L-1:0]       Ie7b7b202a968fe73f6b1e02a044414c5;
wire  [MAX_SUM_WDTH_L-1:0]       I479ab5c0e483c36267d8248340006666;
wire  [MAX_SUM_WDTH_L-1:0]       I777bfe165e25d7fde4fc950f23db7b84;
wire  [MAX_SUM_WDTH_L-1:0]       I146d505a34ddb8d65e0a1769f623a7fd;
reg  [ 0:0]                      I77eae49d321f1d1e39dd7c75829aaedc;
reg  [MAX_SUM_WDTH_L-1:0]        I92169cc57291f20d336a479e392ec271;
wire  [MAX_SUM_WDTH_L-1:0]       Ia85239bddc04bf50bcf037ed2f76d7ac;
wire  [MAX_SUM_WDTH_L-1:0]       Ia7306bacf3c2b180d3261a5c1f0f4a30;
wire  [MAX_SUM_WDTH_L-1:0]       I2018147b86e47af5842c4f29d047d157;
wire  [MAX_SUM_WDTH_L-1:0]       Id17a85459845f8a8be694c4bf1fc29c9;
wire  [MAX_SUM_WDTH_L-1:0]       Ic012b15584d9d25af38f83d0526503da;
reg  [ 0:0]                      I420a4d69a077dc1996ddb4b715d63e15;
reg  [MAX_SUM_WDTH_L-1:0]        I6178b220b469b40dac39168057023a1c;
wire  [MAX_SUM_WDTH_L-1:0]       I7f09bd4a45143a036ce04af11b9927f9;
wire  [MAX_SUM_WDTH_L-1:0]       Ica32f94af6e6f3eaf2b724a2173fa463;
wire  [MAX_SUM_WDTH_L-1:0]       Ib750bb83ddfbbad2a2be8d1c8392b4ff;
wire  [MAX_SUM_WDTH_L-1:0]       I3906ece39480f96020717c6243e8ba4c;
wire  [MAX_SUM_WDTH_L-1:0]       Ie68ce21ade07fa53c30ebf27216b03f9;
reg  [ 0:0]                      I652202a4dc8f102d29334b4811f5628d;
reg  [MAX_SUM_WDTH_L-1:0]        I55342938216a0ea0889f96c2f6c05ce5;
wire  [MAX_SUM_WDTH_L-1:0]       I6cc6fa167c0d2b4b62ddbeecea175ed2;
wire  [MAX_SUM_WDTH_L-1:0]       Ibddf3468ae7c27d5a4b1388e524aa9c2;
wire  [MAX_SUM_WDTH_L-1:0]       Iadcb2b3acaac2e1bb505c65d3cbe4235;
wire  [MAX_SUM_WDTH_L-1:0]       I37cd96b8b0a4939d9a70098fd8bcf452;
reg  [ 0:0]                      I0e33e0cdf39fc4cc99f6696e9f2784de;
reg  [MAX_SUM_WDTH_L-1:0]        Idf28431c76a84a48dd895979d2b11a63;
wire  [MAX_SUM_WDTH_L-1:0]       Ib34b169dcc76daee2d1aa2b2a7513af3;
wire  [MAX_SUM_WDTH_L-1:0]       If36fc316d6ec7c7e09eae77807b37099;
wire  [MAX_SUM_WDTH_L-1:0]       Ifd214c332218ac5c0fe5aded4b952711;
wire  [MAX_SUM_WDTH_L-1:0]       Idcd0fc8f86e2b6f03606b818b8346e5a;
reg  [ 0:0]                      Ib9479328689dec62f900946e56ba0eb4;
reg  [MAX_SUM_WDTH_L-1:0]        I1ef61124c8d62e8f6a82a729fb091694;
wire  [MAX_SUM_WDTH_L-1:0]       If486aa8ac2cfb46f936714812cc760df;
wire  [MAX_SUM_WDTH_L-1:0]       I2d8e5b5fdbda7d599423c38aaace6658;
wire  [MAX_SUM_WDTH_L-1:0]       I6d0878fb7ec75c0a26be4dbba62f80dc;
wire  [MAX_SUM_WDTH_L-1:0]       I16a16ff0e8a6685a09803634da429fd2;
reg  [ 0:0]                      I2728682c0f749d1a9e8afeacdf44bfb7;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8bb96f0372323e6a8072ca56fb9396d;
wire  [MAX_SUM_WDTH_L-1:0]       Idb211abaa54ac26e7379c64a63f7d07c;
wire  [MAX_SUM_WDTH_L-1:0]       I351205eb71acb31b59d2b4470f0ba28c;
wire  [MAX_SUM_WDTH_L-1:0]       If5660c495bf7690252783d888d1ad6e8;
wire  [MAX_SUM_WDTH_L-1:0]       I3a5229cb8e44a15560b5c7bef96e65cc;
reg  [ 0:0]                      I07da3bb5f943db6271fe1867a358df35;
reg  [MAX_SUM_WDTH_L-1:0]        I432f74dda4f6b1cebdf5ad59c659080b;
wire  [MAX_SUM_WDTH_L-1:0]       I889b9b0828e97fe44d8366c5ef71a8f2;
wire  [MAX_SUM_WDTH_L-1:0]       Ie23062e00e39ead706f5b6ead233747d;
wire  [MAX_SUM_WDTH_L-1:0]       I8a2589544c75ecfdc31d28912c639695;
wire  [MAX_SUM_WDTH_L-1:0]       I5c21c59147e9c3a74c7cbbb6f2a23919;
wire  [MAX_SUM_WDTH_L-1:0]       Idacd78e24408e432abbbfb0c447fdde5;
reg  [ 0:0]                      I61fc44808c85a75909b9d9fd4035f147;
reg  [MAX_SUM_WDTH_L-1:0]        Idc689442305acd00f0f32416d8fb3773;
wire  [MAX_SUM_WDTH_L-1:0]       I0e8b171fe5080485a7f4fef83f1f1528;
wire  [MAX_SUM_WDTH_L-1:0]       Ib22c2bd76e6c29cc2f1440885bf24b7b;
wire  [MAX_SUM_WDTH_L-1:0]       I149559fccd9def4ec1ead1fdcff3c7fd;
wire  [MAX_SUM_WDTH_L-1:0]       Icfa8fed3239748abca27a5fc17de79c0;
wire  [MAX_SUM_WDTH_L-1:0]       I2ff115fa483f080d93bada49a9566b33;
reg  [ 0:0]                      Ic5075ee0ad355c20dd45ed594f2a8c3f;
reg  [MAX_SUM_WDTH_L-1:0]        Ida03738adc101c03c2229756bed2469d;
wire  [MAX_SUM_WDTH_L-1:0]       Ibee4f3cd2f516c29ab68e07a640ab65e;
wire  [MAX_SUM_WDTH_L-1:0]       Ie495ab560f59ad038992c573de7d2f5b;
wire  [MAX_SUM_WDTH_L-1:0]       Ibd812def78c3a9c02f9ba45cc0413711;
wire  [MAX_SUM_WDTH_L-1:0]       I98166634dc80201b0cefb01d9559c228;
wire  [MAX_SUM_WDTH_L-1:0]       Ic2f03a980b5f0b042853ca746abab22b;
reg  [ 0:0]                      Ic0a651f45a502ead495cf14f97d65bfc;
reg  [MAX_SUM_WDTH_L-1:0]        I4d14c75f28f3e516c259ea288996131b;
wire  [MAX_SUM_WDTH_L-1:0]       I2807a88097d2683ebdb9e0e785e3af02;
wire  [MAX_SUM_WDTH_L-1:0]       I8bebbb3a676c8506af0768516abcd740;
wire  [MAX_SUM_WDTH_L-1:0]       I31d380f34691c9fe9022035f233b77e2;
wire  [MAX_SUM_WDTH_L-1:0]       I1ffb5675c98ab5b3c62b24eb23441473;
wire  [MAX_SUM_WDTH_L-1:0]       If56424546ec4f3445853538207ea864e;
reg  [ 0:0]                      Ic1c05ea22f708f620f626cc8c5ca309c;
reg  [MAX_SUM_WDTH_L-1:0]        I6e6cbbf430d57f347a0d70558af143d8;
wire  [MAX_SUM_WDTH_L-1:0]       I31a49be4a34d9bac2e0d815097439772;
wire  [MAX_SUM_WDTH_L-1:0]       I6b96a2498078953e87de223aa2236d50;
wire  [MAX_SUM_WDTH_L-1:0]       I79bf36e298a85a42c7432f877055f0b4;
wire  [MAX_SUM_WDTH_L-1:0]       I90c070b9bde5da05e8a5d25d2de3ba6b;
wire  [MAX_SUM_WDTH_L-1:0]       I28d0e4e6d772dd58d845d91952ada300;
reg  [ 0:0]                      I61a18378aadae4556da501ce997321b4;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7487df45118e44acec6b9d07bbd5969;
wire  [MAX_SUM_WDTH_L-1:0]       I7232b4e277acc6f1acefcb606ca24508;
wire  [MAX_SUM_WDTH_L-1:0]       I32da124c433c55f692ffa4734d0dc8fc;
wire  [MAX_SUM_WDTH_L-1:0]       I56e487db14eeb8d93f494d2f11b57a49;
wire  [MAX_SUM_WDTH_L-1:0]       I94d3c02bd5b8e84926d4b3c2f56efeac;
wire  [MAX_SUM_WDTH_L-1:0]       I0c35b2e9176f9a06e26ca67d036411b4;
reg  [ 0:0]                      Ib1fc521709a1ce2198fd8df5b41d0177;
reg  [MAX_SUM_WDTH_L-1:0]        I492f382fea500462b3d0866240fb91b2;
wire  [MAX_SUM_WDTH_L-1:0]       Ia6ee7b70d0b7fe7c346760b1784e50b9;
wire  [MAX_SUM_WDTH_L-1:0]       I7ce57c278c683ad045526e49bcc47412;
wire  [MAX_SUM_WDTH_L-1:0]       Ie3d3e681cac0bb919946ac27057409e2;
wire  [MAX_SUM_WDTH_L-1:0]       I8ea0a8cdd6506c982ad75f23136bcebe;
wire  [MAX_SUM_WDTH_L-1:0]       Ic812f8bc775c5ee6a83e2b9aeb22b2a4;
reg  [ 0:0]                      I1bb5511c9cda1a595c45ecde48e9ebc7;
reg  [MAX_SUM_WDTH_L-1:0]        I3fb3ebddaf28efb56092d19a1b4695de;
wire  [MAX_SUM_WDTH_L-1:0]       I0f0adf7fe957b9a68772bd8a1bc163d4;
wire  [MAX_SUM_WDTH_L-1:0]       If09562f8d82bc1dea7c38ed51523a889;
wire  [MAX_SUM_WDTH_L-1:0]       Ib0fd21d66cd89c4e5c95fbc9c7680b62;
wire  [MAX_SUM_WDTH_L-1:0]       I5a2b2bfadc638fe3fdc31136a8f09a8d;
wire  [MAX_SUM_WDTH_L-1:0]       Ica914d8c556285d6b90b35747065a6e5;
reg  [ 0:0]                      I4a29c37ed36b6e12f1f8e263c92bdbc1;
reg  [MAX_SUM_WDTH_L-1:0]        I22a26b7f0b1c8c16b00597732ce2ab23;
wire  [MAX_SUM_WDTH_L-1:0]       I00c5d739bccb0ab6d05da70fe51aafea;
wire  [MAX_SUM_WDTH_L-1:0]       I18e448761bc014ce490b766183350312;
wire  [MAX_SUM_WDTH_L-1:0]       I1b5920f488e9469bd416a6af3072a30b;
wire  [MAX_SUM_WDTH_L-1:0]       I70b41ffed4b6d88ddff219c567b8e968;
reg  [ 0:0]                      I4bf02a07719402890405fb2e7b679ed9;
reg  [MAX_SUM_WDTH_L-1:0]        I2ac08a2d8c917ecb37fbaf5325cb0473;
wire  [MAX_SUM_WDTH_L-1:0]       I935e083b4561da7d015e98ca7f02854e;
wire  [MAX_SUM_WDTH_L-1:0]       Iaca9ef263bf220d786242b88c994fd21;
wire  [MAX_SUM_WDTH_L-1:0]       I92169291959eb33452b79bfd32618cbc;
wire  [MAX_SUM_WDTH_L-1:0]       I126dabc3ebb9c4157adf62b57f217bd0;
reg  [ 0:0]                      I75bd82990cb60b6d7ccd7aa2982da7aa;
reg  [MAX_SUM_WDTH_L-1:0]        I50ff8f51e75fb9ce3db983c2a0f57196;
wire  [MAX_SUM_WDTH_L-1:0]       If4433b1ef2eb963cd301946958b69884;
wire  [MAX_SUM_WDTH_L-1:0]       I67ac5b9b794787b3c4738c3366689871;
wire  [MAX_SUM_WDTH_L-1:0]       I4f022d70078c412bdbef158f750d3da3;
wire  [MAX_SUM_WDTH_L-1:0]       I6be6165385f6a77aeedb88f2baaa9cab;
reg  [ 0:0]                      Ia6d3e38249f8a1208540b68f54c46769;
reg  [MAX_SUM_WDTH_L-1:0]        I444bc340ffb7ef7b72d4d2e761d58872;
wire  [MAX_SUM_WDTH_L-1:0]       Id1f7fe91547e158e1d39edffb1421ff3;
wire  [MAX_SUM_WDTH_L-1:0]       I7a51924134902612db53941390891245;
wire  [MAX_SUM_WDTH_L-1:0]       I45128b9e29dd2fdd94a78fc5ffdff2b1;
wire  [MAX_SUM_WDTH_L-1:0]       I7f1082408c8ebb5be18e8f71ff9510e5;
reg  [ 0:0]                      Idf548b72357ab28fd956791e84e5d65c;
reg  [MAX_SUM_WDTH_L-1:0]        I039c6cac5830759529595a958b7f65c9;
wire  [MAX_SUM_WDTH_L-1:0]       I655ebf19c2f4b3dde716668f9ce12e59;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc9d493a507122d92af42d858cdc4c61;
wire  [MAX_SUM_WDTH_L-1:0]       Ib3d3103e5ee4feb160a97c7e26f7102b;
wire  [MAX_SUM_WDTH_L-1:0]       I6cc56b119e72175df3b7ce64dc3d9305;
reg  [ 0:0]                      I50b6f2e0ef2831535ac8c18cd7ca9379;
reg  [MAX_SUM_WDTH_L-1:0]        I0584de7d919236ab138e288a27d08ff1;
wire  [MAX_SUM_WDTH_L-1:0]       I57cf4a9378f1cdd94a1a5608dc57e05f;
wire  [MAX_SUM_WDTH_L-1:0]       I4160ab1aa18e8151c0a5c23b9edeb907;
wire  [MAX_SUM_WDTH_L-1:0]       Ia1f183f2d904d006e46399424e06c614;
wire  [MAX_SUM_WDTH_L-1:0]       If979702738671323995e56108bc9376c;
reg  [ 0:0]                      I4003a2515229ca8eb6fefa2bef289ca6;
reg  [MAX_SUM_WDTH_L-1:0]        I086402c82ec67ae09a9e6360c58904b4;
wire  [MAX_SUM_WDTH_L-1:0]       Ibc96fe0a6bf1f95036f97c7d44fab575;
wire  [MAX_SUM_WDTH_L-1:0]       I755a38220a693ba43701d30e7e9508ad;
wire  [MAX_SUM_WDTH_L-1:0]       I896fb82baa9647a14f4b5b1ecfa70a15;
wire  [MAX_SUM_WDTH_L-1:0]       I23d1c973d7a2048353fbb68e4a294c08;
reg  [ 0:0]                      I48672f8b83eef8c406694676746469e7;
reg  [MAX_SUM_WDTH_L-1:0]        I1cefdc831c146187c77f861b3e2d1af0;
wire  [MAX_SUM_WDTH_L-1:0]       If9fd1e08af14f2fd4ca363383f48580a;
wire  [MAX_SUM_WDTH_L-1:0]       I8f3782f78d88a5c3bc93709564999b30;
wire  [MAX_SUM_WDTH_L-1:0]       I986d61d79ce31f4677f3293339db6ad2;
wire  [MAX_SUM_WDTH_L-1:0]       Ica4d93d9fad21316002008ade5106a9d;
reg  [ 0:0]                      Ia14a60c9497c0faf3f1f448ff2abe553;
reg  [MAX_SUM_WDTH_L-1:0]        Ida9c16ae57d17b6faee8a54838860447;
wire  [MAX_SUM_WDTH_L-1:0]       If77592d5d8bed32477fd690341e543d0;
wire  [MAX_SUM_WDTH_L-1:0]       I25b70c6b830cbfe1b41d8f289c751924;
wire  [MAX_SUM_WDTH_L-1:0]       I2a5d65eeffa18dd9af9fe36463dafd7c;
wire  [MAX_SUM_WDTH_L-1:0]       Ibafa6e10bd4edf5d224fdeb2f9adbf98;
reg  [ 0:0]                      I0ef3962dd323e8ec64c4a881bd4b3044;
reg  [MAX_SUM_WDTH_L-1:0]        Ia3b9fb112f39dd0ccbf7555659369efb;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc25402bd879bc5c43b4945b60cd4540;
wire  [MAX_SUM_WDTH_L-1:0]       Iec48da6882325d8a33e0e0e845eb18a0;
wire  [MAX_SUM_WDTH_L-1:0]       I0fd05e46862fdf8e614afaa3fd478602;
wire  [MAX_SUM_WDTH_L-1:0]       I6253a59dca81842d9ab6e58cf204abbf;
reg  [ 0:0]                      Ie9b64c34e31dab63c03b3de4528d53fe;
reg  [MAX_SUM_WDTH_L-1:0]        Ib1bfcdc0c972aafc99116ed8c0511445;
wire  [MAX_SUM_WDTH_L-1:0]       Ib18d64bc58b354358ee6ac16785880e2;
wire  [MAX_SUM_WDTH_L-1:0]       I28689b693a7a5f761a1f252aa3ef3b67;
wire  [MAX_SUM_WDTH_L-1:0]       I1a4e6d12f9776d5e61094e0b5edf71d9;
wire  [MAX_SUM_WDTH_L-1:0]       I8e1ad23b7ac662bb827a83d3709f0adb;
reg  [ 0:0]                      I5941476ded9f6dc25d7394f5d133955b;
reg  [MAX_SUM_WDTH_L-1:0]        I7adff505c50450a04f1717cac1adebe7;
wire  [MAX_SUM_WDTH_L-1:0]       I000ad2287813072cc18dad933758f2ab;
wire  [MAX_SUM_WDTH_L-1:0]       I7bc3698b51b89ac38ba5f4b5428a0c96;
wire  [MAX_SUM_WDTH_L-1:0]       I78aea1705621e2845a331c3e61a8055b;
wire  [MAX_SUM_WDTH_L-1:0]       I0a31314c3580f5f9e61e79c133e5d794;
reg  [ 0:0]                      Ib46c78ff661ee6fb69c704d39235ffe1;
reg  [MAX_SUM_WDTH_L-1:0]        I699feb4382974a02b21cb387c13f7f3f;
wire  [MAX_SUM_WDTH_L-1:0]       I0e274fd7bfc0388fef95a8ceb939ee91;
wire  [MAX_SUM_WDTH_L-1:0]       Id6f39ddcb73d3f4ec081a365d11d1ef4;
wire  [MAX_SUM_WDTH_L-1:0]       I807770bfa86d160459d6ec3c0f4d6a0b;
wire  [MAX_SUM_WDTH_L-1:0]       I31c89b8a11a3090bfd74b112cbc474bb;
reg  [ 0:0]                      Iadabc5abc7dfbc1dd747179ad7e37850;
reg  [MAX_SUM_WDTH_L-1:0]        Idc99c3b23e49aca3c98f0685ea34441c;
wire  [MAX_SUM_WDTH_L-1:0]       I79b82cb1bfc72bd5a9d313b9e9c9203c;
wire  [MAX_SUM_WDTH_L-1:0]       Ib1046ae03c9a77fd2c0b3e9838e9af87;
wire  [MAX_SUM_WDTH_L-1:0]       Ic63723fd43cbbbde51c233a3cca15d3f;
wire  [MAX_SUM_WDTH_L-1:0]       I3abbb59abada1aec6941185f95f738bd;
reg  [ 0:0]                      I97a6b5f0976feceee3a5b5890d4d76a0;
reg  [MAX_SUM_WDTH_L-1:0]        Ib67318fa6954ec8f3247927d34e74f8c;
wire  [MAX_SUM_WDTH_L-1:0]       I8d5bd7039a77ce82ce0f6cbba9c2a076;
wire  [MAX_SUM_WDTH_L-1:0]       I527ad0b9382dd7b6e657dc1a32d8e472;
wire  [MAX_SUM_WDTH_L-1:0]       I8de02f32e14e719f4930d99743c04a20;
wire  [MAX_SUM_WDTH_L-1:0]       I7614dd5e9628c761dd9b2a512cb1da98;
reg  [ 0:0]                      I7217d4790fec9797a1eb8cab1ebce71b;
reg  [MAX_SUM_WDTH_L-1:0]        I8774ce3f11362915c4331d1026e452dd;
wire  [MAX_SUM_WDTH_L-1:0]       Icae7efa4742dd0ad943ee1f67b0c9b14;
wire  [MAX_SUM_WDTH_L-1:0]       Ieb1854b79e9a2bc6cf5aa1c319e8e753;
wire  [MAX_SUM_WDTH_L-1:0]       Iff50b77f300183ca59a67ccbcc9573c4;
wire  [MAX_SUM_WDTH_L-1:0]       I4868604f8178663de759d4c63dc6c4bd;
reg  [ 0:0]                      I3dd024db4130c105a6817e8a4935de0d;
reg  [MAX_SUM_WDTH_L-1:0]        I2392b2d17ffed6073875fbe8e92534cf;
wire  [MAX_SUM_WDTH_L-1:0]       Ife992a151986c58df4cba79b6bc4ac0a;
wire  [MAX_SUM_WDTH_L-1:0]       I9ab973fb74d9fac5d78eb8fc2c7ecf36;
wire  [MAX_SUM_WDTH_L-1:0]       I5ee7916e859b86a98538659401685016;
reg  [ 0:0]                      Iae502e5a5ae518fb7b817afff28b7932;
reg  [MAX_SUM_WDTH_L-1:0]        I3a4f0d3e32596ef05477f494768d4266;
wire  [MAX_SUM_WDTH_L-1:0]       I48c284cefb8cfb5a938a8f23ce4d7f03;
wire  [MAX_SUM_WDTH_L-1:0]       I5c1fc666b77a689478654dd29519f458;
wire  [MAX_SUM_WDTH_L-1:0]       I38bba98b59184c75ba3b27e1dcf52182;
reg  [ 0:0]                      Ib8b2b1d90204af5b100379ecad20fc0f;
reg  [MAX_SUM_WDTH_L-1:0]        Icd08ff59cf6be3ba97698dd55703339e;
wire  [MAX_SUM_WDTH_L-1:0]       I6905b65403c16b0211643227ece536f6;
wire  [MAX_SUM_WDTH_L-1:0]       I3ed34401bba9d5f229bc98480aedd9a5;
wire  [MAX_SUM_WDTH_L-1:0]       Ib4d05804277cddc7f00ac17ac14f5325;
reg  [ 0:0]                      Idf0e651d0b13e167df3c0cc40d149c29;
reg  [MAX_SUM_WDTH_L-1:0]        I985fb7ed22a8476ea322c9e3c2b3851c;
wire  [MAX_SUM_WDTH_L-1:0]       I41babdca6d3fa462849592d37b0a7998;
wire  [MAX_SUM_WDTH_L-1:0]       I58cfec706dc929ebfdeaca6e01b00c0a;
wire  [MAX_SUM_WDTH_L-1:0]       I7efe3c5b2fc69840a79545e0399ce749;
reg  [ 0:0]                      I89daaca029498d05ca62c095db439eb5;
reg  [MAX_SUM_WDTH_L-1:0]        Ib985709316b1b0a9d3fa3c1eaf6c641f;
wire  [MAX_SUM_WDTH_L-1:0]       I70e3eeb2b3966676d16a6aa4c85753ab;
wire  [MAX_SUM_WDTH_L-1:0]       I2a32d545d1e7beecc7531174c7e8dfbc;
wire  [MAX_SUM_WDTH_L-1:0]       Ib8fb40e4ba0ba1f5e9f5a99d1271ed06;
wire  [MAX_SUM_WDTH_L-1:0]       Ica792cb9850a61fa4a8bd8a4b6c6ca05;
reg  [ 0:0]                      I0fe5a34ceda936d0924efdd07fad11e5;
reg  [MAX_SUM_WDTH_L-1:0]        I4be898887dff6e2cebe53f135ece131b;
wire  [MAX_SUM_WDTH_L-1:0]       I779e5997c66649d6d54fd7f0514c47bd;
wire  [MAX_SUM_WDTH_L-1:0]       I5aa578b0c2831453683fa44af1878cb8;
wire  [MAX_SUM_WDTH_L-1:0]       I735d6229ef1a4ecda0a1f1dbdfb53fc1;
wire  [MAX_SUM_WDTH_L-1:0]       I62affd47512c5e8f0979244115624d97;
reg  [ 0:0]                      I7876cbb2b5d8aba3652ec8b218080dff;
reg  [MAX_SUM_WDTH_L-1:0]        I004db04f61fb57aba81e15cc015442b3;
wire  [MAX_SUM_WDTH_L-1:0]       I14fe27afb3df5531b18dc9604e8dbe65;
wire  [MAX_SUM_WDTH_L-1:0]       Ib1b1626c84dad8ad13c058f921ffd57d;
wire  [MAX_SUM_WDTH_L-1:0]       Idf4a4bdddb88c21c5afe10a02373a6eb;
wire  [MAX_SUM_WDTH_L-1:0]       Iadefc2a3d07ed4b2c3c46b2ab5dec252;
reg  [ 0:0]                      If692ff56ce90d22d7af881599c54df75;
reg  [MAX_SUM_WDTH_L-1:0]        I8f7e3dfb2f728d4cd1e79b82b62b0406;
wire  [MAX_SUM_WDTH_L-1:0]       I19315957077b037ffc6415dbb06ef789;
wire  [MAX_SUM_WDTH_L-1:0]       I1f9be09334407fc86c83a7c127e17bbe;
wire  [MAX_SUM_WDTH_L-1:0]       I28e17a5af7a7286a2643100d6d058dc0;
wire  [MAX_SUM_WDTH_L-1:0]       Icb2297c397bfe56be251ffb6b249a020;
reg  [ 0:0]                      I18a7a4fe8931c79df3a69223af46c440;
reg  [MAX_SUM_WDTH_L-1:0]        I991054370345e61638ddaf81785505bd;
wire  [MAX_SUM_WDTH_L-1:0]       I64a48984527d660002f1f82c376c7a84;
wire  [MAX_SUM_WDTH_L-1:0]       I238b5fc70ce9f05b6322a2691b3a0207;
wire  [MAX_SUM_WDTH_L-1:0]       I00c16e7ad3821981032a42d5baa767b3;
wire  [MAX_SUM_WDTH_L-1:0]       I42fd5b094da200b33036e6cb8c7d0286;
reg  [ 0:0]                      I8eec3538b8cc9c046954b6804cc656b0;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa1f503965270d10e7a5c9a15576069b;
wire  [MAX_SUM_WDTH_L-1:0]       I98b7e26a0e9ec9ad750ff87cc0641a73;
wire  [MAX_SUM_WDTH_L-1:0]       I3ec904916870171bf837e162d1030052;
wire  [MAX_SUM_WDTH_L-1:0]       Iedb11b97900b7dd769d31f8a89521975;
wire  [MAX_SUM_WDTH_L-1:0]       Id0dceec6497c9f13ada07138986d4145;
reg  [ 0:0]                      I653767e659590c1676edf6c25fc0e253;
reg  [MAX_SUM_WDTH_L-1:0]        I24f773842a4742fb58d09cae45717b2f;
wire  [MAX_SUM_WDTH_L-1:0]       Ibfe7d9bac29b8838f20cdcfe8ef7da0c;
wire  [MAX_SUM_WDTH_L-1:0]       I4d6c95605595942a34573d6ed55eb326;
wire  [MAX_SUM_WDTH_L-1:0]       Id6d8f32958dfa1a98958a84e7f1aed02;
wire  [MAX_SUM_WDTH_L-1:0]       I971cdf9ddd1bfff5664eec35f22da335;
reg  [ 0:0]                      I5ff863be142b92dff89f7916d0d088c1;
reg  [MAX_SUM_WDTH_L-1:0]        I5bac7e0d778a547a0ae764fe259b6f7a;
wire  [MAX_SUM_WDTH_L-1:0]       Idd8bc1412a0dc5f489ef253a6164ceea;
wire  [MAX_SUM_WDTH_L-1:0]       Idbeec36de0128e5924e214877c82bf11;
wire  [MAX_SUM_WDTH_L-1:0]       I50a9cd240979bc56421bf85011ae99ed;
wire  [MAX_SUM_WDTH_L-1:0]       I6437095f6bad2d4fb2fbe0361f60bba1;
reg  [ 0:0]                      I49f9fd0e0719be527f2a54814dab83ea;
reg  [MAX_SUM_WDTH_L-1:0]        I255577ebee6768871df0224fc1db2db3;
wire  [MAX_SUM_WDTH_L-1:0]       Ie9b6eb3bbac26635aa00c38110958d46;
wire  [MAX_SUM_WDTH_L-1:0]       I9f34e81e3ffb85539a6273babc2a732e;
wire  [MAX_SUM_WDTH_L-1:0]       Id0a1ab8472d704001e0eba0317b117d6;
reg  [ 0:0]                      I945f2476eb599844cbee0cd89038e392;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7fb4af3d3529a32f902a52cf5598474;
wire  [MAX_SUM_WDTH_L-1:0]       I9e632217cd0561d8faa28e4b8850d995;
wire  [MAX_SUM_WDTH_L-1:0]       Iedeb5b7b2fa8acf1ea083102678710ea;
wire  [MAX_SUM_WDTH_L-1:0]       I972431d1f5af0bdf4828e4f85591e358;
reg  [ 0:0]                      Ied0c5f8a9243cd9d93672ad6cc907d21;
reg  [MAX_SUM_WDTH_L-1:0]        I2c98806141f064c9e92935b23a84ede1;
wire  [MAX_SUM_WDTH_L-1:0]       I1f41024b715d8312944ccbf70e95bb40;
wire  [MAX_SUM_WDTH_L-1:0]       Ia6bb5ca05f5d0af452c994dd50004e1d;
wire  [MAX_SUM_WDTH_L-1:0]       I9a1d1d1c862808f9a769cbdb3bc634e1;
reg  [ 0:0]                      I9134c7f579723c7615af60b4344efe76;
reg  [MAX_SUM_WDTH_L-1:0]        I5680847bc8d224fa4ed93b2fc0d841e1;
wire  [MAX_SUM_WDTH_L-1:0]       I9734eb86f4e73ba217739baf5cb1b13c;
wire  [MAX_SUM_WDTH_L-1:0]       Ifc0fe00f86569956df72d8a960337e8c;
wire  [MAX_SUM_WDTH_L-1:0]       I223341a807a1d555f759632f67815159;
reg  [ 0:0]                      Ie92388a9d1e71d73c07ed86e9bf6c887;
reg  [MAX_SUM_WDTH_L-1:0]        I365254279ebb10dd7ba0b3482d5e34cd;
wire  [MAX_SUM_WDTH_L-1:0]       I6c1f5cdf5f2917118941f4af14d67fef;
wire  [MAX_SUM_WDTH_L-1:0]       Ie84e88fd1aa2a0b90aa1715fcd27a329;
wire  [MAX_SUM_WDTH_L-1:0]       I558f70d7039a8bb58d8ea3f72e43dac0;
wire  [MAX_SUM_WDTH_L-1:0]       I9924269ed3de12f1f2a28893c7f95292;
wire  [MAX_SUM_WDTH_L-1:0]       If1153befd1396be2798cc14535ddeb8a;
reg  [ 0:0]                      I6804fecdf59233c6cf14409bf2f1e430;
reg  [MAX_SUM_WDTH_L-1:0]        I57bf4ad773cc058ae1bb7b1911dc3174;
wire  [MAX_SUM_WDTH_L-1:0]       I9bc447b20687fb3e7eff45792bd4dc3a;
wire  [MAX_SUM_WDTH_L-1:0]       If590520f01e452db9867a8d6d5dab29b;
wire  [MAX_SUM_WDTH_L-1:0]       Id93ee7d283016ab9b0aaa21237237c54;
wire  [MAX_SUM_WDTH_L-1:0]       Ic1cf03baabaed466fe532e4db3a9ea78;
wire  [MAX_SUM_WDTH_L-1:0]       If3031f9aa8f6eba90eac12db7839fefd;
reg  [ 0:0]                      I9e777a342bf53eaba0280737ae404bc1;
reg  [MAX_SUM_WDTH_L-1:0]        I57072dfb29c4a3d2e2b40e46e62f0d95;
wire  [MAX_SUM_WDTH_L-1:0]       I0dc2708970ca2b6c092273b6626bacd6;
wire  [MAX_SUM_WDTH_L-1:0]       Ia58944aebf0b4f0a7d76a1444fced9de;
wire  [MAX_SUM_WDTH_L-1:0]       Iedd8e69679d10e05f2889f1d71cf0e7b;
wire  [MAX_SUM_WDTH_L-1:0]       I90f0d471914a2333b9dc14d6d01cf927;
wire  [MAX_SUM_WDTH_L-1:0]       Idceeb22013af64b6bb9f0d773e9ffe9a;
reg  [ 0:0]                      Ied53820aab06b5c3423b1d878c71948f;
reg  [MAX_SUM_WDTH_L-1:0]        Id8cafb6f76321bdaba9711133be7be99;
wire  [MAX_SUM_WDTH_L-1:0]       If43574342e60a625fb6bee5a495e88f3;
wire  [MAX_SUM_WDTH_L-1:0]       Id285f055275014d9f23d35f91879afa1;
wire  [MAX_SUM_WDTH_L-1:0]       I8c803ab08db372802117de4fa4e2a187;
wire  [MAX_SUM_WDTH_L-1:0]       I13ba48a6b360f3cff5f37ce60cb735c6;
wire  [MAX_SUM_WDTH_L-1:0]       I4547cd1dad45dfd01e335e8cf20eadd6;
reg  [ 0:0]                      I24cceded372d782c67b33f3a78b16045;
reg  [MAX_SUM_WDTH_L-1:0]        I6344e71ca2b0fd39d36caedd889c3085;
wire  [MAX_SUM_WDTH_L-1:0]       I0a305655b815b0cc159ac1c5f4ce30f8;
wire  [MAX_SUM_WDTH_L-1:0]       I3633737da6b74284b0ea9a06c3f5875f;
wire  [MAX_SUM_WDTH_L-1:0]       Ia949c1b338d1cba07cf6bb6572c3e322;
reg  [ 0:0]                      I2e78d36bca5bfb016af674c343f9c041;
reg  [MAX_SUM_WDTH_L-1:0]        I0c99a68e0bed90afce18807acf7d55bb;
wire  [MAX_SUM_WDTH_L-1:0]       I9a0185f8400159415bc0ad6c38284041;
wire  [MAX_SUM_WDTH_L-1:0]       I3eeffe43e7deed7ee77a7f5a3bce3cd2;
wire  [MAX_SUM_WDTH_L-1:0]       I85af0c31ca7002ae569d9f5ce39943f7;
reg  [ 0:0]                      I17a9a995de58643dbbfb78604f26198b;
reg  [MAX_SUM_WDTH_L-1:0]        I1c95650979c86310ae2a949961c9db11;
wire  [MAX_SUM_WDTH_L-1:0]       I3dfb8d2fad83fbd807fbfc6330c5b857;
wire  [MAX_SUM_WDTH_L-1:0]       Ic12be21bcba5fa49437cc44dd8a7f064;
wire  [MAX_SUM_WDTH_L-1:0]       I713a384d022d3012e3d0019f5c4ac077;
reg  [ 0:0]                      Iad642c4c62766e8f8bd5a1e9e73bdc80;
reg  [MAX_SUM_WDTH_L-1:0]        I04eaefa5d133e53494fc270b07be7043;
wire  [MAX_SUM_WDTH_L-1:0]       I80550019479d0323d0dd7e7d0f767d83;
wire  [MAX_SUM_WDTH_L-1:0]       Ib8a866f080dd997e0b6c93b6c844d1bc;
wire  [MAX_SUM_WDTH_L-1:0]       Id542de206d736ee3769ea0bd037cb627;
reg  [ 0:0]                      I96f92481be1ac6cf985b8ab387d326bf;
reg  [MAX_SUM_WDTH_L-1:0]        I4a64fa2412eb8058c2dfd9351d7b297d;
wire  [MAX_SUM_WDTH_L-1:0]       I77e6cdb09c92492c3303d0213de9c291;
wire  [MAX_SUM_WDTH_L-1:0]       I788c33a9f94b26f4ce0f515891d06f90;
wire  [MAX_SUM_WDTH_L-1:0]       Iaf7074c2b570a296fe2ea8a5a7097ca0;
wire  [MAX_SUM_WDTH_L-1:0]       I8964c6d3f8e02866a6ad86553ab05d99;
reg  [ 0:0]                      Ie03c09039ccafb427153d2347c1caea8;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8bb2fcb752c6a33254963d1ebb4130d;
wire  [MAX_SUM_WDTH_L-1:0]       I2aa25edaca90c9dae8ed63b48d333c17;
wire  [MAX_SUM_WDTH_L-1:0]       I51a440917c7ae23339bec6f8a745c103;
wire  [MAX_SUM_WDTH_L-1:0]       I56ce875e4619d4d8d6ca2fa0ddee91b1;
wire  [MAX_SUM_WDTH_L-1:0]       I80607da8f92f5a5d2e4798a62a7b1c5c;
reg  [ 0:0]                      Ie7381a8294b4cdf669b9c57cfe4012b5;
reg  [MAX_SUM_WDTH_L-1:0]        Iac05b7e3ae18f948b72c356ccfb8000f;
wire  [MAX_SUM_WDTH_L-1:0]       Ic4dcaa520e26bac40b3876f02074f856;
wire  [MAX_SUM_WDTH_L-1:0]       I3b2714d34081a3b6cccc47fa1638e72e;
wire  [MAX_SUM_WDTH_L-1:0]       I2db1d1ee8f546c00e512875ce2e13cee;
wire  [MAX_SUM_WDTH_L-1:0]       If80a6bb104ff3b2020e909103c104063;
reg  [ 0:0]                      I61c9e3f8e42f869f4c9c1386325100b3;
reg  [MAX_SUM_WDTH_L-1:0]        I27da3f75cca6c49e55db90306aa68e94;
wire  [MAX_SUM_WDTH_L-1:0]       Iadb72cc5444816fbd132256493930bb4;
wire  [MAX_SUM_WDTH_L-1:0]       I3a8ec1ad07bfada3d2c6ffca88b8b678;
wire  [MAX_SUM_WDTH_L-1:0]       I0aa042b86d9f68d22a49b4eb480a9088;
wire  [MAX_SUM_WDTH_L-1:0]       I89a387374771b68d87d7ff2dcc810829;
reg  [ 0:0]                      I24c5b2de59eb1f43fe1efe687231c4b7;
reg  [MAX_SUM_WDTH_L-1:0]        Idc7fed723190098341225fe01ba65ced;
wire  [MAX_SUM_WDTH_L-1:0]       I2935b3d5c3bba4dddfc7ae03fa77b229;
wire  [MAX_SUM_WDTH_L-1:0]       I4e0c0248f4aa97d263d64dfec36e3aa2;
wire  [MAX_SUM_WDTH_L-1:0]       Ia2871d7493b2727d2cb2fbab596b7e6a;
reg  [ 0:0]                      I43d43acde5f831fc32b7bf5f10b9b3a9;
reg  [MAX_SUM_WDTH_L-1:0]        Ife9065805598960919ee4f14c3cc6fd4;
wire  [MAX_SUM_WDTH_L-1:0]       Ie57adae8873946d6c706074b52a49786;
wire  [MAX_SUM_WDTH_L-1:0]       If5ac85646e4b339a19af658f01d0a17f;
wire  [MAX_SUM_WDTH_L-1:0]       I1c092426f34be030b3e020f40517b0e1;
reg  [ 0:0]                      Ib06e93161fc8ca3be232f4261b04feb1;
reg  [MAX_SUM_WDTH_L-1:0]        I717c5c2d6a2be61593492ae5f17a112f;
wire  [MAX_SUM_WDTH_L-1:0]       Ic719b72ad271bc7c077067518e6bbb98;
wire  [MAX_SUM_WDTH_L-1:0]       Ib87362230682c88d68a0ba70e25f3c20;
wire  [MAX_SUM_WDTH_L-1:0]       Ifcf097a102f8dc1f912022fed893d222;
reg  [ 0:0]                      Ia0dd00f83afc805036f2c6a0e38f725e;
reg  [MAX_SUM_WDTH_L-1:0]        I4c31fa8e6eb648439cdae1de1afe0d6f;
wire  [MAX_SUM_WDTH_L-1:0]       I56483ca3fa550dc59bfa347780cfef7b;
wire  [MAX_SUM_WDTH_L-1:0]       I4aa9f61be376458185c3235442c8fda0;
wire  [MAX_SUM_WDTH_L-1:0]       Id91fde1007d47258273299de80721390;
reg  [ 0:0]                      Ib0a0f924fe3757a1e0aade7017ad9277;
reg  [MAX_SUM_WDTH_L-1:0]        Iead549a9af27f1fced7d9c36e7b5c3f5;
wire  [MAX_SUM_WDTH_L-1:0]       Id58498c34aff2e1216c189b9df88822c;
wire  [MAX_SUM_WDTH_L-1:0]       Ib52e0c68caadcf4dd9636a84f5460e53;
wire  [MAX_SUM_WDTH_L-1:0]       Ie19679053b289bb5a0aad570cc81bd14;
wire  [MAX_SUM_WDTH_L-1:0]       I8862c5ef45b723c9abf5d0ab6854a900;
wire  [MAX_SUM_WDTH_L-1:0]       I30db951a07af96a8ddf59360141b9a6a;
reg  [ 0:0]                      I1ca949071d734d230cdb8adda46c9d79;
reg  [MAX_SUM_WDTH_L-1:0]        I10422eb79364e7d0e21e1643d9060331;
wire  [MAX_SUM_WDTH_L-1:0]       I4855a0a0c6426d33014ce6a4c96965ce;
wire  [MAX_SUM_WDTH_L-1:0]       I362e8db1791718290bd33a79b4fc0855;
wire  [MAX_SUM_WDTH_L-1:0]       I773f0508440fb71d73fd82a372cc0a00;
wire  [MAX_SUM_WDTH_L-1:0]       I792891cecae468d7a87e12f2da62a718;
wire  [MAX_SUM_WDTH_L-1:0]       I33303820ad094d7a0ab53bca722fc609;
reg  [ 0:0]                      I40170922c652fa7fa42abc6f580b5e3d;
reg  [MAX_SUM_WDTH_L-1:0]        I914cb87eba8baa40cd515334e59f26b2;
wire  [MAX_SUM_WDTH_L-1:0]       Iff98739de575e25104c0dc30f08912a5;
wire  [MAX_SUM_WDTH_L-1:0]       I1952614b64ea451e9d0646dcce5dd1cd;
wire  [MAX_SUM_WDTH_L-1:0]       I49c1a7d1c20a25496821ad80c7eff790;
wire  [MAX_SUM_WDTH_L-1:0]       Ie2be17a55e79ca76350e033f227800de;
wire  [MAX_SUM_WDTH_L-1:0]       I737a5b06f848cacf0c8da4985c73c66b;
reg  [ 0:0]                      Ib1ad0b531ac9028971d68f533e7ae566;
reg  [MAX_SUM_WDTH_L-1:0]        I32ed679af4ab759901aee43c9d93eb67;
wire  [MAX_SUM_WDTH_L-1:0]       Iab160609bb21501aa55b662d2010357b;
wire  [MAX_SUM_WDTH_L-1:0]       Ief74f1a9d4a43ee5c9def7b83369bb21;
wire  [MAX_SUM_WDTH_L-1:0]       Id144423f50751e661db3860a8487d004;
wire  [MAX_SUM_WDTH_L-1:0]       I623352a4f6705b21d461d6b32e85c12b;
wire  [MAX_SUM_WDTH_L-1:0]       I28d1dc8dc594977b5058b5bb9f6bfc66;
reg  [ 0:0]                      I0ab0170c7ceffbb58377b65d2ad92093;
reg  [MAX_SUM_WDTH_L-1:0]        Id376dfa5141402f4d41a8858180ed87e;
wire  [MAX_SUM_WDTH_L-1:0]       I5371a83bf9d6f334cf8d1c5b082527e9;
wire  [MAX_SUM_WDTH_L-1:0]       If1605d6646fd267e701668a7245b3b44;
wire  [MAX_SUM_WDTH_L-1:0]       Idf5eb1ac2c5bd92fa08ed935ae298255;
reg  [ 0:0]                      I9ac68f228a93bbf4aa4a559b1364e42e;
reg  [MAX_SUM_WDTH_L-1:0]        I98a384bc62ee03f5ad7df20ef2d9af95;
wire  [MAX_SUM_WDTH_L-1:0]       I44ce30330c4d2d6033a0a970dd2bdd68;
wire  [MAX_SUM_WDTH_L-1:0]       Ic101b8f56ea1e25c6b752583a1b01242;
wire  [MAX_SUM_WDTH_L-1:0]       Ib7cf44e681881e55d2d353280a6319d6;
reg  [ 0:0]                      I375c5f7eac92d853e85e0606011f3fb0;
reg  [MAX_SUM_WDTH_L-1:0]        Icfed259ca2bb2732d8e0c26ef67cd4cf;
wire  [MAX_SUM_WDTH_L-1:0]       I35690f724e964248dbb1e80fb1ea49f8;
wire  [MAX_SUM_WDTH_L-1:0]       I5affa2759148a6baf5b9f0cd3122348c;
wire  [MAX_SUM_WDTH_L-1:0]       Iaeea1f06ff0c6e9cfa43ba14420c3adc;
reg  [ 0:0]                      I94f9b1f2e63748c21ec7222c9641366a;
reg  [MAX_SUM_WDTH_L-1:0]        I20861535c450d6e6bf11c45dac120454;
wire  [MAX_SUM_WDTH_L-1:0]       Iac5a23266c3b038b4b54a916dccdf3a8;
wire  [MAX_SUM_WDTH_L-1:0]       Icdfb7f52cc27b1cfcde90a100d29af13;
wire  [MAX_SUM_WDTH_L-1:0]       I71484d7e00efa02a08b54a1405f2902c;
reg  [ 0:0]                      I55500c1d85c4970932be67cc5cd2e023;
reg  [MAX_SUM_WDTH_L-1:0]        I013929385ad819ddfcfcc59c22902ee3;
wire  [MAX_SUM_WDTH_L-1:0]       I68a9b0607e69e8b3dae64689eb288a33;
wire  [MAX_SUM_WDTH_L-1:0]       I2598c48aad48072a7f216b2ab56ee532;
wire  [MAX_SUM_WDTH_L-1:0]       I796e3a193b1b66fa9a04ca60aee11ea1;
wire  [MAX_SUM_WDTH_L-1:0]       Ic96be7e69faf0f43b92618131cf0c98a;
reg  [ 0:0]                      I36b487cd1a57a3a503e587fdefbb19e4;
reg  [MAX_SUM_WDTH_L-1:0]        I34fffcb07fe82f11fe142f7c37f39155;
wire  [MAX_SUM_WDTH_L-1:0]       I648afe4114ce435bf1d13e0ad54425cf;
wire  [MAX_SUM_WDTH_L-1:0]       If05d7e30b4717e0a1bfd20b90d0539bd;
wire  [MAX_SUM_WDTH_L-1:0]       I5fc356af8a62a1d739cb375fb851e90f;
wire  [MAX_SUM_WDTH_L-1:0]       I22f4c5403fbe33d18f97cf21786cdd80;
reg  [ 0:0]                      Icb5350e8c55a2adb370078a7575e28f8;
reg  [MAX_SUM_WDTH_L-1:0]        I61ca60fde05ed88cce714dcd8c13b827;
wire  [MAX_SUM_WDTH_L-1:0]       I9a1b2b9f924099f1e57fa501ba2e33ba;
wire  [MAX_SUM_WDTH_L-1:0]       If6253af4ebc430e4937269a5f4989b29;
wire  [MAX_SUM_WDTH_L-1:0]       I0427d17423548dbb33cf792883b4be8c;
wire  [MAX_SUM_WDTH_L-1:0]       Ie539faf01ae85253e399308fef98afd6;
reg  [ 0:0]                      I8a7a31327c9e4cbd88ce39fea8971caf;
reg  [MAX_SUM_WDTH_L-1:0]        I4907dd45c158dc7e0041c64f1fb388f6;
wire  [MAX_SUM_WDTH_L-1:0]       Iae6e7c42f250cd9223f18f8830fb177d;
wire  [MAX_SUM_WDTH_L-1:0]       Iff47ec1743b59d7f90e9042af7ce44cb;
wire  [MAX_SUM_WDTH_L-1:0]       I1cf4a55ebab332defa32d2922b885285;
wire  [MAX_SUM_WDTH_L-1:0]       I284913858691ad5724073b73a820047a;
reg  [ 0:0]                      Ied069655ed3775819d0bcb722d6d0488;
reg  [MAX_SUM_WDTH_L-1:0]        I2c8f6a9b9f655b317bb0af4d60fdbc4b;
wire  [MAX_SUM_WDTH_L-1:0]       I35626ca53adbbf0a3a71cc6fcf43bcb1;
wire  [MAX_SUM_WDTH_L-1:0]       I0d74ef22d31abcec73c7c582310b1e6d;
wire  [MAX_SUM_WDTH_L-1:0]       I15f4cf1aa0ad5ce2bda52df338e677e3;
wire  [MAX_SUM_WDTH_L-1:0]       I6c5ca5e68c8844bb1617a2288b5bbc37;
reg  [ 0:0]                      I78a5fc80d42e8db1b56cce5f4c97e325;
reg  [MAX_SUM_WDTH_L-1:0]        Ic7dff631559304ec59f0696c66436d62;
wire  [MAX_SUM_WDTH_L-1:0]       I44343a9491069c3c8ea4fbd6255a5a6c;
wire  [MAX_SUM_WDTH_L-1:0]       I1d8318b94d86e1fd28323a5e5684a37b;
wire  [MAX_SUM_WDTH_L-1:0]       I825e83bd88575868f4fcc9a8b8729663;
wire  [MAX_SUM_WDTH_L-1:0]       I3184a16c71cff80c8c90b40e45f114b8;
reg  [ 0:0]                      I3ade7e345432319c1a9c91d4068b3ec9;
reg  [MAX_SUM_WDTH_L-1:0]        I6a239d3e55b4a9a3be9989a85bbec545;
wire  [MAX_SUM_WDTH_L-1:0]       Iae133550f8bad8357a73e7de1372faa3;
wire  [MAX_SUM_WDTH_L-1:0]       Ibccb4a43c410f698e0fff68553326a77;
wire  [MAX_SUM_WDTH_L-1:0]       I72dc7aa294a3af89101ea62a4223170e;
wire  [MAX_SUM_WDTH_L-1:0]       I91eb3e70921e0b141a344bc57dfbc934;
reg  [ 0:0]                      I88aed46f6dad7a81006562a720670654;
reg  [MAX_SUM_WDTH_L-1:0]        I630f905e55f08e7d1569a08e937ad216;
wire  [MAX_SUM_WDTH_L-1:0]       I1986f22f2269cc135c6ed28d35fb0bd1;
wire  [MAX_SUM_WDTH_L-1:0]       Ibef24017bc71de9c002aafa7ce9a784c;
wire  [MAX_SUM_WDTH_L-1:0]       Ieae3ed78fa2c45507066f4e20d96e956;
wire  [MAX_SUM_WDTH_L-1:0]       I730fd25ffc7778fd4bb02d33cb3870d6;
reg  [ 0:0]                      I79e574dc9c7e18b695c9a2619b71b995;
reg  [MAX_SUM_WDTH_L-1:0]        I8d13eb3669785c4279c685763d4f3fad;
wire  [MAX_SUM_WDTH_L-1:0]       I9a32313f2911b797fb0848f7d97e62b9;
wire  [MAX_SUM_WDTH_L-1:0]       I6373e2d64fdb5dd77733b3e4bb405121;
wire  [MAX_SUM_WDTH_L-1:0]       Ib437aa67ab7c13b45d7a4d56ce9e79b8;
wire  [MAX_SUM_WDTH_L-1:0]       I0cb5c7a759f4c75d4a675f9777f15c5f;
reg  [ 0:0]                      I800ef583bec1d46d3d4ffdea6b312ef9;
reg  [MAX_SUM_WDTH_L-1:0]        I25a6f3de9a9a01cbbdd32ed848561aa4;
wire  [MAX_SUM_WDTH_L-1:0]       I0ca91c1426ba14a7b47a081cb3becd19;
wire  [MAX_SUM_WDTH_L-1:0]       I0737e0cc7453e328efab2277bb712ea8;
wire  [MAX_SUM_WDTH_L-1:0]       I456af863661122cc303fccb235f3c7a1;
wire  [MAX_SUM_WDTH_L-1:0]       Idc5916c4800e9f647d51c52444ab6fff;
reg  [ 0:0]                      I56cc5cd6d0a5a4e4601fd48e838fdaf3;
reg  [MAX_SUM_WDTH_L-1:0]        Iba3dd4b2c2c85c4cfe770d9b52ef4634;
wire  [MAX_SUM_WDTH_L-1:0]       I57aca70e2b8d126c120736b2606ed333;
wire  [MAX_SUM_WDTH_L-1:0]       Ic6650a6d092b749b4498c08d69cf815e;
wire  [MAX_SUM_WDTH_L-1:0]       Ic2e3b8f91eb218650c7b9c515c7efe97;
wire  [MAX_SUM_WDTH_L-1:0]       I93a084aa1e6881ab8dc905dcdcdfd7ee;
reg  [ 0:0]                      I21047a3955b8b89bdb9013d571b2bd0d;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1b744387b5200a504e4874e14d2f282;
wire  [MAX_SUM_WDTH_L-1:0]       I8cba172573be52c5a90bd40e6f40a508;
wire  [MAX_SUM_WDTH_L-1:0]       I1cccfd1516af59265731121dde878116;
wire  [MAX_SUM_WDTH_L-1:0]       Ia171bbefe2d20b4c058126c33ef28eb8;
wire  [MAX_SUM_WDTH_L-1:0]       I84bc44a5d53a8f66b985b70c7ec1ae7c;
reg  [ 0:0]                      I56eb529a34b484cd20e29958cd6878eb;
reg  [MAX_SUM_WDTH_L-1:0]        Icf76cb69aedf4db01cd3444f4c4ba471;
wire  [MAX_SUM_WDTH_L-1:0]       I321b104ca3c818018d4b03adfe1110b9;
wire  [MAX_SUM_WDTH_L-1:0]       Ia79b8994da536c86634bf6f54a21145d;
wire  [MAX_SUM_WDTH_L-1:0]       I4df55ce80eec5fee295b5a0ae92bd6c8;
wire  [MAX_SUM_WDTH_L-1:0]       I46593a7956590d870fe680228081a6d2;
reg  [ 0:0]                      I74588df6399af2c1112e3fa557e89e17;
reg  [MAX_SUM_WDTH_L-1:0]        I4857b5b50556c8e7fff4b2d3e08e4b28;
wire  [MAX_SUM_WDTH_L-1:0]       I906e9da31de73ae45579607a014e8b54;
wire  [MAX_SUM_WDTH_L-1:0]       If5dd1a1b9e3fc0e67a85da3183480aed;
wire  [MAX_SUM_WDTH_L-1:0]       Iadfb1571c78c3f0c05e4ef498267df24;
wire  [MAX_SUM_WDTH_L-1:0]       Icebb43b184c2745cc9da9d01b06bc62f;
reg  [ 0:0]                      Ic8eae1a92f46db040eb22d726c3a0e6d;
reg  [MAX_SUM_WDTH_L-1:0]        I0a1e9cf99f1d4725327615f50fcc3ad0;
wire  [MAX_SUM_WDTH_L-1:0]       I6e4b0489ec7333abf2245a1b72a8923d;
wire  [MAX_SUM_WDTH_L-1:0]       I24ac5dd30526c1d3bc7b941103a66804;
wire  [MAX_SUM_WDTH_L-1:0]       I33681b2292c086fe536dae2aec70903a;
wire  [MAX_SUM_WDTH_L-1:0]       Ia373ca76c3b15a4148532b3822f82ba5;
reg  [ 0:0]                      I854a15bc7e9728b01c9a1960f6248dc9;
reg  [MAX_SUM_WDTH_L-1:0]        Ie844f4c446983ce381b0bc4c0e8ef7d7;
wire  [MAX_SUM_WDTH_L-1:0]       I7d08adbaf66cea04be4891db610bca3f;
wire  [MAX_SUM_WDTH_L-1:0]       Ic09ed51b20f411683a801eaad61657a3;
wire  [MAX_SUM_WDTH_L-1:0]       I6a9af8c9009b5de47ebe9ee8b79d3831;
wire  [MAX_SUM_WDTH_L-1:0]       Ife18e8a16d4437161b75a93e3dff1b5b;
reg  [ 0:0]                      Iae332cfd000fd0529684ab787041b5dc;
reg  [MAX_SUM_WDTH_L-1:0]        I6067f47cccceea96ac46ff0d457b25f2;
wire  [MAX_SUM_WDTH_L-1:0]       I0cde86532c8db1a32d9fbe38a40b91b8;
wire  [MAX_SUM_WDTH_L-1:0]       I49c8ec4cd33e6caed8ed7dab779e7ebb;
wire  [MAX_SUM_WDTH_L-1:0]       Idb86f95570587a0711d796aac7004c25;
wire  [MAX_SUM_WDTH_L-1:0]       I2d1373d0b18992fa46a9607a86d21520;
reg  [ 0:0]                      I70148fe95244eebf7f0ec953703398de;
reg  [MAX_SUM_WDTH_L-1:0]        Ifd6fd1f3cbf8884ca7f64bc42278e4fa;
wire  [MAX_SUM_WDTH_L-1:0]       I30f26e090ab14551cbac41883ad8a152;
wire  [MAX_SUM_WDTH_L-1:0]       Ib1b4e41ab25733d1d6dd54e1fe81a419;
wire  [MAX_SUM_WDTH_L-1:0]       I146c0d5154a6de44c0536de873904ccf;
wire  [MAX_SUM_WDTH_L-1:0]       I8eb9d4839a478a4e28b45a549b5682a4;
reg  [ 0:0]                      I24ee2d953e65fefdc73b3d3c4c0ddd05;
reg  [MAX_SUM_WDTH_L-1:0]        Iaec9fd9e79371676bfa8ff14b4feae52;
wire  [MAX_SUM_WDTH_L-1:0]       I2501ef991a59512c43693ba9d7db8571;
wire  [MAX_SUM_WDTH_L-1:0]       I38213f78fd4dc52f9d2c9b7b22136c1c;
wire  [MAX_SUM_WDTH_L-1:0]       I49ce91ac152279af421bbc6c4d9b8087;
wire  [MAX_SUM_WDTH_L-1:0]       I6a2b7bb2cb3ca2ab932c211a68dded55;
reg  [ 0:0]                      Ie3a5f8eec283fd4f682b5d0f909b051c;
reg  [MAX_SUM_WDTH_L-1:0]        I500757c4eda5d3d899aee47b87da585b;
wire  [MAX_SUM_WDTH_L-1:0]       Idaae6ba9da8754615a2c34ef859492db;
wire  [MAX_SUM_WDTH_L-1:0]       Icaca9fc70a3ec6c48c0e41f8168e2bb9;
wire  [MAX_SUM_WDTH_L-1:0]       I4f69b8ff834c7ab3194bc9390ce0f5f6;
wire  [MAX_SUM_WDTH_L-1:0]       I037cb596cd48c5533ed22bc32518d992;
reg  [ 0:0]                      I781d986d7fd6c2fec3a8cf3f29545174;
reg  [MAX_SUM_WDTH_L-1:0]        I47bf091b0fa74ad511a760bad9d2506c;
wire  [MAX_SUM_WDTH_L-1:0]       I94a89577951de90edc4f73b281ad7364;
wire  [MAX_SUM_WDTH_L-1:0]       Ib7493a1a384aebaa7999ff1fb867fc6b;
wire  [MAX_SUM_WDTH_L-1:0]       I2ceb9e423696539135c5bae5cc2d8d98;
reg  [ 0:0]                      Ib4db8131350f8605e00907234aff901d;
reg  [MAX_SUM_WDTH_L-1:0]        Ia4c3d0cd9957f678880de5775de76e0d;
wire  [MAX_SUM_WDTH_L-1:0]       Ia6bbf236436b2ed22bbaae3b8849de6d;
wire  [MAX_SUM_WDTH_L-1:0]       I33cdaee4676d546dd5507df4704ea1f8;
wire  [MAX_SUM_WDTH_L-1:0]       Ia44daa9ddc3e4d377267333813d4675f;
reg  [ 0:0]                      Ie093f0750b60d3aed75705637933f34c;
reg  [MAX_SUM_WDTH_L-1:0]        If5f957fa2f055b1c2c28e8d7cfe3e9ad;
wire  [MAX_SUM_WDTH_L-1:0]       Ie1f8fff3f43426d6bc39e45322a532ca;
wire  [MAX_SUM_WDTH_L-1:0]       I4ee181895efc22862b6e85802a944095;
wire  [MAX_SUM_WDTH_L-1:0]       I5c24ea83cabbb6be089ac084732cb9d6;
reg  [ 0:0]                      Id2fba7c1b3dc7a75a5e0d90494d56962;
reg  [MAX_SUM_WDTH_L-1:0]        I3608378a5da8c66bef58528d56192530;
wire  [MAX_SUM_WDTH_L-1:0]       Ifee2342449a3b3d0036ce2ecbc9ae189;
wire  [MAX_SUM_WDTH_L-1:0]       I70a9a9b8f25066612a50e411ad68e6c4;
wire  [MAX_SUM_WDTH_L-1:0]       I1870059af857c79d444bef948bb536ef;
reg  [ 0:0]                      I9ecee74c445711a376133636ef414666;
reg  [MAX_SUM_WDTH_L-1:0]        Ie6dead855e00ea0a8e6a9b7503aaebb8;
wire  [MAX_SUM_WDTH_L-1:0]       Iafe61ab12e232a1090123a0f16eefaca;
wire  [MAX_SUM_WDTH_L-1:0]       I10ca809fe9a04eaf5d7784ba69314178;
wire  [MAX_SUM_WDTH_L-1:0]       I7a1bd0a115b3a1f85cb9c54840f5bf9b;
wire  [MAX_SUM_WDTH_L-1:0]       I986a564393d944d7d202414431c6d165;
reg  [ 0:0]                      Ifb3cf6b88835d27220df837682c4dc93;
reg  [MAX_SUM_WDTH_L-1:0]        I3bae5e6862e003a8b9a476f72cc6858b;
wire  [MAX_SUM_WDTH_L-1:0]       I464042aaa60a41c7e1faf3d16eeb121d;
wire  [MAX_SUM_WDTH_L-1:0]       I34b9a0bf2b6b562fb36291022ddf5179;
wire  [MAX_SUM_WDTH_L-1:0]       I17dd8612b5c7f9dcc90f17e584aab2d3;
wire  [MAX_SUM_WDTH_L-1:0]       Id77cf7c05844d83e808a694971145261;
reg  [ 0:0]                      I386fbb3bd550891d682e137044e8773a;
reg  [MAX_SUM_WDTH_L-1:0]        I4431adecba8be9e5f21bc6b3e1f8cb10;
wire  [MAX_SUM_WDTH_L-1:0]       I276c1155d766437253f12b25066b84e4;
wire  [MAX_SUM_WDTH_L-1:0]       Id75b386d8076893cb73baca69c3eff59;
wire  [MAX_SUM_WDTH_L-1:0]       If62ddbe87274965cfd83189c6666401e;
wire  [MAX_SUM_WDTH_L-1:0]       I4f73a07452638a610b31e3ee52cb5639;
reg  [ 0:0]                      I7ede7d2e1c2730b3b71340b11e880f5b;
reg  [MAX_SUM_WDTH_L-1:0]        I21c7a2885126d532d00484376588a469;
wire  [MAX_SUM_WDTH_L-1:0]       I2a4faf3344d9bf4ee71da0be8994788a;
wire  [MAX_SUM_WDTH_L-1:0]       I7d7ad0cbb962a47e229fe9d8406e6fe1;
wire  [MAX_SUM_WDTH_L-1:0]       I82988dc2dc83ac61380d2a5cb6551768;
wire  [MAX_SUM_WDTH_L-1:0]       I058c3a9848fd30010e4742d8682081ac;
reg  [ 0:0]                      I64c65fad4a7d958d625c783626808175;
reg  [MAX_SUM_WDTH_L-1:0]        I2c4d7339ff2fe68d060dd8d961dcab8c;
wire  [MAX_SUM_WDTH_L-1:0]       I368121c2534820a7147858c06e58b3fc;
wire  [MAX_SUM_WDTH_L-1:0]       I03d4541eeb1440aa72ee490c49977e32;
wire  [MAX_SUM_WDTH_L-1:0]       I75fdf5a355949a87b768b1e67db674e4;
wire  [MAX_SUM_WDTH_L-1:0]       I088f4a0af0239602d422324549cb9799;
reg  [ 0:0]                      Ib2e0cd0a2b51c3a265bdd20834c0ed2d;
reg  [MAX_SUM_WDTH_L-1:0]        Iee518b15b067eec58cccfa37f7432ea5;
wire  [MAX_SUM_WDTH_L-1:0]       I787fe66b38237caf805ec14970d154c7;
wire  [MAX_SUM_WDTH_L-1:0]       Icef176cff3ae503dbbe2af9ecfc4c859;
wire  [MAX_SUM_WDTH_L-1:0]       Ie0a66e4871bfe94f6716279ecc9ef21c;
wire  [MAX_SUM_WDTH_L-1:0]       I474adf7a975b405c288058139a08be38;
reg  [ 0:0]                      I67be0b66c8d0680eb23290a4b3885af3;
reg  [MAX_SUM_WDTH_L-1:0]        I42145be9c2a80288ba4a2edd91f661a3;
wire  [MAX_SUM_WDTH_L-1:0]       Iebeadb39658f41dcf8719ed413e46144;
wire  [MAX_SUM_WDTH_L-1:0]       Ie018b0d9f05a86207ae09ca2efac54e2;
wire  [MAX_SUM_WDTH_L-1:0]       I51ee69807609fca0f332c8bc31afd632;
wire  [MAX_SUM_WDTH_L-1:0]       Iee1cb471704b2a8718a68ef93fd2e356;
reg  [ 0:0]                      I01148401f7d058614dc1ae6ed3c8bd94;
reg  [MAX_SUM_WDTH_L-1:0]        I9dc297ad41fafcda77f5347f331cfc25;
wire  [MAX_SUM_WDTH_L-1:0]       I1731c0e3be86eec142c3732ee836e4d5;
wire  [MAX_SUM_WDTH_L-1:0]       Id3b8c0ca32331f94fd98c8dae72bb15d;
wire  [MAX_SUM_WDTH_L-1:0]       I6a86b0a82441c6c14436a3e0af6b0fb7;
wire  [MAX_SUM_WDTH_L-1:0]       I8c92ff598084da7a50f7c68da96620b3;
reg  [ 0:0]                      I3394319c370daf6102be00d938d55769;
reg  [MAX_SUM_WDTH_L-1:0]        I846700c79f30ca954cc2933fc94d355b;
wire  [MAX_SUM_WDTH_L-1:0]       I8bd1862e7bc2e83e9863389d532e6623;
wire  [MAX_SUM_WDTH_L-1:0]       I8053269f8bd78a931878c8350693e1d6;
wire  [MAX_SUM_WDTH_L-1:0]       I2ff66cdd7314276232715ef2361ad184;
wire  [MAX_SUM_WDTH_L-1:0]       Icf541c76bfaf37fe6111de037d205f15;
reg  [ 0:0]                      I24d6a334dd15ccdea558f32cd029e6d1;
reg  [MAX_SUM_WDTH_L-1:0]        I8af96a91457316e49e3f7dd5e57c82da;
wire  [MAX_SUM_WDTH_L-1:0]       I68319c8b9febef9f564832429c91b85a;
wire  [MAX_SUM_WDTH_L-1:0]       I127772614218dd7c50d3136b4f174d7a;
wire  [MAX_SUM_WDTH_L-1:0]       Ib8d1aea4ad24c6ceb44f2cc672e1ff90;
wire  [MAX_SUM_WDTH_L-1:0]       I9ca26c8104bf15f48b19dc3256914544;
reg  [ 0:0]                      I3a41f68bca2d7edd1f5738c4fda8e73c;
reg  [MAX_SUM_WDTH_L-1:0]        I7d1c247500d7d32e406b2a5f7e2b745b;
wire  [MAX_SUM_WDTH_L-1:0]       Icc76d9ffc3f3d7b410205eeb8232a33b;
wire  [MAX_SUM_WDTH_L-1:0]       I7fc4551d8a0445f79b87b4ba5f2ffeaa;
wire  [MAX_SUM_WDTH_L-1:0]       I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8;
wire  [MAX_SUM_WDTH_L-1:0]       Ie34c07af9f6adb9e4b636dce3d0682c0;
reg  [ 0:0]                      I9ef1784d165492f3482d14f475732451;
reg  [MAX_SUM_WDTH_L-1:0]        I66d85c030a8864505298919046056305;
wire  [MAX_SUM_WDTH_L-1:0]       Ib869a349250a765d2f8660e0dbdcf312;
wire  [MAX_SUM_WDTH_L-1:0]       I1a4fb631fdc7b5454c266589962ff5f0;
wire  [MAX_SUM_WDTH_L-1:0]       I9de4e0e86e9edcf948d9eddf0401b94a;
wire  [MAX_SUM_WDTH_L-1:0]       Iee7b4838986c962969c00a0bbe53ce0b;
reg  [ 0:0]                      I9d9378337a77515a4e8d04fb88938808;
reg  [MAX_SUM_WDTH_L-1:0]        I4841257ae596d9d3e4eb1e6f886956b0;
wire  [MAX_SUM_WDTH_L-1:0]       Id81b11a8ca1dd8989e36cef637ae6aab;
wire  [MAX_SUM_WDTH_L-1:0]       Ibe96deab015b799fe7f69bae8432952c;
wire  [MAX_SUM_WDTH_L-1:0]       I986b52155cc1470299321a4933241ed7;
wire  [MAX_SUM_WDTH_L-1:0]       I04be63a04f3942ce749cc9bd7540e055;
reg  [ 0:0]                      If0e20ef9aa69b77ae0e58ca3dfc9998f;
reg  [MAX_SUM_WDTH_L-1:0]        Icd6f7ec117f9ab4eda8c5eba41386ffa;
wire  [MAX_SUM_WDTH_L-1:0]       Ia7adea5b0ec86e9fcd427a5468d72b64;
wire  [MAX_SUM_WDTH_L-1:0]       Ie8990d8abd23f8f9f79d7fe38c57fa8c;
wire  [MAX_SUM_WDTH_L-1:0]       I9d2f90ddddbdbb525d5f070f32546b64;
wire  [MAX_SUM_WDTH_L-1:0]       I905256d73bdb63bf860e15687350795f;
reg  [ 0:0]                      Iec2cb48bb1b58f268bf164d5e8a8120f;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc0498839d1d9b6dc853b8e5d7a88fa3;
wire  [MAX_SUM_WDTH_L-1:0]       I9adcfc18e4471209edbe9a379e996067;
wire  [MAX_SUM_WDTH_L-1:0]       I3d7d048348bf833f744a9f73889b7802;
wire  [MAX_SUM_WDTH_L-1:0]       Id619e8d4040014d0e415ff71c5e0591f;
wire  [MAX_SUM_WDTH_L-1:0]       Iaf3de2ef283e03dd72002026e1299224;
reg  [ 0:0]                      Ia4ae7c98720d43a604f28dfc5dd67d50;
reg  [MAX_SUM_WDTH_L-1:0]        I142ebca7f155e287e38ddf45423ab0fd;
wire  [MAX_SUM_WDTH_L-1:0]       I64551529c0028ec145407be7f5dfef71;
wire  [MAX_SUM_WDTH_L-1:0]       I5ebe580a943b65fb16ea722ba101fd05;
wire  [MAX_SUM_WDTH_L-1:0]       I0921901599c43b27e701758026dd3ee1;
wire  [MAX_SUM_WDTH_L-1:0]       I6033532f27c26b2d42bb3ea128f80dfa;

reg  [MAX_SUM_WDTH_L-1:0]        I5deafec6e5f32da1bcf8f7018cf794d8;
reg  [MAX_SUM_WDTH_L-1:0]        I35b3fb2670f3a60d165c1fd10f02c00c;
reg  [MAX_SUM_WDTH_L-1:0]        I68925439e233444a4da44871f31de94a;
reg  [MAX_SUM_WDTH_L-1:0]        I3108702b5ca506422c1ba6174619f193;
reg  [MAX_SUM_WDTH_L-1:0]        Icc8e8f6446ac64350a05f5e1e0541bb9;
reg  [MAX_SUM_WDTH_L-1:0]        Iadebaf3f6cca1ba78feab50ce70c8aef;
reg  [MAX_SUM_WDTH_L-1:0]        I8681cf376dbeceab29279a7637249e7d;
reg  [MAX_SUM_WDTH_L-1:0]        Ie850a07565bed90389bb125ddcd39658;
reg  [MAX_SUM_WDTH_L-1:0]        I97b77743c2311ec629ea24c933b60053;
reg  [MAX_SUM_WDTH_L-1:0]        I07a0a8d41ed8176e92380f2c89c2afdd;
reg  [MAX_SUM_WDTH_L-1:0]        I021842328f948a94159b32903c8bcb68;
reg  [MAX_SUM_WDTH_L-1:0]        Icaf3bd685005a05c8fb334266ea4e4b9;
reg  [MAX_SUM_WDTH_L-1:0]        I92d9e1d7dcf45a4d738c546e959687c3;
reg  [MAX_SUM_WDTH_L-1:0]        I39ca3a8ca714a9726114326ae6bfab0a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9ae20ed5b2a0cad2c37c5bb2ea05ff4;
reg  [MAX_SUM_WDTH_L-1:0]        I8f131eb6138c23fdcb35195703131e64;
reg  [MAX_SUM_WDTH_L-1:0]        Iff77e08da4bcbb85b95fa277b69653a9;
reg  [MAX_SUM_WDTH_L-1:0]        I703e0a4879a39b3b8b0a49de86ca4ff4;
reg  [MAX_SUM_WDTH_L-1:0]        I3da217f6f2d0f515bb9036673d753a88;
reg  [MAX_SUM_WDTH_L-1:0]        Ifcc06d5a010e01a781ae8a9e9e2b31a0;
reg  [MAX_SUM_WDTH_L-1:0]        I42fd611fec087113ba6e35f281bced9c;
reg  [MAX_SUM_WDTH_L-1:0]        I5bb626e7347bb9ae4219cc72244b38f8;
reg  [MAX_SUM_WDTH_L-1:0]        I47e2dac0068652338f94ddffd2dbe88a;
reg  [MAX_SUM_WDTH_L-1:0]        I59a3f06de2984078a4d4c430a2980fe3;
reg  [MAX_SUM_WDTH_L-1:0]        I857b7fd58279b1063a06a4f33b880ba6;
reg  [MAX_SUM_WDTH_L-1:0]        I3901bbda029cd0a41640001c1efd400f;
reg  [MAX_SUM_WDTH_L-1:0]        Ifceeccf10f1d85a32f70c04654a1a1b4;
reg  [MAX_SUM_WDTH_L-1:0]        I2d810c1d1304658edff74921e8d0f388;
reg  [MAX_SUM_WDTH_L-1:0]        I575b0201be445388607ab83465eab8d6;
reg  [MAX_SUM_WDTH_L-1:0]        I7928c5ce0f821df1cb6271d15e19fa22;
reg  [MAX_SUM_WDTH_L-1:0]        I12695a21c942d02a432cf6382d7d7452;
reg  [MAX_SUM_WDTH_L-1:0]        I00d03f0f71b008dad8035bbf251f41bf;
reg  [MAX_SUM_WDTH_L-1:0]        I41afedcbc0f492e3243436cbefdaf609;
reg  [MAX_SUM_WDTH_L-1:0]        I638c4c2708e437a050ed7cbbac516a59;
reg  [MAX_SUM_WDTH_L-1:0]        I6877d3306b1f08c236b5d1b59f0de259;
reg  [MAX_SUM_WDTH_L-1:0]        Ib3e66aa460f39d32110ea6f115785b3d;
reg  [MAX_SUM_WDTH_L-1:0]        I5e603e8392a5322951b3225b65b19446;
reg  [MAX_SUM_WDTH_L-1:0]        If5da7fa1a615e1122445460e33487772;
reg  [MAX_SUM_WDTH_L-1:0]        Ic4153dafafaf7d047478c5d81109437f;
reg  [MAX_SUM_WDTH_L-1:0]        I7b5476007f04e81afc0125e6a8930303;
reg  [MAX_SUM_WDTH_L-1:0]        I3521a18022925249caddb8e37d2c1262;
reg  [MAX_SUM_WDTH_L-1:0]        Ifd0f52d4f814e2bb4c3bd34c1e09bda7;
reg  [MAX_SUM_WDTH_L-1:0]        I8945f6d420c8b373225451defcd2c805;
reg  [MAX_SUM_WDTH_L-1:0]        Ieec6cb6518cc0d9300de0c4f2d32487d;
reg  [MAX_SUM_WDTH_L-1:0]        Ic62eb7e90d703ef994e68587345a4293;
reg  [MAX_SUM_WDTH_L-1:0]        Id3efd8419da986aa89b8ad8e75848cfa;
reg  [MAX_SUM_WDTH_L-1:0]        I40803f10b7c4dc9ae4969739349b0265;
reg  [MAX_SUM_WDTH_L-1:0]        I7d961743fdeaf1e72e4b25c12a1d4c46;
reg  [MAX_SUM_WDTH_L-1:0]        Ifea156f33eb61fece272efe379327f6e;
reg  [MAX_SUM_WDTH_L-1:0]        Ifc99169b3399f3d14121c1a9bce3fc21;
reg  [MAX_SUM_WDTH_L-1:0]        I6536144383cbda6f3b3c564391866906;
reg  [MAX_SUM_WDTH_L-1:0]        Ic21bf9a8a4cd85ec123d7fe142ed49c0;
reg  [MAX_SUM_WDTH_L-1:0]        I1f31fe6a0ca8510bcadbc2069403150b;
reg  [MAX_SUM_WDTH_L-1:0]        I0e40933d00f4a7d9b53b2764aa0da700;
reg  [MAX_SUM_WDTH_L-1:0]        Ic41a6e00bc84bfc1b8194d15bb899c93;
reg  [MAX_SUM_WDTH_L-1:0]        I2832571f2b0a7fbb41d2e8ca7f64e003;
reg  [MAX_SUM_WDTH_L-1:0]        I9593c853e41952e408a809cb24efa4fd;
reg  [MAX_SUM_WDTH_L-1:0]        I6edffbf4136e193dca0fcec3a74e8e9c;
reg  [MAX_SUM_WDTH_L-1:0]        Ibaed50cc2e36ae58945887d11a6ec9e4;
reg  [MAX_SUM_WDTH_L-1:0]        Ie4570cac44f59e6ff46f73a703026479;
reg  [MAX_SUM_WDTH_L-1:0]        Ibaa136d37936687e9dbe4222749d19c3;
reg  [MAX_SUM_WDTH_L-1:0]        If85de3225f45478827b43b89089cd29e;
reg  [MAX_SUM_WDTH_L-1:0]        I0344b86a6e9c036e103a9c1f3651175f;
reg  [MAX_SUM_WDTH_L-1:0]        I5463d13575e0b9fb8a0f6cc8b35d0ce9;
reg  [MAX_SUM_WDTH_L-1:0]        I8a3c63ef122001a29e5abe93c4e1a48f;
reg  [MAX_SUM_WDTH_L-1:0]        I6a79108484fcb192f6d93bfb98e271c4;
reg  [MAX_SUM_WDTH_L-1:0]        I9001e95b71457a2bd09a9846af370b16;
reg  [MAX_SUM_WDTH_L-1:0]        I51620de618db6327358a5cac97e1e97f;
reg  [MAX_SUM_WDTH_L-1:0]        Ib9c58818059af5c5a03e77a5dcef4654;
reg  [MAX_SUM_WDTH_L-1:0]        I8081c71aa01a8d575bfea6ea7f2f595f;
reg  [MAX_SUM_WDTH_L-1:0]        Iad999607ad8d7da0f3b341f83ea030a6;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7291c914d2cb66f547b0a7717f71311;
reg  [MAX_SUM_WDTH_L-1:0]        Ic01018a5f1bc392bbd267016f6612a83;
reg  [MAX_SUM_WDTH_L-1:0]        Ib11dff839e7e532657b32f29fd9b1651;
reg  [MAX_SUM_WDTH_L-1:0]        I251d7ea16dd5407d22a6846ddcfe12d8;
reg  [MAX_SUM_WDTH_L-1:0]        I773797f81f73b9b6e844441142a1bb48;
reg  [MAX_SUM_WDTH_L-1:0]        I853ecadf30fc10a13dd1ffb1f2dfb5d6;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb8b3c91e1d3b890cfe58f32f8ec3ae3;
reg  [MAX_SUM_WDTH_L-1:0]        I3485d69de942d64e56925da522175b51;
reg  [MAX_SUM_WDTH_L-1:0]        Iae42f12bc0475c8b58341d80027a57cb;
reg  [MAX_SUM_WDTH_L-1:0]        I22fe2af25463f87ee7315a9aac32854e;
reg  [MAX_SUM_WDTH_L-1:0]        Idf44ad78c338c39699721ce511691dfd;
reg  [MAX_SUM_WDTH_L-1:0]        I984a657f9265d41318c0290e249e9712;
reg  [MAX_SUM_WDTH_L-1:0]        I915fccfb1d1ada9aa7c8e24c2eebd04c;
reg  [MAX_SUM_WDTH_L-1:0]        I2bdf58ecd0974720631be830efb48dc8;
reg  [MAX_SUM_WDTH_L-1:0]        Ibaedf6246fa43acc8accb5a24d49cc2f;
reg  [MAX_SUM_WDTH_L-1:0]        I904d13524dcdf55478a5266d50e53ff7;
reg  [MAX_SUM_WDTH_L-1:0]        I22d8e5d57c1bc082169437a654d22bba;
reg  [MAX_SUM_WDTH_L-1:0]        I719cdaa2a2e61a0df7f1fd5efe517426;
reg  [MAX_SUM_WDTH_L-1:0]        I8e92a61eb73c41680652936cfcc614ff;
reg  [MAX_SUM_WDTH_L-1:0]        I7ad5af8319f6da469858300f0777b580;
reg  [MAX_SUM_WDTH_L-1:0]        I32be72eaf04e79120a57ea94296a4e56;
reg  [MAX_SUM_WDTH_L-1:0]        Ie756f6a87d85adb40479ce7cf3545556;
reg  [MAX_SUM_WDTH_L-1:0]        I8794c6ce0a3f2e6697372e2c911ba420;
reg  [MAX_SUM_WDTH_L-1:0]        Ic82b1a29b5e63bcc3686a0d4bf1f5c24;
reg  [MAX_SUM_WDTH_L-1:0]        I253ef976058080beab79646af18e2d5b;
reg  [MAX_SUM_WDTH_L-1:0]        I930dd54c36540d75dc870eef89960163;
reg  [MAX_SUM_WDTH_L-1:0]        Iaf7554cd4e8b5ea6155ec61a8d589b86;
reg  [MAX_SUM_WDTH_L-1:0]        I50907c7d1efa0038d81efed82b192891;
reg  [MAX_SUM_WDTH_L-1:0]        If3e9486d2960d164d94641d4f1917416;
reg  [MAX_SUM_WDTH_L-1:0]        I2bec61db45dd79b98d6ebff6c5a4899e;
reg  [MAX_SUM_WDTH_L-1:0]        I7f31647f3ea6ce7bbd211c25cf4828fb;
reg  [MAX_SUM_WDTH_L-1:0]        Ice65387e606faf9c7b884475b489abba;
reg  [MAX_SUM_WDTH_L-1:0]        I63f914927dcf49552e9f3fe0180a30e8;
reg  [MAX_SUM_WDTH_L-1:0]        I742ff5725e3a18acd03454cf9f313f4b;
reg  [MAX_SUM_WDTH_L-1:0]        I84e4b3bc63ec0b0bff7f98f433c1fd67;
reg  [MAX_SUM_WDTH_L-1:0]        I78c6a1428a1f211c5e89b8c76b3dc033;
reg  [MAX_SUM_WDTH_L-1:0]        I9897cbf9d7cab759f99f5f8f4bc125d0;
reg  [MAX_SUM_WDTH_L-1:0]        I9a6c1ff6dde5141849e4aa925140ebb8;
reg  [MAX_SUM_WDTH_L-1:0]        Icc1c25b229393361f1245c40f573b423;
reg  [MAX_SUM_WDTH_L-1:0]        I53b5a72e41ee53037ee3ae040799f401;
reg  [MAX_SUM_WDTH_L-1:0]        I3cc25fb583118f45babf457fe78d5434;
reg  [MAX_SUM_WDTH_L-1:0]        I20c046dd8a1265e12e902275b73417da;
reg  [MAX_SUM_WDTH_L-1:0]        I1b184c9a34aeb6eda813d86556e235d9;
reg  [MAX_SUM_WDTH_L-1:0]        I70e03db993e1d26d5814ff5fcd38ada1;
reg  [MAX_SUM_WDTH_L-1:0]        I119dc168a44950d215af877eb81152fe;
reg  [MAX_SUM_WDTH_L-1:0]        Id717ed42457eb1d3f4e3edbf0dd72c41;
reg  [MAX_SUM_WDTH_L-1:0]        I79d1f852a03bcc11d6121a12d8c5b86d;
reg  [MAX_SUM_WDTH_L-1:0]        I769e650e49f152c0803b06232740691c;
reg  [MAX_SUM_WDTH_L-1:0]        I1ef3c09b8481f14c3526224430a5f4b9;
reg  [MAX_SUM_WDTH_L-1:0]        I2a38d43a7e25050aa672cbf84a409aa8;
reg  [MAX_SUM_WDTH_L-1:0]        I1c2be5e13c462a8a6b07bca311582ce4;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8fd61caf16aa0e504cc7dc8cec6f0b8;
reg  [MAX_SUM_WDTH_L-1:0]        Icd0fe98ca873ad6dacdf80dfdfc450ec;
reg  [MAX_SUM_WDTH_L-1:0]        I94e1ab698dc93ff0764dc5c1e62179fe;
reg  [MAX_SUM_WDTH_L-1:0]        Ifd48363af9abb390a72991fbdd6f7877;
reg  [MAX_SUM_WDTH_L-1:0]        I44f79397a010088e4ecdcb9669f2efbd;
reg  [MAX_SUM_WDTH_L-1:0]        I124b0b7d91cfb42b0d9722f3229c2d53;
reg  [MAX_SUM_WDTH_L-1:0]        Iadf1875c584adc34f7586a146184a763;
reg  [MAX_SUM_WDTH_L-1:0]        I02d3f9982f02ea85f996bf5b5975b930;
reg  [MAX_SUM_WDTH_L-1:0]        Ia6e1b39d83ddce053518c5ae9a5ca33e;
reg  [MAX_SUM_WDTH_L-1:0]        I3308663053f4307d43ac66f43266f706;
reg  [MAX_SUM_WDTH_L-1:0]        I87ad25dff6c0c9ac46b7a129cb575537;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf5d40b7c46b50866f58f6fa23e1861b;
reg  [MAX_SUM_WDTH_L-1:0]        I0e3a9a3b38875156d15f697adaf95410;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3f87d094e71e4a82f60e8d91cdd768b;
reg  [MAX_SUM_WDTH_L-1:0]        I793f52d174cd09fe000e8d0351753592;
reg  [MAX_SUM_WDTH_L-1:0]        I89ea3da7db40e7e6705020462b2d1df1;
reg  [MAX_SUM_WDTH_L-1:0]        Ib2af2f1a928dd824f25b99f0b602753f;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3e887f5f1a64c37a10404d636212b45;
reg  [MAX_SUM_WDTH_L-1:0]        I5c6a004278f155d33d0cc1b576c3b25f;
reg  [MAX_SUM_WDTH_L-1:0]        I6a03a4a548a0906d1a3e9ce47f3454c6;
reg  [MAX_SUM_WDTH_L-1:0]        I542e525074d049197ac3904e6102f0bd;
reg  [MAX_SUM_WDTH_L-1:0]        Ie0307a43ce71ba73d4c8e5ad556bd341;
reg  [MAX_SUM_WDTH_L-1:0]        Ib03e1d3a1f27721e4ea32629c2e86f85;
reg  [MAX_SUM_WDTH_L-1:0]        I782f4ab4666c9f550a2cfc943cedbe77;
reg  [MAX_SUM_WDTH_L-1:0]        Ib991e16161d5c8b3b655e3c7c08b93c4;
reg  [MAX_SUM_WDTH_L-1:0]        I72f8c6bad4bff3b00055aa8824479931;
reg  [MAX_SUM_WDTH_L-1:0]        I58e5100cc1e9b809e93125fe5d08a9d8;
reg  [MAX_SUM_WDTH_L-1:0]        I0aa7056fdacd6022f328a3be49048856;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2f40b5c49a2284fb6a234bf7472130f;
reg  [MAX_SUM_WDTH_L-1:0]        I8da184aee7953890f2c89e40744402f4;
reg  [MAX_SUM_WDTH_L-1:0]        I613ccfc7dad5627cde02fa1720244d01;
reg  [MAX_SUM_WDTH_L-1:0]        I080fc6c99e506e569b97433f3fdc3e60;
reg  [MAX_SUM_WDTH_L-1:0]        I79aa118ef8ac0d9b13723fb1f5a7e4ad;
reg  [MAX_SUM_WDTH_L-1:0]        I7e6e7601245ca5b3a58b91848e25a6d3;
reg  [MAX_SUM_WDTH_L-1:0]        I2792edda66743635b837aa3bec0c58b9;
reg  [MAX_SUM_WDTH_L-1:0]        I085cc29465c945957d00cbcf804e3ae4;
reg  [MAX_SUM_WDTH_L-1:0]        I74a8e879666bb216a331fd2ab723e37c;
reg  [MAX_SUM_WDTH_L-1:0]        I7a90a43ed71e82862457d9fa40bd005c;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1e7b4bd6201baa02b8d59cb0f6ffb8e;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7b7cdc22b22f276b1c021abaa8fb443;
reg  [MAX_SUM_WDTH_L-1:0]        Ib58e33f31be36b28997ba05ef1004573;
reg  [MAX_SUM_WDTH_L-1:0]        Ibec394e82f499e8d2d5a9524f943d6ac;
reg  [MAX_SUM_WDTH_L-1:0]        Ie06ad127e475dc131859992bb5f350a0;
reg  [MAX_SUM_WDTH_L-1:0]        Ic494a58468b6a7dda76923a9475bf173;
reg  [MAX_SUM_WDTH_L-1:0]        Ib82a2db86d03fe8538fa19d06e501dae;
reg  [MAX_SUM_WDTH_L-1:0]        I5b64727fee9d0825a4ea83261992e489;
reg  [MAX_SUM_WDTH_L-1:0]        Ice7e502b9c2b797719448fde8376087a;
reg  [MAX_SUM_WDTH_L-1:0]        I792b4f73ed7139b8761443cbc0833e39;
reg  [MAX_SUM_WDTH_L-1:0]        I278d57d1964cbf3339db450926ef4782;
reg  [MAX_SUM_WDTH_L-1:0]        I9c1a08b61782ef6c72545504693ac54e;
reg  [MAX_SUM_WDTH_L-1:0]        I363594fb91d01abca7a2b7402e352fd0;
reg  [MAX_SUM_WDTH_L-1:0]        Idd284c75a230f4b97d5acb98a8e38b2d;
reg  [MAX_SUM_WDTH_L-1:0]        If040df53a6410b263f5b3dc3090631c4;
reg  [MAX_SUM_WDTH_L-1:0]        I31df60ffcaea9cee63b920478cb058f1;
reg  [MAX_SUM_WDTH_L-1:0]        Icdd2f6ce69b389fbf712e45bdc0a0257;
reg  [MAX_SUM_WDTH_L-1:0]        I8971b250393b397b94db38b9fd0fe501;
reg  [MAX_SUM_WDTH_L-1:0]        I9199e5e8fdc0e2c62ad1d62fc4d873cb;
reg  [MAX_SUM_WDTH_L-1:0]        I6e03f71fdf20db836c5772658a050e9c;
reg  [MAX_SUM_WDTH_L-1:0]        I2ef49f893dbc8581725ca0f6d1c3305c;
reg  [MAX_SUM_WDTH_L-1:0]        I8796f168c892ac60c38a0a7f1e18035e;
reg  [MAX_SUM_WDTH_L-1:0]        I64a26e5117c8f3ab95bf0dfa97427243;
reg  [MAX_SUM_WDTH_L-1:0]        Id7946a0299ced3ba00f6c3e6e664931f;
reg  [MAX_SUM_WDTH_L-1:0]        I5243b90640ea4680de83021601c85c39;
reg  [MAX_SUM_WDTH_L-1:0]        Ic8301fceed328cc031640ecc4ff34803;
reg  [MAX_SUM_WDTH_L-1:0]        I6e852c94b6105af62ee85f8adf77fa55;
reg  [MAX_SUM_WDTH_L-1:0]        I7d98c5c2a54832b6368ce60009208eb0;
reg  [MAX_SUM_WDTH_L-1:0]        I7e42f2281518bead81a6d18d2dcbd1a3;
reg  [MAX_SUM_WDTH_L-1:0]        I63c126c978154f2d68b11f08a938dcb4;
reg  [MAX_SUM_WDTH_L-1:0]        I2ff7719c35578b47720cacd9ddfd92eb;
reg  [MAX_SUM_WDTH_L-1:0]        I480599aef36967a670155dd77120a37d;
reg  [MAX_SUM_WDTH_L-1:0]        Ic000b2c844de484b8f30b7b84dd6234d;
reg  [MAX_SUM_WDTH_L-1:0]        If0e25df151db991185f992eab5d5be99;
reg  [MAX_SUM_WDTH_L-1:0]        I2f533699abb7a997160bf4ee4cda3efb;
reg  [MAX_SUM_WDTH_L-1:0]        If6b33cfc6d34e33fbb18e08fb4d8a5ed;
reg  [MAX_SUM_WDTH_L-1:0]        I2ea5423dc8726fc0217899e0f406a1e9;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf3f4f8a04cbacc9624ca5cc73bf7069;
reg  [MAX_SUM_WDTH_L-1:0]        I9ba53c36934ab1c7f498241a79cfbae8;
reg  [MAX_SUM_WDTH_L-1:0]        I106a25f18536f96782927bf3bc2ccd72;
reg  [MAX_SUM_WDTH_L-1:0]        Ie5cdad65e918679607cc5f816987b736;
reg  [MAX_SUM_WDTH_L-1:0]        Ica6dc9ded8756fd6f82eec4271e246c3;
reg  [MAX_SUM_WDTH_L-1:0]        Ica42ac6ca5813d0d1a67f14d1248437a;
reg  [MAX_SUM_WDTH_L-1:0]        I13dc6cfc75ef846c30e5dc1dc5305d59;
reg  [MAX_SUM_WDTH_L-1:0]        I33e784182dfb4af39715788b1ae98af6;
reg  [MAX_SUM_WDTH_L-1:0]        I9e1a66805348d2e5bbf5e2316187444b;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9619916a96d218cf5eb5f3a4995d0e7;
reg  [MAX_SUM_WDTH_L-1:0]        I02ce7969c51ad141df227ed7d18e74b1;
reg  [MAX_SUM_WDTH_L-1:0]        Idd73461af0d75c4d820f7f8f0f419e0f;
reg  [MAX_SUM_WDTH_L-1:0]        I3df6c2cdccb2a82c58c1d81b00af7786;
reg  [MAX_SUM_WDTH_L-1:0]        I97f441fc5ffb88efeb5ed66b60f07a7c;
reg  [MAX_SUM_WDTH_L-1:0]        I3194a235eb652c8d0e4307cd056e5e72;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc315f6c79ba2bf336ee57f2e5f7d776;
reg  [MAX_SUM_WDTH_L-1:0]        I937a54f5cda99a7079c7fa46b4ea26f6;
reg  [MAX_SUM_WDTH_L-1:0]        I49c99afecc613656cd1469d8c1e98936;
reg  [MAX_SUM_WDTH_L-1:0]        Id76ce0333f43bf7bccf1ce48e25ca69c;
reg  [MAX_SUM_WDTH_L-1:0]        I2c77f9644145219005751f7a4eb71aaa;
reg  [MAX_SUM_WDTH_L-1:0]        I5cecc266272eef88cda88c1df9bcc37e;
reg  [MAX_SUM_WDTH_L-1:0]        I776a0b1b5c14afa21b7fda3c2cacafed;
reg  [MAX_SUM_WDTH_L-1:0]        I84860b1f933339e0f90beeb3d666393b;
reg  [MAX_SUM_WDTH_L-1:0]        Id24581713f1ecb767db39d5154c2f5f4;
reg  [MAX_SUM_WDTH_L-1:0]        Idb0eae2f0e1dae1d56251d64e2c51f9f;
reg  [MAX_SUM_WDTH_L-1:0]        I2e3ca4b130e6d3d92385928a28644452;
reg  [MAX_SUM_WDTH_L-1:0]        I7922d80ae333dcfafde31d294f0eb4d8;
reg  [MAX_SUM_WDTH_L-1:0]        I82de04cd2dfef5616efca4af26d7c561;
reg  [MAX_SUM_WDTH_L-1:0]        I7ce384520525b15d24c2ef6f161213a5;
reg  [MAX_SUM_WDTH_L-1:0]        I56aeea71c7bd19d47620cf36adf3f115;
reg  [MAX_SUM_WDTH_L-1:0]        I138e1a6db0c6649bc023cc36d81d5b47;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5e8b1c4dd9b5dad56b59cc11c87a258;
reg  [MAX_SUM_WDTH_L-1:0]        I86f785e2d5e8d6c08fad1d334c7d244e;
reg  [MAX_SUM_WDTH_L-1:0]        I9a6c8efca218c724da4ee4c1087d58bc;
reg  [MAX_SUM_WDTH_L-1:0]        Ia30e8dbc6974ea94b763842e8dffa633;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa60f45f4d8848eb0b89f5644ec69668;
reg  [MAX_SUM_WDTH_L-1:0]        I0aeb4b93cfa6d62ec41b7e6dd0287dd0;
reg  [MAX_SUM_WDTH_L-1:0]        Ifce1fc978fb5b0187593f46f53c3b469;
reg  [MAX_SUM_WDTH_L-1:0]        If3b6de7c919c5d53a0e191a75bd7e574;
reg  [MAX_SUM_WDTH_L-1:0]        Iecce594e6e99b0c05fc845144a664b07;
reg  [MAX_SUM_WDTH_L-1:0]        I2c8431500ecb25619d2884a2fb4260c0;
reg  [MAX_SUM_WDTH_L-1:0]        I217c710f7ef39035546efcbb043f63f3;
reg  [MAX_SUM_WDTH_L-1:0]        I1b4236130cb1879d885653fdd9eeab4e;
reg  [MAX_SUM_WDTH_L-1:0]        Iae0f7c13f1564d63b4bfdc152ddf4111;
reg  [MAX_SUM_WDTH_L-1:0]        I010592496030d138a3a4245d00069957;
reg  [MAX_SUM_WDTH_L-1:0]        I9d7f47a6289a16448221d61f301586aa;
reg  [MAX_SUM_WDTH_L-1:0]        I7b8ed2953170c4deadaeb33a6ba165d4;
reg  [MAX_SUM_WDTH_L-1:0]        I4efe9eef6a48aeb0a9ba4e0ffd9906c3;
reg  [MAX_SUM_WDTH_L-1:0]        I5a8466bbd83c39dfbeaa6399e3fb3337;
reg  [MAX_SUM_WDTH_L-1:0]        I1ab96ffa948dd09bcc4f748c6c2575d2;
reg  [MAX_SUM_WDTH_L-1:0]        I016f57568eaf00b26f8a22100858c158;
reg  [MAX_SUM_WDTH_L-1:0]        I1fb995e302f4f1ba493ff85f39938175;
reg  [MAX_SUM_WDTH_L-1:0]        Ie643ad235307c60f1ee96dfdcbc8c2a8;
reg  [MAX_SUM_WDTH_L-1:0]        I8dafdf2c780082d8dfc2961b3447f104;
reg  [MAX_SUM_WDTH_L-1:0]        I3a2841a0f5e1b42556f384231ab0717b;
reg  [MAX_SUM_WDTH_L-1:0]        I2b00d0e6facf01274c0c3446bb0e1599;
reg  [MAX_SUM_WDTH_L-1:0]        I2c645d25871b70dae5b2c283695d5130;
reg  [MAX_SUM_WDTH_L-1:0]        I540a0e8968a6a82aca775a81ef82b520;
reg  [MAX_SUM_WDTH_L-1:0]        I5b95bbc82e6d8d87421efe3f17b97ea5;
reg  [MAX_SUM_WDTH_L-1:0]        Iad81f5e5e728ffdec6296b2aff668d75;
reg  [MAX_SUM_WDTH_L-1:0]        I960a618f63372da74581b8c352f3e618;
reg  [MAX_SUM_WDTH_L-1:0]        I4f5325f1601acde10018d1fd0aff4d35;
reg  [MAX_SUM_WDTH_L-1:0]        Ib297101fe456520e72cd9d208af44eea;
reg  [MAX_SUM_WDTH_L-1:0]        I73a21342321a9d81a0fa5308149d72b0;
reg  [MAX_SUM_WDTH_L-1:0]        I2a486524f4f53b3454ee02a8892d4fa3;
reg  [MAX_SUM_WDTH_L-1:0]        Ic6c4e4e6a9ba43a3354f9f3192ab069e;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3cdee3560bd06aed84dac5fcd2a259a;
reg  [MAX_SUM_WDTH_L-1:0]        I584febaa4c440fd9353108af36d3a5c6;
reg  [MAX_SUM_WDTH_L-1:0]        I515e78507d7419ca14d77b6d52f75a78;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9578453a57d2b3b9c3b98844044b5f0;
reg  [MAX_SUM_WDTH_L-1:0]        I1e58b3062097a46d8d590232b40278cf;
reg  [MAX_SUM_WDTH_L-1:0]        I3af126eb28c67797ce625b0d82943833;
reg  [MAX_SUM_WDTH_L-1:0]        I130ee1a8acacf4cae8818cd8320d050d;
reg  [MAX_SUM_WDTH_L-1:0]        Idf92dd09c29ce8e921b2b34089550586;
reg  [MAX_SUM_WDTH_L-1:0]        Iba74a64cc1d2ec3c83a4061db298ad37;
reg  [MAX_SUM_WDTH_L-1:0]        I01364c233ca541914d790354515aa5c1;
reg  [MAX_SUM_WDTH_L-1:0]        Ic6a8297308a63ed3113008a3cdc76358;
reg  [MAX_SUM_WDTH_L-1:0]        I6c7ee9d0bd684a7f54bed3d52452219d;
reg  [MAX_SUM_WDTH_L-1:0]        I985ea87550ec8a222e6af621589e186d;
reg  [MAX_SUM_WDTH_L-1:0]        I6836a7d1e006d7f7556edf8b31aea32e;
reg  [MAX_SUM_WDTH_L-1:0]        Ia7a356a18af18ec131b9df46019f3e58;
reg  [MAX_SUM_WDTH_L-1:0]        If3a7e111247232c47ceccb5e05338312;
reg  [MAX_SUM_WDTH_L-1:0]        I5f38d1665294b2d3c18f9cd888ff60f1;
reg  [MAX_SUM_WDTH_L-1:0]        I10290b9576bf3d8caf90583a388226b7;
reg  [MAX_SUM_WDTH_L-1:0]        Ief36236305fc1521c5bb4c60753a676a;
reg  [MAX_SUM_WDTH_L-1:0]        Ibaa0539fbf5ccc979511c09c061cf494;
reg  [MAX_SUM_WDTH_L-1:0]        I95664ffd0ff13c2893421032149f24d2;
reg  [MAX_SUM_WDTH_L-1:0]        Ie390153b3b7985dc63d65913de215377;
reg  [MAX_SUM_WDTH_L-1:0]        I704147dda658f4a03627dacc1c91dd48;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb09672d505898f081aa13c95fcb88b5;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb5cb89097dd11bf292d5b5a2422175b;
reg  [MAX_SUM_WDTH_L-1:0]        I4a305956b18d6ad6901d2c17e99f2bab;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf5bb3b9eb1812383db9634fa9a27ad3;
reg  [MAX_SUM_WDTH_L-1:0]        I66b37d055c3735f011095ee4b1ad02ed;
reg  [MAX_SUM_WDTH_L-1:0]        I43e71dd694d97217e242f267248cd594;
reg  [MAX_SUM_WDTH_L-1:0]        I4baa925db1ec733bd4bd25d9dc873e23;
reg  [MAX_SUM_WDTH_L-1:0]        I547928c9db7acc531af251264d576ffb;
reg  [MAX_SUM_WDTH_L-1:0]        Ie4ce634b2fb62a20781f8a2e8fddc762;
reg  [MAX_SUM_WDTH_L-1:0]        I0e90e96ffa64c2874d79110b622994bf;
reg  [MAX_SUM_WDTH_L-1:0]        I767e37e3c6f4224eb07adeda480ce253;
reg  [MAX_SUM_WDTH_L-1:0]        I75fcaf2c65b7e63adac834054850c6d6;
reg  [MAX_SUM_WDTH_L-1:0]        I5f1de2dfbd79204ab2db9b686d6a6862;
reg  [MAX_SUM_WDTH_L-1:0]        I8d01de6be4091dca2589cef625c05229;
reg  [MAX_SUM_WDTH_L-1:0]        Ic09e773899fdd208c0fdd874933b2cec;
reg  [MAX_SUM_WDTH_L-1:0]        I24a3f9fd851c4af70ef66bfcee44af65;
reg  [MAX_SUM_WDTH_L-1:0]        Idd31807ecd603db8c719349a2be1be40;
reg  [MAX_SUM_WDTH_L-1:0]        Iaf680cae40d1adf7649da12b31a2be0d;
reg  [MAX_SUM_WDTH_L-1:0]        I22d948171c1a66f7a28d5e51007700ea;
reg  [MAX_SUM_WDTH_L-1:0]        I3954318b2392a82f2da71a0ca1504497;
reg  [MAX_SUM_WDTH_L-1:0]        I15c78b909cbd04fe25820d777655d829;
reg  [MAX_SUM_WDTH_L-1:0]        Ia529c5ec88a9f6c14ceda5cad56b346d;
reg  [MAX_SUM_WDTH_L-1:0]        I5b73c81f28901705f6ee26d63847db0a;
reg  [MAX_SUM_WDTH_L-1:0]        I1a9bd3f728db23b679639e5657ced179;
reg  [MAX_SUM_WDTH_L-1:0]        I57ca72784a7c91cecbd694ddd08bcb98;
reg  [MAX_SUM_WDTH_L-1:0]        I50f31ecd3f2b498cc7b759efa057f12f;
reg  [MAX_SUM_WDTH_L-1:0]        I8ccaf29848defdd264f522642968fa29;
reg  [MAX_SUM_WDTH_L-1:0]        I808ea92ee1340876cf1d2c47255dc2fe;
reg  [MAX_SUM_WDTH_L-1:0]        I3da806790125328b626be1949f71267a;
reg  [MAX_SUM_WDTH_L-1:0]        I55e59bc1daeb8b2be3d7a1e4b272df93;
reg  [MAX_SUM_WDTH_L-1:0]        Ib0ffadc6a0091ceff91ad1fa435413a6;
reg  [MAX_SUM_WDTH_L-1:0]        Ic863f139e6bed2d06789a07c6dedf6f8;
reg  [MAX_SUM_WDTH_L-1:0]        Id0e8f6ada5060a911090f76cfaa3c6bf;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb8c9b8fc9b58f5f8a6ad342934804a8;
reg  [MAX_SUM_WDTH_L-1:0]        I9323a188737ca54c2dd553cd99bd416c;
reg  [MAX_SUM_WDTH_L-1:0]        I2694cef38855f496e7ca12f42dfdb9fc;
reg  [MAX_SUM_WDTH_L-1:0]        I75790b4c0b1f6c7935f5cfbea26407d1;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8b366c47e56a49fc53ea4a9e1ebbd99;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1c86256df2bc6c4dad41237eca41986;
reg  [MAX_SUM_WDTH_L-1:0]        I7c9e3f97a94f9a078c209a1b84ff916d;
reg  [MAX_SUM_WDTH_L-1:0]        Idde839d34403fdbba62671b83801ea8d;
reg  [MAX_SUM_WDTH_L-1:0]        I824e23c3e43434e0a7bf8c8b8e0de597;
reg  [MAX_SUM_WDTH_L-1:0]        I0f83a2c488c229e971030fc66ce212f5;
reg  [MAX_SUM_WDTH_L-1:0]        I8fdda3dea7a63fd6e57f70365d7b6571;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa2fc30c14c549339edc65c3670d90a0;
reg  [MAX_SUM_WDTH_L-1:0]        If69bb1bfa10ca7dd37ba57485c3429e7;
reg  [MAX_SUM_WDTH_L-1:0]        I2ab0738fa2d5916d77a81b9da2315376;
reg  [MAX_SUM_WDTH_L-1:0]        I50a9ce776ad2ccd8048b56ce101c80d2;
reg  [MAX_SUM_WDTH_L-1:0]        I9c9d0332ee7ad6a3488b7e39bcb06ca2;
reg  [MAX_SUM_WDTH_L-1:0]        Idc155814976f0aef9b56b2bb3d52b3a5;
reg  [MAX_SUM_WDTH_L-1:0]        I2e02fbd496d08acb3ad3359b49b9f680;
reg  [MAX_SUM_WDTH_L-1:0]        If0f8b3dfce99a5a75c2105d45ccad985;
reg  [MAX_SUM_WDTH_L-1:0]        I6790223e6a7cf136a7e2b261ba4fdb0a;
reg  [MAX_SUM_WDTH_L-1:0]        I6a9643afea7a6cc9b94806ccc8e84c0f;
reg  [MAX_SUM_WDTH_L-1:0]        Id3d19d7c2b941930478a7ab01049e390;
reg  [MAX_SUM_WDTH_L-1:0]        Ib0a25312d51cb6aa1741f7e425bc5cd8;
reg  [MAX_SUM_WDTH_L-1:0]        I44dd1b66f5a9a6b0b976d3d61d6c5cbe;
reg  [MAX_SUM_WDTH_L-1:0]        I3ee456f2f0e7f447ae92b7523136adb5;
reg  [MAX_SUM_WDTH_L-1:0]        Ic110e2a08b550acd3c8bda4a1bc2bbae;
reg  [MAX_SUM_WDTH_L-1:0]        I3f87162d2874effd66a82f821aa6c73a;
reg  [MAX_SUM_WDTH_L-1:0]        I660ea6d341fcb38f108270c08d82473b;
reg  [MAX_SUM_WDTH_L-1:0]        Ic128d603fc08affd2f3d0ab3425710e5;
reg  [MAX_SUM_WDTH_L-1:0]        Id5372641727970383a59e08f550814b4;
reg  [MAX_SUM_WDTH_L-1:0]        Ie99ad992d66880542dcd330ef6ccee04;
reg  [MAX_SUM_WDTH_L-1:0]        I9ed0b194f7d210d57c54b289e01c75e6;
reg  [MAX_SUM_WDTH_L-1:0]        I227828831c4ad21b06ed00fb5781b0e3;
reg  [MAX_SUM_WDTH_L-1:0]        I09d5ad12cb836adfbb4833ee80fad2c9;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa9c94ee94e4beb2e7c8d2d57150df41;
reg  [MAX_SUM_WDTH_L-1:0]        Icb88e59e194db215382e8e949603a9be;
reg  [MAX_SUM_WDTH_L-1:0]        Id4ebd28aaf1076acec266666f88a02ad;
reg  [MAX_SUM_WDTH_L-1:0]        Idf0a0bd862167392357501b3233a8d8c;
reg  [MAX_SUM_WDTH_L-1:0]        If94cdb867ea0fc2c5578b16aacb1acfc;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8c066b0700941a4fa739820ff12b948;
reg  [MAX_SUM_WDTH_L-1:0]        I11e0f8dc46b286bafb05f901f968e1ad;
reg  [MAX_SUM_WDTH_L-1:0]        I608537f5639d5e0cd3e80453e21f6f85;
reg  [MAX_SUM_WDTH_L-1:0]        I0e9d8db1bb6347c9507b645132308b3a;
reg  [MAX_SUM_WDTH_L-1:0]        I17033b417fa383a2db41d157df33d9de;
reg  [MAX_SUM_WDTH_L-1:0]        Ib7f45dbcad513b4dafee60f33622b0c3;
reg  [MAX_SUM_WDTH_L-1:0]        Ibfbd8e00e00272f32428c7b4a3c53050;
reg  [MAX_SUM_WDTH_L-1:0]        I27973d1d4e07eaa49608d6f6975d0a93;
reg  [MAX_SUM_WDTH_L-1:0]        If77fcedbcf99f89045de87e5cae45d8a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8f8691820e7a560db8116f38dae5d49;
reg  [MAX_SUM_WDTH_L-1:0]        If0b19af59ad851aded19970494514034;
reg  [MAX_SUM_WDTH_L-1:0]        I98b8e05818925a4b65082fa57affde83;
reg  [MAX_SUM_WDTH_L-1:0]        I69317e8c556ed67630829c990f8b74db;
reg  [MAX_SUM_WDTH_L-1:0]        I9147d103cf235310393f9339f1cbb376;
reg  [MAX_SUM_WDTH_L-1:0]        Ibe0b2cab6e2d3f3cc8baf3623ff50988;
reg  [MAX_SUM_WDTH_L-1:0]        Idc64f1443dd2497dfaa223cda3fbd682;
reg  [MAX_SUM_WDTH_L-1:0]        I6e37e92b812099985436851da8a6ccb2;
reg  [MAX_SUM_WDTH_L-1:0]        I057df2bf67d5580275654bdc28b40027;
reg  [MAX_SUM_WDTH_L-1:0]        Ie87a151c8b90942a899b8167bcb34afb;
reg  [MAX_SUM_WDTH_L-1:0]        I735752035af159b48f53d8302bb33c21;
reg  [MAX_SUM_WDTH_L-1:0]        I1f26bc7cb30a9659a638e2ab65e1f187;
reg  [MAX_SUM_WDTH_L-1:0]        If39a50e88c4a7c43428c1d15b0bfbbcc;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf966c12f049d603361ad32f55b0a2c8;
reg  [MAX_SUM_WDTH_L-1:0]        Ie1b3ed6d3fdae47669d3c4cb8af8d969;
reg  [MAX_SUM_WDTH_L-1:0]        I4ec6c8d9e87224ecbe7c69d92f9419c8;
reg  [MAX_SUM_WDTH_L-1:0]        I2acb34de8c3fc53117a7ea4f9ce7dd2b;
reg  [MAX_SUM_WDTH_L-1:0]        I7fa4009267e80ea7eb71194843c3b22b;
reg  [MAX_SUM_WDTH_L-1:0]        I6854329daadea2734e52180a41f56bcc;
reg  [MAX_SUM_WDTH_L-1:0]        Ifca16aebaf75b2990188de201e4536fd;
reg  [MAX_SUM_WDTH_L-1:0]        I46cc26afc8475f2fb290eefc95a542eb;
reg  [MAX_SUM_WDTH_L-1:0]        Id746d6515cec9e60e7478898a09787e5;
reg  [MAX_SUM_WDTH_L-1:0]        I09a3ad636db96e00adac78c3c94bdaaa;
reg  [MAX_SUM_WDTH_L-1:0]        I28b3baa225a5fd602c9fee9c948ae58b;
reg  [MAX_SUM_WDTH_L-1:0]        Ibe12ef0f56d875c7a44030882deb0e29;
reg  [MAX_SUM_WDTH_L-1:0]        I9bd9979e4acc4944227a4bd62b910c1d;
reg  [MAX_SUM_WDTH_L-1:0]        Idcfa802f458499150055dbe4b1ce8146;
reg  [MAX_SUM_WDTH_L-1:0]        Iee010958cc3e9389cb8ecacff84fccee;
reg  [MAX_SUM_WDTH_L-1:0]        I3d74b31096917c53757c829a67cf06df;
reg  [MAX_SUM_WDTH_L-1:0]        Ic27031a9654db9459815fe0ca35408db;
reg  [MAX_SUM_WDTH_L-1:0]        Idf6ead2c37f75f3cde1d4b40cd73db00;
reg  [MAX_SUM_WDTH_L-1:0]        I66a56161cd0ed67f65834b9eb0e94d17;
reg  [MAX_SUM_WDTH_L-1:0]        If6de990e26ca9e8efc009188f8a5a4d9;
reg  [MAX_SUM_WDTH_L-1:0]        I8d866786bb2dea06f5b30f6ea80cff17;
reg  [MAX_SUM_WDTH_L-1:0]        I01ca9a1d4901ec9b2a64300617ce4cd1;
reg  [MAX_SUM_WDTH_L-1:0]        I2dbead35e15afb9affaa6ad4edd3829e;
reg  [MAX_SUM_WDTH_L-1:0]        I83c57653e24cc09214075b04b06bad83;
reg  [MAX_SUM_WDTH_L-1:0]        I56b9c1f555b24c2dc197168decfdb8d1;
reg  [MAX_SUM_WDTH_L-1:0]        Id5c48111f1b93de2cfe89f92fd182b43;
reg  [MAX_SUM_WDTH_L-1:0]        I32908c3c90ed6488357ce4869e8a1721;
reg  [MAX_SUM_WDTH_L-1:0]        I16b4601f2e07e6cecdb5a030178e75c0;
reg  [MAX_SUM_WDTH_L-1:0]        I0ae08a41ebd0e6b402a4980478087bb5;
reg  [MAX_SUM_WDTH_L-1:0]        Icb57267a66f117943e964dd6420d7a58;
reg  [MAX_SUM_WDTH_L-1:0]        Icfa47fb87b74106cd3814adfce909424;
reg  [MAX_SUM_WDTH_L-1:0]        I63067cef0e1a348a3e6d8cd9bd88b907;
reg  [MAX_SUM_WDTH_L-1:0]        I10aa5ba0f53632578c0e1cefa4bf4fde;
reg  [MAX_SUM_WDTH_L-1:0]        I427c0215d0ac047e8402c20610676752;
reg  [MAX_SUM_WDTH_L-1:0]        Icf4efa87688bd1b80437686eb0126057;
reg  [MAX_SUM_WDTH_L-1:0]        Ic373f785ddd1bf8eccce263df5a82c87;
reg  [MAX_SUM_WDTH_L-1:0]        I56f8e8d2d7052af26528530d389b6dc1;
reg  [MAX_SUM_WDTH_L-1:0]        Ifb145bc18d435fb66779e7415417bc0f;
reg  [MAX_SUM_WDTH_L-1:0]        I62a6e0c9952d6c6e6095e2364df93078;
reg  [MAX_SUM_WDTH_L-1:0]        Id6405c2b2b9aea6bc457f1064d5f3ffa;
reg  [MAX_SUM_WDTH_L-1:0]        I079df9611bd81f672f2ae028bf267995;
reg  [MAX_SUM_WDTH_L-1:0]        I096b226cc511363946a39307a7d97867;
reg  [MAX_SUM_WDTH_L-1:0]        I4cc42c5a75ef339510ee0e86fb44e16a;
reg  [MAX_SUM_WDTH_L-1:0]        I680c01c3327cb9372a42c1ec5b4193e3;
reg  [MAX_SUM_WDTH_L-1:0]        I83451a072082194ecb3f9419edd728b3;
reg  [MAX_SUM_WDTH_L-1:0]        I52ad85b6a1c822ca8c2459bde8fbd510;
reg  [MAX_SUM_WDTH_L-1:0]        I1c44d2ef638825862061a8ee1a0a2f95;
reg  [MAX_SUM_WDTH_L-1:0]        I8fa1fd425809cc39cd8e2785773c1d7a;
reg  [MAX_SUM_WDTH_L-1:0]        Ifa22335f04d35680eb8cfec8f862f357;
reg  [MAX_SUM_WDTH_L-1:0]        I6aff673c27811b81530453906312aa9c;
reg  [MAX_SUM_WDTH_L-1:0]        If674ac0540f457a21235664c213d4923;
reg  [MAX_SUM_WDTH_L-1:0]        Iac223ac498bdcf2cb2514582aeaf76f3;
reg  [MAX_SUM_WDTH_L-1:0]        I7f40931ab78ededfcb52ccaac9b81282;
reg  [MAX_SUM_WDTH_L-1:0]        Iab7c8dad0ca20eb0988fbd99f25591a8;
reg  [MAX_SUM_WDTH_L-1:0]        I3cb5f890a5bd3daaae34c8dfb6ecfc49;
reg  [MAX_SUM_WDTH_L-1:0]        Id80e145586d7e539a6514dd67ebabf6a;
reg  [MAX_SUM_WDTH_L-1:0]        I01e09bc554768f30dc490041d19b4da2;
reg  [MAX_SUM_WDTH_L-1:0]        I0196f7df6f834ae20c4fdd127e66104d;
reg  [MAX_SUM_WDTH_L-1:0]        I4669c4f256c123a0fcceb55c1e72193a;
reg  [MAX_SUM_WDTH_L-1:0]        I4a02ffa2a79df824f406909aa189a404;
reg  [MAX_SUM_WDTH_L-1:0]        I3117e5029119e70846dff61d746699e7;
reg  [MAX_SUM_WDTH_L-1:0]        I1e4e705b3bda1451fc384cd934c0bb52;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5bea8e0072de3de2c8431ea6a35dd51;
reg  [MAX_SUM_WDTH_L-1:0]        I7d9d94022ea95ea01cddc237f3df8cb8;
reg  [MAX_SUM_WDTH_L-1:0]        I3f0f9aab07427fa81fc3096c6b6d3d6d;
reg  [MAX_SUM_WDTH_L-1:0]        I12a7983041f9c298d533bad58f41d24b;
reg  [MAX_SUM_WDTH_L-1:0]        I78503880e5c96ec0a03c75266b1226e8;
reg  [MAX_SUM_WDTH_L-1:0]        I8adeae445b33f634977957bb1a2259aa;
reg  [MAX_SUM_WDTH_L-1:0]        I73bd13f381d15e0b0198b60cee44bb42;
reg  [MAX_SUM_WDTH_L-1:0]        Ic8b651c2b043a4a6e4cd259774322230;
reg  [MAX_SUM_WDTH_L-1:0]        I76979d7df582f9306e796a03cb540963;
reg  [MAX_SUM_WDTH_L-1:0]        If61d4585986757a525c54589ec93d8c6;
reg  [MAX_SUM_WDTH_L-1:0]        I1bc5766a4a3cc2b468ab8ef62eab691c;
reg  [MAX_SUM_WDTH_L-1:0]        I21585169e5fceda643bd03fddf8153be;
reg  [MAX_SUM_WDTH_L-1:0]        Idb2990946f60939136b3bfddbc7b1671;
reg  [MAX_SUM_WDTH_L-1:0]        Icfbf703890f684bfc96decc429deaa04;
reg  [MAX_SUM_WDTH_L-1:0]        Id5bb42639a1c1c1d67df1c89a14a2bfc;
reg  [MAX_SUM_WDTH_L-1:0]        I55b8ef91d667c1c1d9e58dbc86a2288a;
reg  [MAX_SUM_WDTH_L-1:0]        I17ff683da41b469c8c8b82ee32a7378a;
reg  [MAX_SUM_WDTH_L-1:0]        I51f10296c38872338ec7df35ccd520d8;
reg  [MAX_SUM_WDTH_L-1:0]        Ia59ff33765ddf4aeb17f90a70c01d76c;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf97abffb1ec40f2f0e099a814e04ab2;
reg  [MAX_SUM_WDTH_L-1:0]        I3efc3271e18a1e350473dcf3375088aa;
reg  [MAX_SUM_WDTH_L-1:0]        I1efd1220ea9100f2fb4f169ceaf462a5;
reg  [MAX_SUM_WDTH_L-1:0]        I9af399f27c8e2b62b7f3fc6481ef9318;
reg  [MAX_SUM_WDTH_L-1:0]        I171bb4ee9be2f92e4d82997108572426;
reg  [MAX_SUM_WDTH_L-1:0]        Ib13cd76c20fcaf95f26f4914380c4fcf;
reg  [MAX_SUM_WDTH_L-1:0]        Iafb219f1c8c6883e01fbfb4c887c8d6a;
reg  [MAX_SUM_WDTH_L-1:0]        I94fc9b0bdd2b0a89a9f6351f1fdd4ff5;
reg  [MAX_SUM_WDTH_L-1:0]        Ia9ceb45f33402293c162cef4037ba007;
reg  [MAX_SUM_WDTH_L-1:0]        I0fa4e12e62e8a30b3b8045143b344b4f;
reg  [MAX_SUM_WDTH_L-1:0]        Icec1c637d24ca277bb2e488257e92a40;
reg  [MAX_SUM_WDTH_L-1:0]        Ie9aca08b988fad20904545fe070defd5;
reg  [MAX_SUM_WDTH_L-1:0]        Ie82304b2c8583f967649475e309e68fa;
reg  [MAX_SUM_WDTH_L-1:0]        I60da0fb8a2c0669d5f9037ae99b23565;
reg  [MAX_SUM_WDTH_L-1:0]        Id8c19a3547c17ed513d2d857adc66885;
reg  [MAX_SUM_WDTH_L-1:0]        Id74984743844e9495ea0f528a391f4b8;
reg  [MAX_SUM_WDTH_L-1:0]        I9edcdd5b927b3f6b3a4c7cacebeb4a82;
reg  [MAX_SUM_WDTH_L-1:0]        Ic89597a95f50382cd3a2730896735d55;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb7d203dfc75bf6211b09ab94877f93d;
reg  [MAX_SUM_WDTH_L-1:0]        Id2f2e6837c83973cb2173454433acb88;
reg  [MAX_SUM_WDTH_L-1:0]        I1259d5918f8d65b4b22ccfef22fe3afa;
reg  [MAX_SUM_WDTH_L-1:0]        Ib84e8c6e7fd9d7762e6e7e508d5ee40a;
reg  [MAX_SUM_WDTH_L-1:0]        Ia032017912715abde99ffdf5ba732c5f;
reg  [MAX_SUM_WDTH_L-1:0]        I55c310bfefb635448ef9c25c5d15987e;
reg  [MAX_SUM_WDTH_L-1:0]        I92c0f229cf7fdb2cc0fe4d84f4d9b11d;
reg  [MAX_SUM_WDTH_L-1:0]        I5570eb486d238fd96f9a59b174f5a22a;
reg  [MAX_SUM_WDTH_L-1:0]        If6f01d24acf4a8b38bdbb1b366cd9a47;
reg  [MAX_SUM_WDTH_L-1:0]        Iff29fff36064aa4f9d339d4c62956e61;
reg  [MAX_SUM_WDTH_L-1:0]        I818d7cae6f1b80ac452dbfc073ccfe7a;
reg  [MAX_SUM_WDTH_L-1:0]        I77ecfe991c6ec778495d7d5e5e442eca;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7c6a56e8b6f7756bb5a24bdfd6a855e;
reg  [MAX_SUM_WDTH_L-1:0]        I9f9bc8eb8b2978a3dc529c34516fdf75;
reg  [MAX_SUM_WDTH_L-1:0]        Ie3c0e5a4b00a92357a5d37e527d59b61;
reg  [MAX_SUM_WDTH_L-1:0]        I9b9a9486420e7d4aa105c48dd50aa74d;
reg  [MAX_SUM_WDTH_L-1:0]        Id12199a504f7aa298fffaaedd1aacc99;
reg  [MAX_SUM_WDTH_L-1:0]        I813691fd8ea36626d32c8d2562163f32;
reg  [MAX_SUM_WDTH_L-1:0]        I5fd3aaddc3eb8afeb82768b45e2d53d7;
reg  [MAX_SUM_WDTH_L-1:0]        I1ac281eab6c7459e835fe992142b7857;
reg  [MAX_SUM_WDTH_L-1:0]        I49e5078c9161e8bee00fb76bc00b5288;
reg  [MAX_SUM_WDTH_L-1:0]        Ia697adf14616bf50d6e8178596b9fa7e;
reg  [MAX_SUM_WDTH_L-1:0]        Iff3128a26dabe63b015dc6afc98a85a9;
reg  [MAX_SUM_WDTH_L-1:0]        Ifc04708ee5a7cc2b3f1850db778fa42e;
reg  [MAX_SUM_WDTH_L-1:0]        Ia405859c9dff67905b2e91bcbc06259e;
reg  [MAX_SUM_WDTH_L-1:0]        I2fec8f62b28575e8f3af756db66fa232;
reg  [MAX_SUM_WDTH_L-1:0]        I98e97c02477032ead66dc50f3f274e5a;
reg  [MAX_SUM_WDTH_L-1:0]        I9f2dc5add3a4d1e6eb3116c741cd2f82;
reg  [MAX_SUM_WDTH_L-1:0]        Ie122f7d8a48d7ad29d998b6a14b8e70f;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5576c996062391f44066d893dd5cb91;
reg  [MAX_SUM_WDTH_L-1:0]        If931597aab866a74c3a3ffb1cd429583;
reg  [MAX_SUM_WDTH_L-1:0]        I79878bd69ed53785b8a5f025a2a00a4f;
reg  [MAX_SUM_WDTH_L-1:0]        Iefb0a20652954fc2002154ea874c120a;
reg  [MAX_SUM_WDTH_L-1:0]        I646ca66e4e9f24b4fb75b38bf293b4cc;
reg  [MAX_SUM_WDTH_L-1:0]        I051f0d4c44123e3637b84a32c9a00a75;
reg  [MAX_SUM_WDTH_L-1:0]        I1876f9ec3f6f637ee40cdad7cc347f6f;
reg  [MAX_SUM_WDTH_L-1:0]        Ic3d6b8dbec6cf92a9b6a17fb2f75dcd4;
reg  [MAX_SUM_WDTH_L-1:0]        I7d89f1db7b1015d34363ad781374de58;
reg  [MAX_SUM_WDTH_L-1:0]        Ife217ec4da1f1477bce034cb3545160f;
reg  [MAX_SUM_WDTH_L-1:0]        Idc5e5e98508c94b87a760f8eb36fad41;
reg  [MAX_SUM_WDTH_L-1:0]        I9e72b0c823f297535f13a1b3072c2776;
reg  [MAX_SUM_WDTH_L-1:0]        Ia81da7c58d6636ab70e0cf3e263a12c0;
reg  [MAX_SUM_WDTH_L-1:0]        Ibfc69ef08382c79e30cfafd89bfeff69;
reg  [MAX_SUM_WDTH_L-1:0]        I2d2afa9165b7121dc8289e9e6cdab5de;
reg  [MAX_SUM_WDTH_L-1:0]        I065052693fd8ca87614feb60f7ef37c3;
reg  [MAX_SUM_WDTH_L-1:0]        I13344a81551374f665cbc17c7e94296a;
reg  [MAX_SUM_WDTH_L-1:0]        If5a1d2de0715fa87d191ee5f48171676;
reg  [MAX_SUM_WDTH_L-1:0]        I02b256f74ee86b42ff1eba5e3d242737;
reg  [MAX_SUM_WDTH_L-1:0]        Ic113fc051eefaef846f440e98f2f8913;
reg  [MAX_SUM_WDTH_L-1:0]        Iabeab9bdd0bd82dd145218b563b5dac1;
reg  [MAX_SUM_WDTH_L-1:0]        If9ce0a09e3a4e816dda002a24319ac0b;
reg  [MAX_SUM_WDTH_L-1:0]        Ib5a7d72c36e41754033a64fbe0718784;
reg  [MAX_SUM_WDTH_L-1:0]        I41df12c7dee8526abf92b8e98965fa06;
reg  [MAX_SUM_WDTH_L-1:0]        I83dfbd224e7465a6fd769e407182829a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie57bba5092ec318456365b81b36aaa65;
reg  [MAX_SUM_WDTH_L-1:0]        Ibcf043d24474ab8c1002d15fde2d7da2;
reg  [MAX_SUM_WDTH_L-1:0]        I2e3385871c6ed8cf9519f273c8a19fda;
reg  [MAX_SUM_WDTH_L-1:0]        I664917b9f44515bf556d69ade4ca408c;
reg  [MAX_SUM_WDTH_L-1:0]        I28deacdec0fbd0bce49b654c2620ac38;
reg  [MAX_SUM_WDTH_L-1:0]        Ibdfc4852c620f573f929584e6b816f35;
reg  [MAX_SUM_WDTH_L-1:0]        I5a69b2bbb63ab919ea2270503cd326f1;
reg  [MAX_SUM_WDTH_L-1:0]        I2eccd8d60a19481fa595566f51c7aa4e;
reg  [MAX_SUM_WDTH_L-1:0]        I49eb4bba42440657fe04b711eedfa67f;
reg  [MAX_SUM_WDTH_L-1:0]        I9ed8323951af0de78ae89153cbf9e9eb;
reg  [MAX_SUM_WDTH_L-1:0]        I1d00816529836546b514f54b1275d39e;
reg  [MAX_SUM_WDTH_L-1:0]        Icc58b9a24fb9ef7e8fa5f13a2cc0a0cb;
reg  [MAX_SUM_WDTH_L-1:0]        I9339aef608b029175b488e82f5b3f1bb;
reg  [MAX_SUM_WDTH_L-1:0]        Ibd2f24860b701ab46e0c436d774e43f9;
reg  [MAX_SUM_WDTH_L-1:0]        I37fe66ec8927f27f646b304500400ccf;
reg  [MAX_SUM_WDTH_L-1:0]        I4bd6a48f494cf633a857b8ccbd67af68;
reg  [MAX_SUM_WDTH_L-1:0]        Icd7a7566438dc67e77f138ac814844f0;
reg  [MAX_SUM_WDTH_L-1:0]        Ic3d4239413333883dd926c7a42c0a87f;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8298d1ead61bc00eb31599b3087d769;
reg  [MAX_SUM_WDTH_L-1:0]        I23dbe33ce46f94d3dff1e6d391305609;
reg  [MAX_SUM_WDTH_L-1:0]        I138286817f424c76e8a4f30540b0530b;
reg  [MAX_SUM_WDTH_L-1:0]        I30c645a78b900306864a1ab23e923bde;
reg  [MAX_SUM_WDTH_L-1:0]        Id88681d0fe3ea62530166938503db05a;
reg  [MAX_SUM_WDTH_L-1:0]        I808008402174fa4edf42783135c0c3a9;
reg  [MAX_SUM_WDTH_L-1:0]        I3ad4d02ea2e52a49b6fa4f1da9b58149;
reg  [MAX_SUM_WDTH_L-1:0]        I39486eecb7bbfecf26573a7a5876feb9;
reg  [MAX_SUM_WDTH_L-1:0]        I21e8ea20029fb2cb62103405b81b21b0;
reg  [MAX_SUM_WDTH_L-1:0]        Id0b67fa451e276889e02779ddb667904;
reg  [MAX_SUM_WDTH_L-1:0]        Ic328d25a58ec4559b753da3bcff938de;
reg  [MAX_SUM_WDTH_L-1:0]        I49c44c2f2522e086c2db8a00647ba35c;
reg  [MAX_SUM_WDTH_L-1:0]        Id4152a04385391294f4b8a18df2cb9ee;
reg  [MAX_SUM_WDTH_L-1:0]        I5b0213a3df61e94fd0b744a8141f7502;
reg  [MAX_SUM_WDTH_L-1:0]        If0ad11ed403cbbed68614b01e2a3793e;
reg  [MAX_SUM_WDTH_L-1:0]        Icfa1170bc73534bee13778bc3b88a2f7;
reg  [MAX_SUM_WDTH_L-1:0]        Ife1bd938a0dd06d8d3cf30ff41a303b2;
reg  [MAX_SUM_WDTH_L-1:0]        I4a09cb1b99b476fa6fae0bc44c41a041;
reg  [MAX_SUM_WDTH_L-1:0]        Ie08cf323944813e4b9e2d59a680ffe8d;
reg  [MAX_SUM_WDTH_L-1:0]        I85fc307fb52d58550eeecd33bc4207a4;
reg  [MAX_SUM_WDTH_L-1:0]        Id00dd13741fe621d0a240bdc92318f55;
reg  [MAX_SUM_WDTH_L-1:0]        Idc8e891fd432df75a4eb133ce35ecec4;
reg  [MAX_SUM_WDTH_L-1:0]        I2a51cada20cbd14f7d5a289599e68b53;
reg  [MAX_SUM_WDTH_L-1:0]        I65a701d1e083e501544bb0fce24f0c4e;
reg  [MAX_SUM_WDTH_L-1:0]        If3020a9109ac83274b5bafac18d176de;
reg  [MAX_SUM_WDTH_L-1:0]        Iaa6bd55038c2ae911e4df08f707c55f5;
reg  [MAX_SUM_WDTH_L-1:0]        Id49065cedf20e13abac8971534bb8b0e;
reg  [MAX_SUM_WDTH_L-1:0]        I0bb64952d77b59803a561e14b950b9b1;
reg  [MAX_SUM_WDTH_L-1:0]        I01e295a6ab88c6f34b44efcc32a23233;
reg  [MAX_SUM_WDTH_L-1:0]        I2acf864d587b7681ca0fb6e2e2bea617;
reg  [MAX_SUM_WDTH_L-1:0]        Idfd0410b37713e8808f8bea81e2af881;
reg  [MAX_SUM_WDTH_L-1:0]        I02861f333b5adfd4962356cdf5a11f23;
reg  [MAX_SUM_WDTH_L-1:0]        I4ddbc3daa65b111cb0d45e13d62cc292;
reg  [MAX_SUM_WDTH_L-1:0]        Id363d158feb8fec19b5f3d73d84f0068;
reg  [MAX_SUM_WDTH_L-1:0]        I8ec9b7a6e65e727abbed336ce240a4cf;
reg  [MAX_SUM_WDTH_L-1:0]        I128fa1e99b7eb9b6905c2cfd26b95ab4;
reg  [MAX_SUM_WDTH_L-1:0]        I93d459b6da42a205c91c48622f0c5032;
reg  [MAX_SUM_WDTH_L-1:0]        I1243cc8d5dddf7dd65b40c0b3b958b9e;
reg  [MAX_SUM_WDTH_L-1:0]        I238df7e09d42bc93a972da349a00f511;
reg  [MAX_SUM_WDTH_L-1:0]        Ic658b2afdc7331653fc84d6372d47418;
reg  [MAX_SUM_WDTH_L-1:0]        If39be111eb101c9c983fe0baa9a1cb18;
reg  [MAX_SUM_WDTH_L-1:0]        I9d19d5b7d8b256c1707de97a4549c458;
reg  [MAX_SUM_WDTH_L-1:0]        I6c2fffe204091f7f64aea16b0ac98769;
reg  [MAX_SUM_WDTH_L-1:0]        Ic4ba4d2e5c12d9f1dd233d64929f1072;
reg  [MAX_SUM_WDTH_L-1:0]        Ia9dec5831998d472d11429e5a7e60ed8;
reg  [MAX_SUM_WDTH_L-1:0]        Ieaaf52c1e663f260292bc1529718d681;
reg  [MAX_SUM_WDTH_L-1:0]        I37061896a09588a73445deed73d3746c;
reg  [MAX_SUM_WDTH_L-1:0]        I02f25b80945b6f58193fb37add3da2d8;
reg  [MAX_SUM_WDTH_L-1:0]        I19045602bb77f12666ebd44f813db2c5;
reg  [MAX_SUM_WDTH_L-1:0]        I4abdc8d5318d2922696a8aaee46ffa59;
reg  [MAX_SUM_WDTH_L-1:0]        Ie139f2048f346d82623c8fc6d40c9acc;
reg  [MAX_SUM_WDTH_L-1:0]        I8d99c96e203fafc81d13ce5aee925d75;
reg  [MAX_SUM_WDTH_L-1:0]        I37b0bdeb3cc54d6a97720c4912c67832;
reg  [MAX_SUM_WDTH_L-1:0]        I08257e9e6c74c60448e22fb9855f0825;
reg  [MAX_SUM_WDTH_L-1:0]        I32188cca2fc715698fc05b0fc6506434;
reg  [MAX_SUM_WDTH_L-1:0]        I88f1cbab9b8fa3802345f745d024931c;
reg  [MAX_SUM_WDTH_L-1:0]        Idf548c0e78bd221bf9f612f27002fae0;
reg  [MAX_SUM_WDTH_L-1:0]        Iedfd2e04f5740d283388639dde3ecdb5;
reg  [MAX_SUM_WDTH_L-1:0]        I7088c83eacff6f1dfb134f79d469c8f1;
reg  [MAX_SUM_WDTH_L-1:0]        I6f8431671331f4ca7ea19656e0677cd4;
reg  [MAX_SUM_WDTH_L-1:0]        I1e31259e267e04920cbbd16bd7aa18bc;
reg  [MAX_SUM_WDTH_L-1:0]        If54d9f8088e67e44cfa3026f5a520fd7;
reg  [MAX_SUM_WDTH_L-1:0]        I6fd2c0746407b23aec5dff1e083f5fca;
reg  [MAX_SUM_WDTH_L-1:0]        Ib2147a19b44d361da628a628fbfaa988;
reg  [MAX_SUM_WDTH_L-1:0]        Ie804d1f4b241a2de3e9d9c7c876d914a;
reg  [MAX_SUM_WDTH_L-1:0]        I6cd1e6db57e06d8f5e60a31f48ae4809;
reg  [MAX_SUM_WDTH_L-1:0]        I3e0e8832d5338423284ac4b2a0c5f3f5;
reg  [MAX_SUM_WDTH_L-1:0]        I6ac006d79e95e222cdc66754b67a08ed;
reg  [MAX_SUM_WDTH_L-1:0]        I29087dda1a527842aeb3d35d66c853cb;
reg  [MAX_SUM_WDTH_L-1:0]        Ia67e5920bbac700dfee52cd96b15963e;
reg  [MAX_SUM_WDTH_L-1:0]        I1f6ecd894d90547f661e7a3888d048bb;
reg  [MAX_SUM_WDTH_L-1:0]        I3112e793c6e79e1f5da2776e69a34e3c;
reg  [MAX_SUM_WDTH_L-1:0]        I79152f32b45ed5b4a5302f6460707b01;
reg  [MAX_SUM_WDTH_L-1:0]        I3d16e7d6b190639b88a217f19ac63233;
reg  [MAX_SUM_WDTH_L-1:0]        Ia1be780c686163cea54b62d6ede72dc6;
reg  [MAX_SUM_WDTH_L-1:0]        Ic398c31a2a6ca89d0236534589a5919b;
reg  [MAX_SUM_WDTH_L-1:0]        Ie91c3202bc957b350d1915000564392f;
reg  [MAX_SUM_WDTH_L-1:0]        I687957f5300b0d4f50d6893cc556bf25;
reg  [MAX_SUM_WDTH_L-1:0]        I7816b368e8e8b8dd69383b2c9327120d;
reg  [MAX_SUM_WDTH_L-1:0]        I5f021f4a664205afbe0761af4c8914f1;
reg  [MAX_SUM_WDTH_L-1:0]        I69728004b59b5206a03a8e2087834f7d;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbe1d623f8f5f3aa7fc70197acc6df5e;
reg  [MAX_SUM_WDTH_L-1:0]        I4cb9f74288811592fd97fdff52bd6fe7;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb471dbccd39d41e951e98348812e343;
reg  [MAX_SUM_WDTH_L-1:0]        I7f37d68f8ddcf8b4d5e99fb51eada873;
reg  [MAX_SUM_WDTH_L-1:0]        I72ded7153883418a712ef967439d2159;
reg  [MAX_SUM_WDTH_L-1:0]        Ie071e08299bff6bbdbe1f84703aaec08;
reg  [MAX_SUM_WDTH_L-1:0]        I1b79aa38a39ccfc839260af89aa78e7a;
reg  [MAX_SUM_WDTH_L-1:0]        I7384296e4190d83fb9d9a92cf965125b;
reg  [MAX_SUM_WDTH_L-1:0]        Ie03034ce6233ca24effe53a2c0c8f6f3;
reg  [MAX_SUM_WDTH_L-1:0]        Ic298f77f42fc1d41cce684790036ecfe;
reg  [MAX_SUM_WDTH_L-1:0]        I805269f95afbeb6b93182f68868d08eb;
reg  [MAX_SUM_WDTH_L-1:0]        I881328804c45b06767af51e11182b27b;
reg  [MAX_SUM_WDTH_L-1:0]        I958993626e6e44e12f7c1e8026914680;
reg  [MAX_SUM_WDTH_L-1:0]        If31528d1fc3a083ebc364e75cdd9c71f;
reg  [MAX_SUM_WDTH_L-1:0]        I4703b8d5a9033027889bfa8685e09e4f;
reg  [MAX_SUM_WDTH_L-1:0]        I22d8e84d2db4b07111b7fdc6eef34cc8;
reg  [MAX_SUM_WDTH_L-1:0]        I8b7c6df3b5ea575caab7820c95974608;
reg  [MAX_SUM_WDTH_L-1:0]        Ia8aa76bccf7eb310a9356e8b7ea1609d;
reg  [MAX_SUM_WDTH_L-1:0]        If9de547bf469b8424f1625e990f72b04;
reg  [MAX_SUM_WDTH_L-1:0]        I27d51b2015ea9af9bc345adabdb07b6f;
reg  [MAX_SUM_WDTH_L-1:0]        I93dddce2a0dc01ecb3039fac5cf04011;
reg  [MAX_SUM_WDTH_L-1:0]        I746da2c1d5a620eb7e749f72f0f04a06;
reg  [MAX_SUM_WDTH_L-1:0]        I1e15f8d6fdb4ac732768d0cf73af829e;
reg  [MAX_SUM_WDTH_L-1:0]        Ib719e667d7ba857f4f7432a245f4a30f;
reg  [MAX_SUM_WDTH_L-1:0]        I4c6eec4a0c46e4f5d7c9734df48a16bb;
reg  [MAX_SUM_WDTH_L-1:0]        I95623ec1fd5516040a9492aae0fc2b70;
reg  [MAX_SUM_WDTH_L-1:0]        I69017b49c11de463fe6d881e5c96a1aa;
reg  [MAX_SUM_WDTH_L-1:0]        I4fb9ed32471aa614ce6923f6a2279b36;
reg  [MAX_SUM_WDTH_L-1:0]        I2f0bc217c8a39d71adc1fc45c10b81c3;
reg  [MAX_SUM_WDTH_L-1:0]        I0f1c6bb577ea2b8b2ab636e64378544b;
reg  [MAX_SUM_WDTH_L-1:0]        I7a248af9d606c566e03977e985c280e0;
reg  [MAX_SUM_WDTH_L-1:0]        I0bf9d47bff47277de1e72518e8d88362;
reg  [MAX_SUM_WDTH_L-1:0]        I24b6f4f68f291dc50caf03dc902282cf;
reg  [MAX_SUM_WDTH_L-1:0]        I79335b28eea15735f760b7a8b803e93a;
reg  [MAX_SUM_WDTH_L-1:0]        I0b14b34b06cfa90539c2abca5639abec;
reg  [MAX_SUM_WDTH_L-1:0]        I26878777354945712f834740b17dabcb;
reg  [MAX_SUM_WDTH_L-1:0]        I6cc5daed4de5950c02c0a57b993e22fc;
reg  [MAX_SUM_WDTH_L-1:0]        I52c382d5b0c4829127c011fae402ce04;
reg  [MAX_SUM_WDTH_L-1:0]        I46ea9871e867034daa2d0501038f15e0;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb8a202599550e87831647a93a14181a;
reg  [MAX_SUM_WDTH_L-1:0]        Ibb79f2ce0b6028ebb638fc6661444cf1;
reg  [MAX_SUM_WDTH_L-1:0]        I0d0c07d65eda2eee01df9c330c0d6f4a;
reg  [MAX_SUM_WDTH_L-1:0]        Ie6940736944bac9be609b8d58b2cb13c;
reg  [MAX_SUM_WDTH_L-1:0]        I472a71363435cb3ec054e00f9123ae64;
reg  [MAX_SUM_WDTH_L-1:0]        I553223e9166dcbddd1a51d0f92d68f28;
reg  [MAX_SUM_WDTH_L-1:0]        I495309d795905a53b0a3d3daa4f1f9d0;
reg  [MAX_SUM_WDTH_L-1:0]        I21d358fd7673c4392f4e4b3d3a858b2c;
reg  [MAX_SUM_WDTH_L-1:0]        Ia1a60175112362f015c5531f7c48b90b;
reg  [MAX_SUM_WDTH_L-1:0]        I5644ece811bddcec04c9e3559c86109d;
reg  [MAX_SUM_WDTH_L-1:0]        I37d2f9d3f05cb90e2d45bd578299885c;
reg  [MAX_SUM_WDTH_L-1:0]        Ie7d10f3c0f8b0add66d2cdd4435ccc88;
reg  [MAX_SUM_WDTH_L-1:0]        I3c37396a1cef2f9e42b8ccc126db6eda;
reg  [MAX_SUM_WDTH_L-1:0]        I2f82390734079b8d289d48a6682cc624;
reg  [MAX_SUM_WDTH_L-1:0]        I9061728c3163ae684e8c5aec3e807868;
reg  [MAX_SUM_WDTH_L-1:0]        I672d7ecc28a788c2602aff76187aa568;
reg  [MAX_SUM_WDTH_L-1:0]        I660b2fe99cd0bcaac34e9540118b54bc;
reg  [MAX_SUM_WDTH_L-1:0]        I6aa263fc2a061d2c4059b08309f860f4;
reg  [MAX_SUM_WDTH_L-1:0]        If3aef2d755013d195fd44f734365d7dc;
reg  [MAX_SUM_WDTH_L-1:0]        I3ad2e0bbff17683824f575deff82c6bc;
reg  [MAX_SUM_WDTH_L-1:0]        I5087dc4b32d29bfd7bad49026fa58a5d;
reg  [MAX_SUM_WDTH_L-1:0]        I8a7d893f3ef6d6a93ba552320d901599;
reg  [MAX_SUM_WDTH_L-1:0]        Ic057537712e09fa794918e5cde87e084;
reg  [MAX_SUM_WDTH_L-1:0]        I0cbab5173052c450504e3a7d15ffda52;
reg  [MAX_SUM_WDTH_L-1:0]        I81ee40feb7abd0fec3faee653f778f5f;
reg  [MAX_SUM_WDTH_L-1:0]        Ia344347a85d4e6afafa2ee3487e65def;
reg  [MAX_SUM_WDTH_L-1:0]        I038fce1597157a3d95bd9579cc2dcbc6;
reg  [MAX_SUM_WDTH_L-1:0]        I546585b819c289d855cd098818792e90;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc3a6609765818327e79519f3e348494;
reg  [MAX_SUM_WDTH_L-1:0]        Id1c71a2a34f9e6239559d28fe2780907;
reg  [MAX_SUM_WDTH_L-1:0]        I1cd6cf5f8119d5e6b4ca40694399b1c2;
reg  [MAX_SUM_WDTH_L-1:0]        I15e2a1b4356785d73e2ab5d51f1f5ec0;
reg  [MAX_SUM_WDTH_L-1:0]        I803aeb29e66384bfc62744a841bcc83e;
reg  [MAX_SUM_WDTH_L-1:0]        Ib6e220dd4f54410239dd0c791d84a700;
reg  [MAX_SUM_WDTH_L-1:0]        I8a009007fec23f4d492b0da1b6b404fa;
reg  [MAX_SUM_WDTH_L-1:0]        I5f89adcb1ba235a74639eca119fb2655;
reg  [MAX_SUM_WDTH_L-1:0]        I8fd2b001ff154e4760ead2df355c80da;
reg  [MAX_SUM_WDTH_L-1:0]        I581569cc2e63bc68a8466b07ca471b25;
reg  [MAX_SUM_WDTH_L-1:0]        Ia9cfdea21a65b0270de42cef7ebbf822;
reg  [MAX_SUM_WDTH_L-1:0]        Id66a233d2e312aff939549dfa96a8cf0;
reg  [MAX_SUM_WDTH_L-1:0]        Ie479c12c25a1964c3804936d45725bdc;
reg  [MAX_SUM_WDTH_L-1:0]        Ie30d8770ab7e6643fcb67463f6999125;
reg  [MAX_SUM_WDTH_L-1:0]        I4a17ff532c9341e80f7ed0626f728054;
reg  [MAX_SUM_WDTH_L-1:0]        I597bc1ec224007a78c25f7eea24c2c3e;
reg  [MAX_SUM_WDTH_L-1:0]        If198ec15fcf66e97e69f88f718979c2b;
reg  [MAX_SUM_WDTH_L-1:0]        I6aa13ef29cf7e86ec83affca4fa11e42;
reg  [MAX_SUM_WDTH_L-1:0]        Ide136b08f4b6211bca8cccf494a0baa5;
reg  [MAX_SUM_WDTH_L-1:0]        Ieeab247764c23256749776b0a164314d;
reg  [MAX_SUM_WDTH_L-1:0]        I210e9ff7f4588185bd712915954543ce;
reg  [MAX_SUM_WDTH_L-1:0]        I59186d5219833d6dd2e813a2910a61f5;
reg  [MAX_SUM_WDTH_L-1:0]        I0c8b2bb61a9c3a67ac7e03e40be2b98e;
reg  [MAX_SUM_WDTH_L-1:0]        Ide24c1f9033e7057262da1bc4762b840;
reg  [MAX_SUM_WDTH_L-1:0]        I4677558b9faf190e7960cfa9b8ee00fd;
reg  [MAX_SUM_WDTH_L-1:0]        Ie38ab94215851e531d2100b6602d5fa5;
reg  [MAX_SUM_WDTH_L-1:0]        I3f5119e8fac99376aa38e4765b8b0f99;
reg  [MAX_SUM_WDTH_L-1:0]        Ie8040301d224f78c1fd18bfe9e29e5ba;
reg  [MAX_SUM_WDTH_L-1:0]        Ied989966cebf0d730633606c5182a249;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8818bc4ca106ae38cacd5c20083aa08;
reg  [MAX_SUM_WDTH_L-1:0]        Ibf08556fc39044222321912e84a4436b;
reg  [MAX_SUM_WDTH_L-1:0]        I985e2740ac0f656da8f9dd973bca99e6;
reg  [MAX_SUM_WDTH_L-1:0]        I73012d2d9f6f237bc50bbffc199e012b;
reg  [MAX_SUM_WDTH_L-1:0]        Iefd0d59e58623b14437b17297fdbf4ff;
reg  [MAX_SUM_WDTH_L-1:0]        I68d2443e98f2fd3fa3baf96f98e1f4bc;
reg  [MAX_SUM_WDTH_L-1:0]        Ia2d1b6833cd8ed02f05281e508e4d716;
reg  [MAX_SUM_WDTH_L-1:0]        I512e2251bef73108eb0f3e01e79ca3fb;
reg  [MAX_SUM_WDTH_L-1:0]        I9bf64811d14ca8b4c633342ad22669a3;
reg  [MAX_SUM_WDTH_L-1:0]        I45a910acd40d5b9417bdfdc50cddf241;
reg  [MAX_SUM_WDTH_L-1:0]        Ibbcf5c5f4528b03508b506c43e4511c4;
reg  [MAX_SUM_WDTH_L-1:0]        I2b8b54048e164ef2f1c072517fdfe400;
reg  [MAX_SUM_WDTH_L-1:0]        Ia48d8883fe4f685477da6b4b05ecd387;
reg  [MAX_SUM_WDTH_L-1:0]        I276395da1f3f1ae246b082408be2cb80;
reg  [MAX_SUM_WDTH_L-1:0]        I4d0e2e01d9abf9ce839fe650abfaaddd;
reg  [MAX_SUM_WDTH_L-1:0]        I7e4e7909094f762c54137cbee99255e5;
reg  [MAX_SUM_WDTH_L-1:0]        I761255e100d161b25645ca3a5187e82a;
reg  [MAX_SUM_WDTH_L-1:0]        Icc2ce1fa3cde69256378ec3f4a07b0fc;
reg  [MAX_SUM_WDTH_L-1:0]        Idd99afa80ca23644675d3edd60e74fe4;
reg  [MAX_SUM_WDTH_L-1:0]        I486bcb4fb0af80c98c2ea21ac64f7a90;
reg  [MAX_SUM_WDTH_L-1:0]        I759cca2c0003fc2c2af7709c5ebc59f7;
reg  [MAX_SUM_WDTH_L-1:0]        I1d5ce9f132cd1f46e96b511c77234e21;
reg  [MAX_SUM_WDTH_L-1:0]        I032e26ea05e88c6d325a810b67e82306;
reg  [MAX_SUM_WDTH_L-1:0]        I0f72df5225a1fec2f276fd3c9138e8c3;
reg  [MAX_SUM_WDTH_L-1:0]        I0d18cf087b2335f1b9e1a621acd5379f;
reg  [MAX_SUM_WDTH_L-1:0]        I7684fc23c57105e856050a45640f2bfd;
reg  [MAX_SUM_WDTH_L-1:0]        If778767ab80e59e940deeaa8a0dac99a;
reg  [MAX_SUM_WDTH_L-1:0]        Idaf86833beb8c334f99291db9302ed29;
reg  [MAX_SUM_WDTH_L-1:0]        I6610e8d41cea10498d95850440ce388b;
reg  [MAX_SUM_WDTH_L-1:0]        Ibc653e701eb995e828c8180efaa122c9;
reg  [MAX_SUM_WDTH_L-1:0]        I21d36c49c9c766139b4b01df7c00a8f3;
reg  [MAX_SUM_WDTH_L-1:0]        I0e4ffded936d7ccfc32b410aec617df8;
reg  [MAX_SUM_WDTH_L-1:0]        I1a5745021323efb5327d0b893962e852;
reg  [MAX_SUM_WDTH_L-1:0]        I65547afdcd7fedb7b44bd51358eec4d2;
reg  [MAX_SUM_WDTH_L-1:0]        Iada3eb71e94ff6a6f4e5c702e83036ed;
reg  [MAX_SUM_WDTH_L-1:0]        I077404a911da16d707a326f18717dc7a;
reg  [MAX_SUM_WDTH_L-1:0]        I6da1e92759c96aab8b9207a9acb244ab;
reg  [MAX_SUM_WDTH_L-1:0]        If7110182720ffa279b1cec1305cf9889;
reg  [MAX_SUM_WDTH_L-1:0]        If0e20ea1696ff84329b9928d7f9e3381;
reg  [MAX_SUM_WDTH_L-1:0]        I4e69ae6e73a856d4e26203fb9acf3565;
reg  [MAX_SUM_WDTH_L-1:0]        I64c939aa568669b4567c21be09ad0e94;
reg  [MAX_SUM_WDTH_L-1:0]        Ia88eb16f68265e322509d541eb457993;
reg  [MAX_SUM_WDTH_L-1:0]        I916f75e5a3858a420ab5cd4c43b13921;
reg  [MAX_SUM_WDTH_L-1:0]        Id076f99460a8f73a9fd43467216e8f8e;
reg  [MAX_SUM_WDTH_L-1:0]        Ib4d7aeb8544fbdc36575a55b9f67f2dc;
reg  [MAX_SUM_WDTH_L-1:0]        If65d2514892fb7ee64fa4dc37fc0fed3;
reg  [MAX_SUM_WDTH_L-1:0]        Ibef07e48768252e9b41baf067bb1ff5d;
reg  [MAX_SUM_WDTH_L-1:0]        Ib8fb61fa9cb8e92bc57c53a567891895;
reg  [MAX_SUM_WDTH_L-1:0]        Id8f5f32cd0757b4d6861d17fcbd6e8d0;
reg  [MAX_SUM_WDTH_L-1:0]        I8be241f29e7eb258e9b3501430820b0d;
reg  [MAX_SUM_WDTH_L-1:0]        Ica8a188ea43e2f28e70b8ea4e2431dc3;
reg  [MAX_SUM_WDTH_L-1:0]        I83ceb726e57d52698b57dc39ce585897;
reg  [MAX_SUM_WDTH_L-1:0]        Ic88e7e05d83ff800b4a941ae4b424557;
reg  [MAX_SUM_WDTH_L-1:0]        I7de81aaac1e5776dfb60eed2d12d4f6d;
reg  [MAX_SUM_WDTH_L-1:0]        I37058036bd9f4331387ee4a9348541e2;
reg  [MAX_SUM_WDTH_L-1:0]        I570f85838c418d8501c8ccdc38a53f00;
reg  [MAX_SUM_WDTH_L-1:0]        I4aa6f0c0f5163b944f11328888af73e0;
reg  [MAX_SUM_WDTH_L-1:0]        Ic7fc1f38ad4e9b2cb472ae75bc3c100c;
reg  [MAX_SUM_WDTH_L-1:0]        Ibace8d2fba25834c83b1e57195c81086;
reg  [MAX_SUM_WDTH_L-1:0]        Iefc1488e3eb60b99ae08d904a15c5242;



assign I97afe24956b7f87cd431f048202bab67 =  ~I5deafec6e5f32da1bcf8f7018cf794d8+ 1'b1 ;
assign I117235e3ac8e68e4c1ab34db1612aba0 =  ~I35b3fb2670f3a60d165c1fd10f02c00c+ 1'b1 ;
assign Ifd700cc9d18f99b63f1947f3ae631976 =  ~I68925439e233444a4da44871f31de94a+ 1'b1 ;
assign Ifffbe3d1007fb07a20d3b37902b3ec95 =  ~I3108702b5ca506422c1ba6174619f193+ 1'b1 ;
assign If5443777169422ea6e1e3f709b970e05 =  ~Icc8e8f6446ac64350a05f5e1e0541bb9+ 1'b1 ;
assign Ifaf9fc93e4609d818aa46751754c17f1 =  ~Iadebaf3f6cca1ba78feab50ce70c8aef+ 1'b1 ;
assign I419caf964986c655df84d043badc37c9 =  ~I8681cf376dbeceab29279a7637249e7d+ 1'b1 ;
assign I3095214ac0e6c1323e75ee4ec85e6821 =  ~Ie850a07565bed90389bb125ddcd39658+ 1'b1 ;
assign Ided9739bf63937933250a6d0c37535f9 =  ~I97b77743c2311ec629ea24c933b60053+ 1'b1 ;
assign Id0f139b9f3848b45554ac8429230eea2 =  ~I07a0a8d41ed8176e92380f2c89c2afdd+ 1'b1 ;
assign Id9feed58cf9565255abfd0bf7e3ec068 =  ~I021842328f948a94159b32903c8bcb68+ 1'b1 ;
assign I30a3be3b5f6ad1880a917eb35659a1bf =  ~Icaf3bd685005a05c8fb334266ea4e4b9+ 1'b1 ;
assign Ie8148d9aa962a733eb65877b902a187d =  ~I92d9e1d7dcf45a4d738c546e959687c3+ 1'b1 ;
assign I69e98cf3e679183aef6005bb582b18dc =  ~I39ca3a8ca714a9726114326ae6bfab0a+ 1'b1 ;
assign I7f42a504fc61c9548acebdd8b1858eaa =  ~Ie9ae20ed5b2a0cad2c37c5bb2ea05ff4+ 1'b1 ;
assign I08b1b4639b5a9ca509b943b977f6d4bb =  ~I8f131eb6138c23fdcb35195703131e64+ 1'b1 ;
assign I8d7296627d886566783e79c01b9fa423 =  ~Iff77e08da4bcbb85b95fa277b69653a9+ 1'b1 ;
assign I4fc4c97229a8b1f631a3b505941159e4 =  ~I703e0a4879a39b3b8b0a49de86ca4ff4+ 1'b1 ;
assign Ib9b16bf51891c328dba2699eb9bcef95 =  ~I3da217f6f2d0f515bb9036673d753a88+ 1'b1 ;
assign I6c30501ec81fce286817788d614a7824 =  ~Ifcc06d5a010e01a781ae8a9e9e2b31a0+ 1'b1 ;
assign Ia4d4f37baec48121a88808075dd655ef =  ~I42fd611fec087113ba6e35f281bced9c+ 1'b1 ;
assign I385495ea2bf6442a95ab7561456254ac =  ~I5bb626e7347bb9ae4219cc72244b38f8+ 1'b1 ;
assign I5128e03d383c226befa6f7422f3a6f04 =  ~I47e2dac0068652338f94ddffd2dbe88a+ 1'b1 ;
assign Ib208908bab4c20713cd17e20139c8db3 =  ~I59a3f06de2984078a4d4c430a2980fe3+ 1'b1 ;
assign Id939992b99a11c09f4688c10ca1a34d1 =  ~I857b7fd58279b1063a06a4f33b880ba6+ 1'b1 ;
assign I823453ccb90d5b2b2d9dfc6e8358224d =  ~I3901bbda029cd0a41640001c1efd400f+ 1'b1 ;
assign I279c5c00b92eb1b872b5afa168b0306e =  ~Ifceeccf10f1d85a32f70c04654a1a1b4+ 1'b1 ;
assign I66f25b1c3c0eb226295179adcca2c3d2 =  ~I2d810c1d1304658edff74921e8d0f388+ 1'b1 ;
assign I3068627e91b667d14cd3e55a9371931a =  ~I575b0201be445388607ab83465eab8d6+ 1'b1 ;
assign I44c4e0a2d8a7289f8660b81a9ecfa19b =  ~I7928c5ce0f821df1cb6271d15e19fa22+ 1'b1 ;
assign Ibe868e258dc87f0dd1460ba6b8354671 =  ~I12695a21c942d02a432cf6382d7d7452+ 1'b1 ;
assign Idc3083c3021200345e3edd35a9d4725a =  ~I00d03f0f71b008dad8035bbf251f41bf+ 1'b1 ;
assign I320d4f19a5b18c23ff407508d47caa77 =  ~I41afedcbc0f492e3243436cbefdaf609+ 1'b1 ;
assign I16becf3c92615d98d5ec51ee9641cc0a =  ~I638c4c2708e437a050ed7cbbac516a59+ 1'b1 ;
assign Ifbfacc3b3a0128119943bcbf80176612 =  ~I6877d3306b1f08c236b5d1b59f0de259+ 1'b1 ;
assign I6b4f670c9e8e25984e8891f2440322ab =  ~Ib3e66aa460f39d32110ea6f115785b3d+ 1'b1 ;
assign I19bf0990a30c72421f231772b8627e8e =  ~I5e603e8392a5322951b3225b65b19446+ 1'b1 ;
assign I3ec3eb096ebe3ee8a47e1cba6487b997 =  ~If5da7fa1a615e1122445460e33487772+ 1'b1 ;
assign I7379ef16405c461ac44b66c4315df831 =  ~Ic4153dafafaf7d047478c5d81109437f+ 1'b1 ;
assign I79db45b23d21d533a1f9a6e8f94d403d =  ~I7b5476007f04e81afc0125e6a8930303+ 1'b1 ;
assign I0979534730cc2b53547d413dbb6b75f4 =  ~I3521a18022925249caddb8e37d2c1262+ 1'b1 ;
assign I5aa2f9c0667d1a6e871efbd4d2bad3a8 =  ~Ifd0f52d4f814e2bb4c3bd34c1e09bda7+ 1'b1 ;
assign Iadb28dc990ccf2dd3099544de16b8f16 =  ~I8945f6d420c8b373225451defcd2c805+ 1'b1 ;
assign I1f71aebf698788d6ada66891e9ea756f =  ~Ieec6cb6518cc0d9300de0c4f2d32487d+ 1'b1 ;
assign Ib234e9cf7e7616a1ebc6ab99df2a7ccb =  ~Ic62eb7e90d703ef994e68587345a4293+ 1'b1 ;
assign I297d1edcc583ea4d69da780150f0620c =  ~Id3efd8419da986aa89b8ad8e75848cfa+ 1'b1 ;
assign Ib0a717cbb4fe38a3fc85520ca0826fd9 =  ~I40803f10b7c4dc9ae4969739349b0265+ 1'b1 ;
assign I037ecd5945b1f1280b4469d73fe1c7ff =  ~I7d961743fdeaf1e72e4b25c12a1d4c46+ 1'b1 ;
assign I367ff6b11b884e02a3065fc7fe811e15 =  ~Ifea156f33eb61fece272efe379327f6e+ 1'b1 ;
assign I6fab19692b512166fe9c74b5e987788d =  ~Ifc99169b3399f3d14121c1a9bce3fc21+ 1'b1 ;
assign I04dd73af505f618ccdb209b3cf97ceec =  ~I6536144383cbda6f3b3c564391866906+ 1'b1 ;
assign If8c559905d4120488d431719c4e8ce24 =  ~Ic21bf9a8a4cd85ec123d7fe142ed49c0+ 1'b1 ;
assign I20ed4f6f14e20ce3f0e106d1b7782fcd =  ~I1f31fe6a0ca8510bcadbc2069403150b+ 1'b1 ;
assign Ib10626ffa126188c5bf1fc8399107b26 =  ~I0e40933d00f4a7d9b53b2764aa0da700+ 1'b1 ;
assign I29007c52357ac7afbda39d72a5bb60af =  ~Ic41a6e00bc84bfc1b8194d15bb899c93+ 1'b1 ;
assign I66d367c046611f145e607a90911cf499 =  ~I2832571f2b0a7fbb41d2e8ca7f64e003+ 1'b1 ;
assign I9c4c2556f6170a8df61d909855a846ed =  ~I9593c853e41952e408a809cb24efa4fd+ 1'b1 ;
assign I6fadc3e8d995bb4317bf7b4377c3c2c5 =  ~I6edffbf4136e193dca0fcec3a74e8e9c+ 1'b1 ;
assign I99b20e911c189e0616f02376ab736e91 =  ~Ibaed50cc2e36ae58945887d11a6ec9e4+ 1'b1 ;
assign I5793c12f5dbdd8245dbb202d550ca960 =  ~Ie4570cac44f59e6ff46f73a703026479+ 1'b1 ;
assign Id0660e9637cad1ce1a73d37188060154 =  ~Ibaa136d37936687e9dbe4222749d19c3+ 1'b1 ;
assign If5a7af7ca023e1393526e888f4220a44 =  ~If85de3225f45478827b43b89089cd29e+ 1'b1 ;
assign Id043eb50634e803e53adc1168379a5d0 =  ~I0344b86a6e9c036e103a9c1f3651175f+ 1'b1 ;
assign I1f866dd0b129267550aea1a267d9c91e =  ~I5463d13575e0b9fb8a0f6cc8b35d0ce9+ 1'b1 ;
assign I8c4da05c08210fe33139c3d3e5d75d58 =  ~I8a3c63ef122001a29e5abe93c4e1a48f+ 1'b1 ;
assign Ib41f7b823681fdd084b6d8436a407aa8 =  ~I6a79108484fcb192f6d93bfb98e271c4+ 1'b1 ;
assign Ic5b50a785b7acac7e3be4095aa92e50a =  ~I9001e95b71457a2bd09a9846af370b16+ 1'b1 ;
assign I3ffbe03796b66d00d47fd918be60ab89 =  ~I51620de618db6327358a5cac97e1e97f+ 1'b1 ;
assign Ifc92a916da938ef6164db250be635f88 =  ~Ib9c58818059af5c5a03e77a5dcef4654+ 1'b1 ;
assign I8ccd42508ce7d5bd897c2cf0c54caeb3 =  ~I8081c71aa01a8d575bfea6ea7f2f595f+ 1'b1 ;
assign I4920e7e82749cc036b58a7cd0a03e327 =  ~Iad999607ad8d7da0f3b341f83ea030a6+ 1'b1 ;
assign Ie1040b2aa91f272e4449c4b5f9f8f575 =  ~Ie7291c914d2cb66f547b0a7717f71311+ 1'b1 ;
assign I65968fb0f63d52ad96cd8fa270126a1b =  ~Ic01018a5f1bc392bbd267016f6612a83+ 1'b1 ;
assign I839ac8ee59f51d4c3de92ba5cb26e788 =  ~Ib11dff839e7e532657b32f29fd9b1651+ 1'b1 ;
assign I33cd95f1919318a0f3df5df7310d64c6 =  ~I251d7ea16dd5407d22a6846ddcfe12d8+ 1'b1 ;
assign I4933e8d16fba26cd797b25a9ac2a2de8 =  ~I773797f81f73b9b6e844441142a1bb48+ 1'b1 ;
assign I218f7578eb748e31d0002052f30c5842 =  ~I853ecadf30fc10a13dd1ffb1f2dfb5d6+ 1'b1 ;
assign I2a808d1c42ad758ae3baaaee8129dfb2 =  ~Ibb8b3c91e1d3b890cfe58f32f8ec3ae3+ 1'b1 ;
assign I4e851fd3c114af87f5e8c68c02594e3a =  ~I3485d69de942d64e56925da522175b51+ 1'b1 ;
assign I0da40f88adc46e90f616acdcdb8e0e2c =  ~Iae42f12bc0475c8b58341d80027a57cb+ 1'b1 ;
assign I0dee7767e472a5fd71250ae6c57cc8b5 =  ~I22fe2af25463f87ee7315a9aac32854e+ 1'b1 ;
assign I9f40be7552b3dd625e5bce0befc5a548 =  ~Idf44ad78c338c39699721ce511691dfd+ 1'b1 ;
assign I8fdf98ffd757c8845ed6ffa4ddd1a16b =  ~I984a657f9265d41318c0290e249e9712+ 1'b1 ;
assign I8103b777314a4fa471e0898fde9cde08 =  ~I915fccfb1d1ada9aa7c8e24c2eebd04c+ 1'b1 ;
assign If6c3ee8e0d7dea58043d5be0f4630873 =  ~I2bdf58ecd0974720631be830efb48dc8+ 1'b1 ;
assign I711a5171f591f472cdbfc9a0f5e1aa17 =  ~Ibaedf6246fa43acc8accb5a24d49cc2f+ 1'b1 ;
assign Ic30bc38184dfbbd694af52640692709d =  ~I904d13524dcdf55478a5266d50e53ff7+ 1'b1 ;
assign I422f6fd1d273a3834d04b04ab8e2812d =  ~I22d8e5d57c1bc082169437a654d22bba+ 1'b1 ;
assign Ia0fdc60b90ad18b6585ec1ad4e89e80b =  ~I719cdaa2a2e61a0df7f1fd5efe517426+ 1'b1 ;
assign I7809fe7a30d041a7e569ffe890242df8 =  ~I8e92a61eb73c41680652936cfcc614ff+ 1'b1 ;
assign I672b14ec1b3c4797545f266727505a85 =  ~I7ad5af8319f6da469858300f0777b580+ 1'b1 ;
assign If9620d20ebaae6245a2c386d9bf5fdb1 =  ~I32be72eaf04e79120a57ea94296a4e56+ 1'b1 ;
assign Ic74e22bffd88f32eefe499cde0fafa8a =  ~Ie756f6a87d85adb40479ce7cf3545556+ 1'b1 ;
assign I76d38ce67387bd76ab45c9cba7d18b31 =  ~I8794c6ce0a3f2e6697372e2c911ba420+ 1'b1 ;
assign I44413c6f6f6493f8a86abf6eb32604f6 =  ~Ic82b1a29b5e63bcc3686a0d4bf1f5c24+ 1'b1 ;
assign I67f632fca617fe06565ddcaaee8fa8b8 =  ~I253ef976058080beab79646af18e2d5b+ 1'b1 ;
assign I3fd38a71ce6aa3db1d7a5a9f8a991e12 =  ~I930dd54c36540d75dc870eef89960163+ 1'b1 ;
assign I63e5718bf7d8771ef90b91be73d73264 =  ~Iaf7554cd4e8b5ea6155ec61a8d589b86+ 1'b1 ;
assign Ie385e1aeb2b0dcf6d2454be3d7708b27 =  ~I50907c7d1efa0038d81efed82b192891+ 1'b1 ;
assign Ib2d1b7e105b25b492b45da72536d7578 =  ~If3e9486d2960d164d94641d4f1917416+ 1'b1 ;
assign I588abf5ef4c583f0fec422736a0ce6a0 =  ~I2bec61db45dd79b98d6ebff6c5a4899e+ 1'b1 ;
assign I58bb95c56c7be17c263a2161210d7d8d =  ~I7f31647f3ea6ce7bbd211c25cf4828fb+ 1'b1 ;
assign Ifaf0e1f21b3bd7393c475b5126540a72 =  ~Ice65387e606faf9c7b884475b489abba+ 1'b1 ;
assign I7027db9e0450724a6d417d708f1043f2 =  ~I63f914927dcf49552e9f3fe0180a30e8+ 1'b1 ;
assign Iebcb7206d8860b5094459c5d10b4efed =  ~I742ff5725e3a18acd03454cf9f313f4b+ 1'b1 ;
assign I6bbf2b47a7dc50e66a3d8d258d6e31fb =  ~I84e4b3bc63ec0b0bff7f98f433c1fd67+ 1'b1 ;
assign I8459abaa907f5afcd11884b1ec8c06c5 =  ~I78c6a1428a1f211c5e89b8c76b3dc033+ 1'b1 ;
assign Ia16ae2f6ef5000d47b6b84ed058252aa =  ~I9897cbf9d7cab759f99f5f8f4bc125d0+ 1'b1 ;
assign Ica32690dbc9ea110fefdce92260b125c =  ~I9a6c1ff6dde5141849e4aa925140ebb8+ 1'b1 ;
assign Ic431d9383cce30b1889c92e2be4cb9d0 =  ~Icc1c25b229393361f1245c40f573b423+ 1'b1 ;
assign Ib9cca4c0e58373c26d5fd9f51f793898 =  ~I53b5a72e41ee53037ee3ae040799f401+ 1'b1 ;
assign I99bf0bc8ac20832b3724b2753f6ca449 =  ~I3cc25fb583118f45babf457fe78d5434+ 1'b1 ;
assign Ie701008f3c60c51ed72c5f964a8fc36e =  ~I20c046dd8a1265e12e902275b73417da+ 1'b1 ;
assign I3e2d78f8307a1787f8b2eccba94c7557 =  ~I1b184c9a34aeb6eda813d86556e235d9+ 1'b1 ;
assign Ic1b4444ab0df9745d29bf893d9b83168 =  ~I70e03db993e1d26d5814ff5fcd38ada1+ 1'b1 ;
assign I5f52dbf600656a8f5dc6b6b8a45ccebe =  ~I119dc168a44950d215af877eb81152fe+ 1'b1 ;
assign I7f307af79f45ad4b9511e3961c917078 =  ~Id717ed42457eb1d3f4e3edbf0dd72c41+ 1'b1 ;
assign Ie17a5be2a16d2efb98c976d7ee882535 =  ~I79d1f852a03bcc11d6121a12d8c5b86d+ 1'b1 ;
assign I5f19d2adff2f34a4bebe03f929a09c49 =  ~I769e650e49f152c0803b06232740691c+ 1'b1 ;
assign I3cd69aeed9e869a2096d6dced5c209a0 =  ~I1ef3c09b8481f14c3526224430a5f4b9+ 1'b1 ;
assign I359b6a22c9568a13b81670c741281393 =  ~I2a38d43a7e25050aa672cbf84a409aa8+ 1'b1 ;
assign I24ba99614df383c38bbac50ae8b4487e =  ~I1c2be5e13c462a8a6b07bca311582ce4+ 1'b1 ;
assign I7498bee46de6b1c946ce95fdcc89f6e5 =  ~Ie8fd61caf16aa0e504cc7dc8cec6f0b8+ 1'b1 ;
assign I0f644f42cabf871b71e5a82871bc7b5d =  ~Icd0fe98ca873ad6dacdf80dfdfc450ec+ 1'b1 ;
assign I71f9e059726a6cac8bdf0efcc0eadd2b =  ~I94e1ab698dc93ff0764dc5c1e62179fe+ 1'b1 ;
assign I0c9b2c1da30bfab514bbb556ae7bd4c4 =  ~Ifd48363af9abb390a72991fbdd6f7877+ 1'b1 ;
assign I7918b2e37e96aee94fbccca7e0f75fc4 =  ~I44f79397a010088e4ecdcb9669f2efbd+ 1'b1 ;
assign I76eebd77eb77e0abcbc727d2c511370a =  ~I124b0b7d91cfb42b0d9722f3229c2d53+ 1'b1 ;
assign Ibb2288e62110bae5b2d3fe901974e5c7 =  ~Iadf1875c584adc34f7586a146184a763+ 1'b1 ;
assign I080f931dfef9d8adfb1dc1ee073eb64c =  ~I02d3f9982f02ea85f996bf5b5975b930+ 1'b1 ;
assign Ide1106431e3565158bd81ccd6b18f3a1 =  ~Ia6e1b39d83ddce053518c5ae9a5ca33e+ 1'b1 ;
assign I63df19931e8d28666cccd79922cbd418 =  ~I3308663053f4307d43ac66f43266f706+ 1'b1 ;
assign I9a7e4a59447048de90446f877eb06627 =  ~I87ad25dff6c0c9ac46b7a129cb575537+ 1'b1 ;
assign I0917e92ed84363ca92fd2074acd74eba =  ~Ibf5d40b7c46b50866f58f6fa23e1861b+ 1'b1 ;
assign Ie3eefdf7b5561a90a6ddd9e6aa432509 =  ~I0e3a9a3b38875156d15f697adaf95410+ 1'b1 ;
assign I56eeb10d11e886cff629457a640a1c76 =  ~Ie3f87d094e71e4a82f60e8d91cdd768b+ 1'b1 ;
assign I7a9eea89c4e76d856df44b6bdc332840 =  ~I793f52d174cd09fe000e8d0351753592+ 1'b1 ;
assign If8d8f4333e893788fcb9ec54256e5b7a =  ~I89ea3da7db40e7e6705020462b2d1df1+ 1'b1 ;
assign Ie4af0e7e04778d85f5dee73da33376a8 =  ~Ib2af2f1a928dd824f25b99f0b602753f+ 1'b1 ;
assign I019a4e997adf54f5f5ca651f80b7901b =  ~Ie3e887f5f1a64c37a10404d636212b45+ 1'b1 ;
assign I10294667f09abbfd4e2f757c414072fc =  ~I5c6a004278f155d33d0cc1b576c3b25f+ 1'b1 ;
assign Id4e8ab8f15b36bd27d1e4ebc5cbe1495 =  ~I6a03a4a548a0906d1a3e9ce47f3454c6+ 1'b1 ;
assign I6c93588ca9e7c623d75314da39e89a91 =  ~I542e525074d049197ac3904e6102f0bd+ 1'b1 ;
assign I1020412efc78d12a9ebcbaeb83e5dcea =  ~Ie0307a43ce71ba73d4c8e5ad556bd341+ 1'b1 ;
assign Id0b574f35a83dcfd4481a10043cd1884 =  ~Ib03e1d3a1f27721e4ea32629c2e86f85+ 1'b1 ;
assign Ifc577e5c2c7288373a8c5e3969ac1589 =  ~I782f4ab4666c9f550a2cfc943cedbe77+ 1'b1 ;
assign Id18a1a17c1cf6e8a2492aa73b62898f2 =  ~Ib991e16161d5c8b3b655e3c7c08b93c4+ 1'b1 ;
assign Id8ce8f636723b9f119bb86c25017e6b3 =  ~I72f8c6bad4bff3b00055aa8824479931+ 1'b1 ;
assign Ic29a18d8d504a2d5280c1d7771346518 =  ~I58e5100cc1e9b809e93125fe5d08a9d8+ 1'b1 ;
assign I96a79193aa2956b8f901d5fcc9cf65cf =  ~I0aa7056fdacd6022f328a3be49048856+ 1'b1 ;
assign I8c97a246c749fbef029f8b1671c772bd =  ~Ia2f40b5c49a2284fb6a234bf7472130f+ 1'b1 ;
assign If9ba9d221909ce7499725f6fd7d519f8 =  ~I8da184aee7953890f2c89e40744402f4+ 1'b1 ;
assign I53a7878f44253f0f1a82d9d27b1a44c3 =  ~I613ccfc7dad5627cde02fa1720244d01+ 1'b1 ;
assign Ie0e928125f9d3d17d123d97e00f1fc34 =  ~I080fc6c99e506e569b97433f3fdc3e60+ 1'b1 ;
assign I2bd0f77efeca09eebe82ea234e9fe638 =  ~I79aa118ef8ac0d9b13723fb1f5a7e4ad+ 1'b1 ;
assign I94f2e7ef9b3463bd598dc9049f6fb0ef =  ~I7e6e7601245ca5b3a58b91848e25a6d3+ 1'b1 ;
assign I6dc16510af6b61b79b339d0fce77ac24 =  ~I2792edda66743635b837aa3bec0c58b9+ 1'b1 ;
assign Ic655e213ab81f5d61a018d3ed7016b12 =  ~I085cc29465c945957d00cbcf804e3ae4+ 1'b1 ;
assign I2ffc4a604025a2f5c4e273c1d070a725 =  ~I74a8e879666bb216a331fd2ab723e37c+ 1'b1 ;
assign I1c76818a9a3b688ca897aa479f7d807f =  ~I7a90a43ed71e82862457d9fa40bd005c+ 1'b1 ;
assign I3bfee9d3d88f0569010a4e0101200c19 =  ~Ie1e7b4bd6201baa02b8d59cb0f6ffb8e+ 1'b1 ;
assign I5d4738755a26beb6d0f61dd3dec0f804 =  ~Ib7b7cdc22b22f276b1c021abaa8fb443+ 1'b1 ;
assign I2f3c800091275bcb72d1a2a38fba53f3 =  ~Ib58e33f31be36b28997ba05ef1004573+ 1'b1 ;
assign I378e67cca7c4ff6325683f8346963210 =  ~Ibec394e82f499e8d2d5a9524f943d6ac+ 1'b1 ;
assign I04c8915a7f4bbde003f7facc84435c1a =  ~Ie06ad127e475dc131859992bb5f350a0+ 1'b1 ;
assign I3f50b10072f38b6addee6845e6df9118 =  ~Ic494a58468b6a7dda76923a9475bf173+ 1'b1 ;
assign Icc60eb18ba740036d2a17f98f15cfb98 =  ~Ib82a2db86d03fe8538fa19d06e501dae+ 1'b1 ;
assign I1677daa18aa8b226753b1a887b9420d1 =  ~I5b64727fee9d0825a4ea83261992e489+ 1'b1 ;
assign I36bc2d4c9a4480daa9b0944c08b50738 =  ~Ice7e502b9c2b797719448fde8376087a+ 1'b1 ;
assign I38419a6905f50135a6783aacca0384dd =  ~I792b4f73ed7139b8761443cbc0833e39+ 1'b1 ;
assign Ib48892dcb0715987289662a14672611e =  ~I278d57d1964cbf3339db450926ef4782+ 1'b1 ;
assign Icd9c94f929dbc71c9b836fda3019630b =  ~I9c1a08b61782ef6c72545504693ac54e+ 1'b1 ;
assign I5d0249d9a772805b3fba3f3c7f5d35bd =  ~I363594fb91d01abca7a2b7402e352fd0+ 1'b1 ;
assign Ie97341deb6fb24d49eb8b96bd0fd3f35 =  ~Idd284c75a230f4b97d5acb98a8e38b2d+ 1'b1 ;
assign I17dd788f9d8e91307b6b1ab7488f9ce2 =  ~If040df53a6410b263f5b3dc3090631c4+ 1'b1 ;
assign I92ae370022ed107b152b10fd0aa3d2b7 =  ~I31df60ffcaea9cee63b920478cb058f1+ 1'b1 ;
assign Iebb39f0d19ec1208bbfba6cf67a3bfc7 =  ~Icdd2f6ce69b389fbf712e45bdc0a0257+ 1'b1 ;
assign I81861f6bb8bbbab6e93407cfb4a852b8 =  ~I8971b250393b397b94db38b9fd0fe501+ 1'b1 ;
assign I217b2e3ca0a534fc5b1910adf3c1b57d =  ~I9199e5e8fdc0e2c62ad1d62fc4d873cb+ 1'b1 ;
assign I8429b08891dc56af24c72ce1b7725457 =  ~I6e03f71fdf20db836c5772658a050e9c+ 1'b1 ;
assign If96747262303f6c5c6b129e39224bd23 =  ~I2ef49f893dbc8581725ca0f6d1c3305c+ 1'b1 ;
assign If7012457af15c405baeaa1710319b541 =  ~I8796f168c892ac60c38a0a7f1e18035e+ 1'b1 ;
assign Ia0a0229ef71b85195352bb664ea4e4e3 =  ~I64a26e5117c8f3ab95bf0dfa97427243+ 1'b1 ;
assign I42aeb7c23accc2ca874c7f8221c3af93 =  ~Id7946a0299ced3ba00f6c3e6e664931f+ 1'b1 ;
assign I7df6a95bf51f40693c439c6df36510d4 =  ~I5243b90640ea4680de83021601c85c39+ 1'b1 ;
assign I8fe65f9c344d7ec8657f192abefc3fb6 =  ~Ic8301fceed328cc031640ecc4ff34803+ 1'b1 ;
assign I4d75c95d34d8d8aeeb528456bbe136e1 =  ~I6e852c94b6105af62ee85f8adf77fa55+ 1'b1 ;
assign I43746054a38c9521f8da9db9d0e91f99 =  ~I7d98c5c2a54832b6368ce60009208eb0+ 1'b1 ;
assign I0430ac2a4b2b2e2fc7f8154bf946553c =  ~I7e42f2281518bead81a6d18d2dcbd1a3+ 1'b1 ;
assign I25dc807fd55b81c9f24fd0d1edcaa758 =  ~I63c126c978154f2d68b11f08a938dcb4+ 1'b1 ;
assign I7881184f1779b9fd4fdf329c5f7664da =  ~I2ff7719c35578b47720cacd9ddfd92eb+ 1'b1 ;
assign I8e6de2d692a307ee8a5a4b2a9265a633 =  ~I480599aef36967a670155dd77120a37d+ 1'b1 ;
assign I54b2b18ab051b468808a3d0fc4bc893f =  ~Ic000b2c844de484b8f30b7b84dd6234d+ 1'b1 ;
assign I37ee86e2ca32832862cb57efe76bbedf =  ~If0e25df151db991185f992eab5d5be99+ 1'b1 ;
assign Ic95f2fc697574803c0f7fa35c2609f0c =  ~I2f533699abb7a997160bf4ee4cda3efb+ 1'b1 ;
assign I933a30c52c9bec5172530b2d739a3b63 =  ~If6b33cfc6d34e33fbb18e08fb4d8a5ed+ 1'b1 ;
assign I7bbd7df18f85197c22fe8cfe37312af6 =  ~I2ea5423dc8726fc0217899e0f406a1e9+ 1'b1 ;
assign I50d5ada7c91c7af16492c6b41151b68f =  ~Ibf3f4f8a04cbacc9624ca5cc73bf7069+ 1'b1 ;
assign I32c8e7996b3473d4906c40018799a16b =  ~I9ba53c36934ab1c7f498241a79cfbae8+ 1'b1 ;
assign Ic0eacd5a4812ad7ae3fa251ab2db4694 =  ~I106a25f18536f96782927bf3bc2ccd72+ 1'b1 ;
assign Ideecf8ab87d28a840cd93851169ab05b =  ~Ie5cdad65e918679607cc5f816987b736+ 1'b1 ;
assign I1ac6775eb38457b7962241d2e7336b0d =  ~Ica6dc9ded8756fd6f82eec4271e246c3+ 1'b1 ;
assign I2ecaa89698604fddd863d7e28d643a57 =  ~Ica42ac6ca5813d0d1a67f14d1248437a+ 1'b1 ;
assign I273e0fe9c51c8549c8dfff393ca2e4e1 =  ~I13dc6cfc75ef846c30e5dc1dc5305d59+ 1'b1 ;
assign Ifb1fc76002f6920a1f44c7b1bbcd0020 =  ~I33e784182dfb4af39715788b1ae98af6+ 1'b1 ;
assign Idf6d4e3aa753aa396a9bffb27732f851 =  ~I9e1a66805348d2e5bbf5e2316187444b+ 1'b1 ;
assign If14ca1f5d1c2977f9da79eaebaad1bf9 =  ~Ie9619916a96d218cf5eb5f3a4995d0e7+ 1'b1 ;
assign If8f1505d9f10e30bd3320f500d34932f =  ~I02ce7969c51ad141df227ed7d18e74b1+ 1'b1 ;
assign Id32aa77c6406b35a00168bb5452b12fb =  ~Idd73461af0d75c4d820f7f8f0f419e0f+ 1'b1 ;
assign I9a73686acefeb361337511f6943b036b =  ~I3df6c2cdccb2a82c58c1d81b00af7786+ 1'b1 ;
assign Ib6eb7ce5a070f3a87bcf0e18be8c855d =  ~I97f441fc5ffb88efeb5ed66b60f07a7c+ 1'b1 ;
assign If69b0b717c35d33fc8c0e59b07eb9edc =  ~I3194a235eb652c8d0e4307cd056e5e72+ 1'b1 ;
assign Ibb0d73078b779585e6b0e228391ecb96 =  ~Ibc315f6c79ba2bf336ee57f2e5f7d776+ 1'b1 ;
assign I2894546e399fe3e33d7579772a1310df =  ~I937a54f5cda99a7079c7fa46b4ea26f6+ 1'b1 ;
assign I97f99a266267859aed199b278a430417 =  ~I49c99afecc613656cd1469d8c1e98936+ 1'b1 ;
assign Ie18cc792329941a3654322376a937d8d =  ~Id76ce0333f43bf7bccf1ce48e25ca69c+ 1'b1 ;
assign Ie914a99f08d60b74c3c36a632a4ca9b0 =  ~I2c77f9644145219005751f7a4eb71aaa+ 1'b1 ;
assign I82916e9dc3894ad88e12de01a68d6aa5 =  ~I5cecc266272eef88cda88c1df9bcc37e+ 1'b1 ;
assign I6cbf576b3d652e34c0221f8316b5a392 =  ~I776a0b1b5c14afa21b7fda3c2cacafed+ 1'b1 ;
assign I9141b2516d7f855cd186472780af7b67 =  ~I84860b1f933339e0f90beeb3d666393b+ 1'b1 ;
assign I07bf32ed72de9c02abf700c64853af61 =  ~Id24581713f1ecb767db39d5154c2f5f4+ 1'b1 ;
assign I52663a2999fb9571834d517538691b6f =  ~Idb0eae2f0e1dae1d56251d64e2c51f9f+ 1'b1 ;
assign I8dcb88c94506367aabe8d7ed62cc56c2 =  ~I2e3ca4b130e6d3d92385928a28644452+ 1'b1 ;
assign Ie676a4bee61154145391d9cc473fe91d =  ~I7922d80ae333dcfafde31d294f0eb4d8+ 1'b1 ;
assign I9502c8fbf6b48749bf9f84a89a937dfe =  ~I82de04cd2dfef5616efca4af26d7c561+ 1'b1 ;
assign I0c91e540e7106f32ae59491d8ed1853e =  ~I7ce384520525b15d24c2ef6f161213a5+ 1'b1 ;
assign Iddfb8a8e261389eb4a2a10880c19446a =  ~I56aeea71c7bd19d47620cf36adf3f115+ 1'b1 ;
assign If0d55f861d4b3f0970c529024ca142d5 =  ~I138e1a6db0c6649bc023cc36d81d5b47+ 1'b1 ;
assign Ib054f5d3f5cbb29a053d0e50c23cb3a8 =  ~Ib5e8b1c4dd9b5dad56b59cc11c87a258+ 1'b1 ;
assign I1d65e9f97e93de8cc2a5dd532f8e482a =  ~I86f785e2d5e8d6c08fad1d334c7d244e+ 1'b1 ;
assign I3bdeab8c87325d46e45d9e2d44756934 =  ~I9a6c8efca218c724da4ee4c1087d58bc+ 1'b1 ;
assign If9228f7ecf19c41f4bbd8dabd0d5816c =  ~Ia30e8dbc6974ea94b763842e8dffa633+ 1'b1 ;
assign I9e3edee214c4937d2aa462d3cffa624b =  ~Ifa60f45f4d8848eb0b89f5644ec69668+ 1'b1 ;
assign I9fcbbd2e81b006b50e2d35ed2627bf83 =  ~I0aeb4b93cfa6d62ec41b7e6dd0287dd0+ 1'b1 ;
assign Ie16f3d50ad5e5581ca099549db7232d2 =  ~Ifce1fc978fb5b0187593f46f53c3b469+ 1'b1 ;
assign I6345e93f3fa7f5eb2008dd41742afc2d =  ~If3b6de7c919c5d53a0e191a75bd7e574+ 1'b1 ;
assign I698b93e10073b5d29357cde4bcac9dbe =  ~Iecce594e6e99b0c05fc845144a664b07+ 1'b1 ;
assign Ie7ced910d84655790823e6173a5a314a =  ~I2c8431500ecb25619d2884a2fb4260c0+ 1'b1 ;
assign If6e3b6fd1810f6964e9024329d7cb3e3 =  ~I217c710f7ef39035546efcbb043f63f3+ 1'b1 ;
assign If1045908c6d7476bd5507e57d08c406c =  ~I1b4236130cb1879d885653fdd9eeab4e+ 1'b1 ;
assign I4d4f6705ed77a16ff31b34bae0d8b6d9 =  ~Iae0f7c13f1564d63b4bfdc152ddf4111+ 1'b1 ;
assign I70a492396580ac1143d8a2f4b181e873 =  ~I010592496030d138a3a4245d00069957+ 1'b1 ;
assign I2fade32b5bdf245fa15289620dae2670 =  ~I9d7f47a6289a16448221d61f301586aa+ 1'b1 ;
assign Ie0dc166f57fea074496241a32cdb6015 =  ~I7b8ed2953170c4deadaeb33a6ba165d4+ 1'b1 ;
assign If6a2518891412caa6d6d507082501f1e =  ~I4efe9eef6a48aeb0a9ba4e0ffd9906c3+ 1'b1 ;
assign Ic9912e5a838a377b26a19d22148a64df =  ~I5a8466bbd83c39dfbeaa6399e3fb3337+ 1'b1 ;
assign Ibc0fca22d16444bc17877106ca772c31 =  ~I1ab96ffa948dd09bcc4f748c6c2575d2+ 1'b1 ;
assign Ie4291d233597d5d676a80fd62d9bd208 =  ~I016f57568eaf00b26f8a22100858c158+ 1'b1 ;
assign Ifc13b798d76aa70ec1877c275fb31d36 =  ~I1fb995e302f4f1ba493ff85f39938175+ 1'b1 ;
assign I57d6637f0bdab578a790e4a12ccaa16b =  ~Ie643ad235307c60f1ee96dfdcbc8c2a8+ 1'b1 ;
assign If8ea04fe685b4f20cdaf9a84984d56fe =  ~I8dafdf2c780082d8dfc2961b3447f104+ 1'b1 ;
assign Ie0c86f20c28bcbe410b191b90d29bf76 =  ~I3a2841a0f5e1b42556f384231ab0717b+ 1'b1 ;
assign I3dc5d3f66726e15968a70cbf3d3b656a =  ~I2b00d0e6facf01274c0c3446bb0e1599+ 1'b1 ;
assign Id674686e7ac37fd6f63846f9a9cede19 =  ~I2c645d25871b70dae5b2c283695d5130+ 1'b1 ;
assign Ie2ed9668d13d219c60f2e0614488cd42 =  ~I540a0e8968a6a82aca775a81ef82b520+ 1'b1 ;
assign I98abc995ff89934534543be93c6e3ffa =  ~I5b95bbc82e6d8d87421efe3f17b97ea5+ 1'b1 ;
assign I579cf9386ab7b08efa204d735335e462 =  ~Iad81f5e5e728ffdec6296b2aff668d75+ 1'b1 ;
assign I9efa4d729d10a6b7cc335fb765ed032c =  ~I960a618f63372da74581b8c352f3e618+ 1'b1 ;
assign If9191ebc8e88d4e75f0f35897ebb1421 =  ~I4f5325f1601acde10018d1fd0aff4d35+ 1'b1 ;
assign I3511287cfe69d5cedc5a8fbcad708437 =  ~Ib297101fe456520e72cd9d208af44eea+ 1'b1 ;
assign I91812179d44cb675b90d477f33ec48ad =  ~I73a21342321a9d81a0fa5308149d72b0+ 1'b1 ;
assign Idb04a1aae91fdc477ca38ed66789ee88 =  ~I2a486524f4f53b3454ee02a8892d4fa3+ 1'b1 ;
assign I566054aece562960590ee28b157e4a3e =  ~Ic6c4e4e6a9ba43a3354f9f3192ab069e+ 1'b1 ;
assign I7b2ffb762cd9ef7aa8ba224efb75c46c =  ~Ie3cdee3560bd06aed84dac5fcd2a259a+ 1'b1 ;
assign Id90bbb642b0f4434d8a148a28b6b2f65 =  ~I584febaa4c440fd9353108af36d3a5c6+ 1'b1 ;
assign Ia4e297e35d484b15adce7e1d67f582b0 =  ~I515e78507d7419ca14d77b6d52f75a78+ 1'b1 ;
assign I84996b1d03b692f6f736fb04c7f91e83 =  ~Ie9578453a57d2b3b9c3b98844044b5f0+ 1'b1 ;
assign I83078cc7857fc17b30f640854a4d6be5 =  ~I1e58b3062097a46d8d590232b40278cf+ 1'b1 ;
assign I94bb467129904032736fb13dd636c600 =  ~I3af126eb28c67797ce625b0d82943833+ 1'b1 ;
assign Ifa76758b50f439170ecd6d86ff898bc4 =  ~I130ee1a8acacf4cae8818cd8320d050d+ 1'b1 ;
assign I9d831dd976e8cd5d8f6a6818601e6424 =  ~Idf92dd09c29ce8e921b2b34089550586+ 1'b1 ;
assign I474774ae149804412ed4aaf1cdcaba88 =  ~Iba74a64cc1d2ec3c83a4061db298ad37+ 1'b1 ;
assign I964cdcb4e6b49a62d30c2a2540851317 =  ~I01364c233ca541914d790354515aa5c1+ 1'b1 ;
assign I6df268bc9f85ce88674a9165664ea84a =  ~Ic6a8297308a63ed3113008a3cdc76358+ 1'b1 ;
assign I74fdcbe9f49f7bce1f5e31d956c5883c =  ~I6c7ee9d0bd684a7f54bed3d52452219d+ 1'b1 ;
assign I4a1b8453cb7a21745d5f74ad05653ed2 =  ~I985ea87550ec8a222e6af621589e186d+ 1'b1 ;
assign I9c53b478b2011fac0615a152fe60d5b6 =  ~I6836a7d1e006d7f7556edf8b31aea32e+ 1'b1 ;
assign Id75dbed8f1a5befda32c60b994681013 =  ~Ia7a356a18af18ec131b9df46019f3e58+ 1'b1 ;
assign I378a59323b74623c5524f854d6e11226 =  ~If3a7e111247232c47ceccb5e05338312+ 1'b1 ;
assign I080bf885464a0cc948a4450e9f7d1d26 =  ~I5f38d1665294b2d3c18f9cd888ff60f1+ 1'b1 ;
assign If769e73adea227de1fd85c2e89d0ba08 =  ~I10290b9576bf3d8caf90583a388226b7+ 1'b1 ;
assign Ifa6a34b83225e9d9b28b14874c4444e3 =  ~Ief36236305fc1521c5bb4c60753a676a+ 1'b1 ;
assign I584b1d4d6fb7ee4f20ad9c96715cdf90 =  ~Ibaa0539fbf5ccc979511c09c061cf494+ 1'b1 ;
assign I265f9b91fbb62164e589dcf96818c4f5 =  ~I95664ffd0ff13c2893421032149f24d2+ 1'b1 ;
assign I3d59a47c88227734cf6fc0d6fd30db11 =  ~Ie390153b3b7985dc63d65913de215377+ 1'b1 ;
assign I6144b6df2c87ea0948d730343b42129f =  ~I704147dda658f4a03627dacc1c91dd48+ 1'b1 ;
assign Ia7ca7400e36ea572fba8e19bcc81ecbd =  ~Ifb09672d505898f081aa13c95fcb88b5+ 1'b1 ;
assign I302e61b49accf5db556b87517f2341f5 =  ~Ibb5cb89097dd11bf292d5b5a2422175b+ 1'b1 ;
assign I5d9af1abff6efe3a55c6568d936b6ec7 =  ~I4a305956b18d6ad6901d2c17e99f2bab+ 1'b1 ;
assign I8cde0aa611c476b5112edeb8f17f15bf =  ~Ibf5bb3b9eb1812383db9634fa9a27ad3+ 1'b1 ;
assign Icaa40ec40d6d26cdf70bb5ae7d492e47 =  ~I66b37d055c3735f011095ee4b1ad02ed+ 1'b1 ;
assign I8346f15d822cacfeecbe5d75412cb53f =  ~I43e71dd694d97217e242f267248cd594+ 1'b1 ;
assign I5ee364aab320ab40c0f65feda6f53b18 =  ~I4baa925db1ec733bd4bd25d9dc873e23+ 1'b1 ;
assign I1f0ecba054900f96cd7100741191c5f4 =  ~I547928c9db7acc531af251264d576ffb+ 1'b1 ;
assign I4faf2caf62966416118a54015908c889 =  ~Ie4ce634b2fb62a20781f8a2e8fddc762+ 1'b1 ;
assign Idd0329980a36f87859150530ab44b52d =  ~I0e90e96ffa64c2874d79110b622994bf+ 1'b1 ;
assign Ie66bc10dde27f08813d4d347fd7cf6ce =  ~I767e37e3c6f4224eb07adeda480ce253+ 1'b1 ;
assign Ie1d8b3ea7c6603cebf2f9adb776910b7 =  ~I75fcaf2c65b7e63adac834054850c6d6+ 1'b1 ;
assign Ia37488e9a50cf5cc08de74ade676db96 =  ~I5f1de2dfbd79204ab2db9b686d6a6862+ 1'b1 ;
assign I08aa45211cab01d567cd5eb172fd2f0c =  ~I8d01de6be4091dca2589cef625c05229+ 1'b1 ;
assign If4ff0c63ec1deb46412858e496451a01 =  ~Ic09e773899fdd208c0fdd874933b2cec+ 1'b1 ;
assign Ife7bfd15fc4c392b5d2288d9a4e879b3 =  ~I24a3f9fd851c4af70ef66bfcee44af65+ 1'b1 ;
assign I24ac26debafd03c7333d174e8725afd6 =  ~Idd31807ecd603db8c719349a2be1be40+ 1'b1 ;
assign I99d80ad68e2563d0f78a0e3bb82c5328 =  ~Iaf680cae40d1adf7649da12b31a2be0d+ 1'b1 ;
assign I9943733ef305983c629565c881054bbf =  ~I22d948171c1a66f7a28d5e51007700ea+ 1'b1 ;
assign I7cb4420bc55c03a6500f5228d31fe43c =  ~I3954318b2392a82f2da71a0ca1504497+ 1'b1 ;
assign Ic4d19dec464359c0a9fa75148fe90c73 =  ~I15c78b909cbd04fe25820d777655d829+ 1'b1 ;
assign I44993416e1d22613dbd78402c37a934d =  ~Ia529c5ec88a9f6c14ceda5cad56b346d+ 1'b1 ;
assign Ibc9b94a9dea471805cb442ac6904bc97 =  ~I5b73c81f28901705f6ee26d63847db0a+ 1'b1 ;
assign I917d9f9b144d3bffafc77bddae7fba6b =  ~I1a9bd3f728db23b679639e5657ced179+ 1'b1 ;
assign Ibc91c6c3d56bb8a14e22909c43ffec51 =  ~I57ca72784a7c91cecbd694ddd08bcb98+ 1'b1 ;
assign If7c2d3eddd96b47b6c2aea8b27c8c7f4 =  ~I50f31ecd3f2b498cc7b759efa057f12f+ 1'b1 ;
assign I4df093ed94d26b058e97db550e347e3c =  ~I8ccaf29848defdd264f522642968fa29+ 1'b1 ;
assign Ie90303b0326bee4ab203a8cf1e643da9 =  ~I808ea92ee1340876cf1d2c47255dc2fe+ 1'b1 ;
assign I19030d352fd059156ee42c66f9270beb =  ~I3da806790125328b626be1949f71267a+ 1'b1 ;
assign I36767a902c53a384128ae1443cf88963 =  ~I55e59bc1daeb8b2be3d7a1e4b272df93+ 1'b1 ;
assign I868dffa3f07407f7996bb5bc596939b7 =  ~Ib0ffadc6a0091ceff91ad1fa435413a6+ 1'b1 ;
assign I7d928be164d0dce8b1322ff230c053e9 =  ~Ic863f139e6bed2d06789a07c6dedf6f8+ 1'b1 ;
assign I98be4971a8a9a08abb3ebe474d7f0c6d =  ~Id0e8f6ada5060a911090f76cfaa3c6bf+ 1'b1 ;
assign I779e70dea33201e9237f29681ffd5e27 =  ~Ibb8c9b8fc9b58f5f8a6ad342934804a8+ 1'b1 ;
assign Ie2262914042172ab7e08599278f36af5 =  ~I9323a188737ca54c2dd553cd99bd416c+ 1'b1 ;
assign I4001323da8f7956cdd480ac2d56df929 =  ~I2694cef38855f496e7ca12f42dfdb9fc+ 1'b1 ;
assign Ib1cd6731034887a0a55e405c9db3e8de =  ~I75790b4c0b1f6c7935f5cfbea26407d1+ 1'b1 ;
assign I51aa496e8c03944c28a908102514e6f8 =  ~Ib8b366c47e56a49fc53ea4a9e1ebbd99+ 1'b1 ;
assign I6415f3996318472532e161510ccc8ca3 =  ~Ie1c86256df2bc6c4dad41237eca41986+ 1'b1 ;
assign Ia11b671b59240988737979328c472812 =  ~I7c9e3f97a94f9a078c209a1b84ff916d+ 1'b1 ;
assign Id4fabe0165a117a402dc14f2f3ec626a =  ~Idde839d34403fdbba62671b83801ea8d+ 1'b1 ;
assign I57238f501ab7278b308d76211ced8cf7 =  ~I824e23c3e43434e0a7bf8c8b8e0de597+ 1'b1 ;
assign I9b257f8556ca4e5402637f01081b78e1 =  ~I0f83a2c488c229e971030fc66ce212f5+ 1'b1 ;
assign I2e093412a9fa3972cea01664389d8c27 =  ~I8fdda3dea7a63fd6e57f70365d7b6571+ 1'b1 ;
assign I17907fd8c6975c8c642535ff929221a6 =  ~Ifa2fc30c14c549339edc65c3670d90a0+ 1'b1 ;
assign I3c6577b04ad56d864bbaa2c048323c11 =  ~If69bb1bfa10ca7dd37ba57485c3429e7+ 1'b1 ;
assign I6f0c341c05eaa8f35bbce4521f6e8f94 =  ~I2ab0738fa2d5916d77a81b9da2315376+ 1'b1 ;
assign Ib72ba950ecf9ae2668374f6633a67ca7 =  ~I50a9ce776ad2ccd8048b56ce101c80d2+ 1'b1 ;
assign I3d7c72d725f4563bb562e2992093cb02 =  ~I9c9d0332ee7ad6a3488b7e39bcb06ca2+ 1'b1 ;
assign I813c881ac61a59041be3be78f6a466c8 =  ~Idc155814976f0aef9b56b2bb3d52b3a5+ 1'b1 ;
assign I866510e7dc721fa5aac312bc5ab5ba0a =  ~I2e02fbd496d08acb3ad3359b49b9f680+ 1'b1 ;
assign Ib4432359f97849dff6ad3e0f044157bd =  ~If0f8b3dfce99a5a75c2105d45ccad985+ 1'b1 ;
assign Ic86aa6eb1b4dcc2520309089b43292e6 =  ~I6790223e6a7cf136a7e2b261ba4fdb0a+ 1'b1 ;
assign I0731115afe5c15bcf131f7ef4f05802b =  ~I6a9643afea7a6cc9b94806ccc8e84c0f+ 1'b1 ;
assign Ib080b8fd34385aa7986dace4afd95267 =  ~Id3d19d7c2b941930478a7ab01049e390+ 1'b1 ;
assign I134890b77451d0b78afc7402a6a28048 =  ~Ib0a25312d51cb6aa1741f7e425bc5cd8+ 1'b1 ;
assign I956da75f13433c1dd7a3cbd3b78922c1 =  ~I44dd1b66f5a9a6b0b976d3d61d6c5cbe+ 1'b1 ;
assign I440b26c9f1b9ccf70f97c9d5f732d38e =  ~I3ee456f2f0e7f447ae92b7523136adb5+ 1'b1 ;
assign I5e3a441faca44bffc4368d96d8fb0bfd =  ~Ic110e2a08b550acd3c8bda4a1bc2bbae+ 1'b1 ;
assign I21d7ba25247a87a1a9c245d0d1f553b0 =  ~I3f87162d2874effd66a82f821aa6c73a+ 1'b1 ;
assign I55aafa8162cfc4fccfae68cf78cd1c2b =  ~I660ea6d341fcb38f108270c08d82473b+ 1'b1 ;
assign Ib99c25f0d8d6493cac4d5c816884c704 =  ~Ic128d603fc08affd2f3d0ab3425710e5+ 1'b1 ;
assign Iee7c9f0a0e8ca127efee008b4874edbd =  ~Id5372641727970383a59e08f550814b4+ 1'b1 ;
assign I17b4a3baae65161387f472037ffc6fc4 =  ~Ie99ad992d66880542dcd330ef6ccee04+ 1'b1 ;
assign Ie7b7b202a968fe73f6b1e02a044414c5 =  ~I9ed0b194f7d210d57c54b289e01c75e6+ 1'b1 ;
assign I479ab5c0e483c36267d8248340006666 =  ~I227828831c4ad21b06ed00fb5781b0e3+ 1'b1 ;
assign I777bfe165e25d7fde4fc950f23db7b84 =  ~I09d5ad12cb836adfbb4833ee80fad2c9+ 1'b1 ;
assign I146d505a34ddb8d65e0a1769f623a7fd =  ~Ifa9c94ee94e4beb2e7c8d2d57150df41+ 1'b1 ;
assign Ia85239bddc04bf50bcf037ed2f76d7ac =  ~Icb88e59e194db215382e8e949603a9be+ 1'b1 ;
assign Ia7306bacf3c2b180d3261a5c1f0f4a30 =  ~Id4ebd28aaf1076acec266666f88a02ad+ 1'b1 ;
assign I2018147b86e47af5842c4f29d047d157 =  ~Idf0a0bd862167392357501b3233a8d8c+ 1'b1 ;
assign Id17a85459845f8a8be694c4bf1fc29c9 =  ~If94cdb867ea0fc2c5578b16aacb1acfc+ 1'b1 ;
assign Ic012b15584d9d25af38f83d0526503da =  ~Ib8c066b0700941a4fa739820ff12b948+ 1'b1 ;
assign I7f09bd4a45143a036ce04af11b9927f9 =  ~I11e0f8dc46b286bafb05f901f968e1ad+ 1'b1 ;
assign Ica32f94af6e6f3eaf2b724a2173fa463 =  ~I608537f5639d5e0cd3e80453e21f6f85+ 1'b1 ;
assign Ib750bb83ddfbbad2a2be8d1c8392b4ff =  ~I0e9d8db1bb6347c9507b645132308b3a+ 1'b1 ;
assign I3906ece39480f96020717c6243e8ba4c =  ~I17033b417fa383a2db41d157df33d9de+ 1'b1 ;
assign Ie68ce21ade07fa53c30ebf27216b03f9 =  ~Ib7f45dbcad513b4dafee60f33622b0c3+ 1'b1 ;
assign I6cc6fa167c0d2b4b62ddbeecea175ed2 =  ~Ibfbd8e00e00272f32428c7b4a3c53050+ 1'b1 ;
assign Ibddf3468ae7c27d5a4b1388e524aa9c2 =  ~I27973d1d4e07eaa49608d6f6975d0a93+ 1'b1 ;
assign Iadcb2b3acaac2e1bb505c65d3cbe4235 =  ~If77fcedbcf99f89045de87e5cae45d8a+ 1'b1 ;
assign I37cd96b8b0a4939d9a70098fd8bcf452 =  ~Ie8f8691820e7a560db8116f38dae5d49+ 1'b1 ;
assign Ib34b169dcc76daee2d1aa2b2a7513af3 =  ~If0b19af59ad851aded19970494514034+ 1'b1 ;
assign If36fc316d6ec7c7e09eae77807b37099 =  ~I98b8e05818925a4b65082fa57affde83+ 1'b1 ;
assign Ifd214c332218ac5c0fe5aded4b952711 =  ~I69317e8c556ed67630829c990f8b74db+ 1'b1 ;
assign Idcd0fc8f86e2b6f03606b818b8346e5a =  ~I9147d103cf235310393f9339f1cbb376+ 1'b1 ;
assign If486aa8ac2cfb46f936714812cc760df =  ~Ibe0b2cab6e2d3f3cc8baf3623ff50988+ 1'b1 ;
assign I2d8e5b5fdbda7d599423c38aaace6658 =  ~Idc64f1443dd2497dfaa223cda3fbd682+ 1'b1 ;
assign I6d0878fb7ec75c0a26be4dbba62f80dc =  ~I6e37e92b812099985436851da8a6ccb2+ 1'b1 ;
assign I16a16ff0e8a6685a09803634da429fd2 =  ~I057df2bf67d5580275654bdc28b40027+ 1'b1 ;
assign Idb211abaa54ac26e7379c64a63f7d07c =  ~Ie87a151c8b90942a899b8167bcb34afb+ 1'b1 ;
assign I351205eb71acb31b59d2b4470f0ba28c =  ~I735752035af159b48f53d8302bb33c21+ 1'b1 ;
assign If5660c495bf7690252783d888d1ad6e8 =  ~I1f26bc7cb30a9659a638e2ab65e1f187+ 1'b1 ;
assign I3a5229cb8e44a15560b5c7bef96e65cc =  ~If39a50e88c4a7c43428c1d15b0bfbbcc+ 1'b1 ;
assign I889b9b0828e97fe44d8366c5ef71a8f2 =  ~Ibf966c12f049d603361ad32f55b0a2c8+ 1'b1 ;
assign Ie23062e00e39ead706f5b6ead233747d =  ~Ie1b3ed6d3fdae47669d3c4cb8af8d969+ 1'b1 ;
assign I8a2589544c75ecfdc31d28912c639695 =  ~I4ec6c8d9e87224ecbe7c69d92f9419c8+ 1'b1 ;
assign I5c21c59147e9c3a74c7cbbb6f2a23919 =  ~I2acb34de8c3fc53117a7ea4f9ce7dd2b+ 1'b1 ;
assign Idacd78e24408e432abbbfb0c447fdde5 =  ~I7fa4009267e80ea7eb71194843c3b22b+ 1'b1 ;
assign I0e8b171fe5080485a7f4fef83f1f1528 =  ~I6854329daadea2734e52180a41f56bcc+ 1'b1 ;
assign Ib22c2bd76e6c29cc2f1440885bf24b7b =  ~Ifca16aebaf75b2990188de201e4536fd+ 1'b1 ;
assign I149559fccd9def4ec1ead1fdcff3c7fd =  ~I46cc26afc8475f2fb290eefc95a542eb+ 1'b1 ;
assign Icfa8fed3239748abca27a5fc17de79c0 =  ~Id746d6515cec9e60e7478898a09787e5+ 1'b1 ;
assign I2ff115fa483f080d93bada49a9566b33 =  ~I09a3ad636db96e00adac78c3c94bdaaa+ 1'b1 ;
assign Ibee4f3cd2f516c29ab68e07a640ab65e =  ~I28b3baa225a5fd602c9fee9c948ae58b+ 1'b1 ;
assign Ie495ab560f59ad038992c573de7d2f5b =  ~Ibe12ef0f56d875c7a44030882deb0e29+ 1'b1 ;
assign Ibd812def78c3a9c02f9ba45cc0413711 =  ~I9bd9979e4acc4944227a4bd62b910c1d+ 1'b1 ;
assign I98166634dc80201b0cefb01d9559c228 =  ~Idcfa802f458499150055dbe4b1ce8146+ 1'b1 ;
assign Ic2f03a980b5f0b042853ca746abab22b =  ~Iee010958cc3e9389cb8ecacff84fccee+ 1'b1 ;
assign I2807a88097d2683ebdb9e0e785e3af02 =  ~I3d74b31096917c53757c829a67cf06df+ 1'b1 ;
assign I8bebbb3a676c8506af0768516abcd740 =  ~Ic27031a9654db9459815fe0ca35408db+ 1'b1 ;
assign I31d380f34691c9fe9022035f233b77e2 =  ~Idf6ead2c37f75f3cde1d4b40cd73db00+ 1'b1 ;
assign I1ffb5675c98ab5b3c62b24eb23441473 =  ~I66a56161cd0ed67f65834b9eb0e94d17+ 1'b1 ;
assign If56424546ec4f3445853538207ea864e =  ~If6de990e26ca9e8efc009188f8a5a4d9+ 1'b1 ;
assign I31a49be4a34d9bac2e0d815097439772 =  ~I8d866786bb2dea06f5b30f6ea80cff17+ 1'b1 ;
assign I6b96a2498078953e87de223aa2236d50 =  ~I01ca9a1d4901ec9b2a64300617ce4cd1+ 1'b1 ;
assign I79bf36e298a85a42c7432f877055f0b4 =  ~I2dbead35e15afb9affaa6ad4edd3829e+ 1'b1 ;
assign I90c070b9bde5da05e8a5d25d2de3ba6b =  ~I83c57653e24cc09214075b04b06bad83+ 1'b1 ;
assign I28d0e4e6d772dd58d845d91952ada300 =  ~I56b9c1f555b24c2dc197168decfdb8d1+ 1'b1 ;
assign I7232b4e277acc6f1acefcb606ca24508 =  ~Id5c48111f1b93de2cfe89f92fd182b43+ 1'b1 ;
assign I32da124c433c55f692ffa4734d0dc8fc =  ~I32908c3c90ed6488357ce4869e8a1721+ 1'b1 ;
assign I56e487db14eeb8d93f494d2f11b57a49 =  ~I16b4601f2e07e6cecdb5a030178e75c0+ 1'b1 ;
assign I94d3c02bd5b8e84926d4b3c2f56efeac =  ~I0ae08a41ebd0e6b402a4980478087bb5+ 1'b1 ;
assign I0c35b2e9176f9a06e26ca67d036411b4 =  ~Icb57267a66f117943e964dd6420d7a58+ 1'b1 ;
assign Ia6ee7b70d0b7fe7c346760b1784e50b9 =  ~Icfa47fb87b74106cd3814adfce909424+ 1'b1 ;
assign I7ce57c278c683ad045526e49bcc47412 =  ~I63067cef0e1a348a3e6d8cd9bd88b907+ 1'b1 ;
assign Ie3d3e681cac0bb919946ac27057409e2 =  ~I10aa5ba0f53632578c0e1cefa4bf4fde+ 1'b1 ;
assign I8ea0a8cdd6506c982ad75f23136bcebe =  ~I427c0215d0ac047e8402c20610676752+ 1'b1 ;
assign Ic812f8bc775c5ee6a83e2b9aeb22b2a4 =  ~Icf4efa87688bd1b80437686eb0126057+ 1'b1 ;
assign I0f0adf7fe957b9a68772bd8a1bc163d4 =  ~Ic373f785ddd1bf8eccce263df5a82c87+ 1'b1 ;
assign If09562f8d82bc1dea7c38ed51523a889 =  ~I56f8e8d2d7052af26528530d389b6dc1+ 1'b1 ;
assign Ib0fd21d66cd89c4e5c95fbc9c7680b62 =  ~Ifb145bc18d435fb66779e7415417bc0f+ 1'b1 ;
assign I5a2b2bfadc638fe3fdc31136a8f09a8d =  ~I62a6e0c9952d6c6e6095e2364df93078+ 1'b1 ;
assign Ica914d8c556285d6b90b35747065a6e5 =  ~Id6405c2b2b9aea6bc457f1064d5f3ffa+ 1'b1 ;
assign I00c5d739bccb0ab6d05da70fe51aafea =  ~I079df9611bd81f672f2ae028bf267995+ 1'b1 ;
assign I18e448761bc014ce490b766183350312 =  ~I096b226cc511363946a39307a7d97867+ 1'b1 ;
assign I1b5920f488e9469bd416a6af3072a30b =  ~I4cc42c5a75ef339510ee0e86fb44e16a+ 1'b1 ;
assign I70b41ffed4b6d88ddff219c567b8e968 =  ~I680c01c3327cb9372a42c1ec5b4193e3+ 1'b1 ;
assign I935e083b4561da7d015e98ca7f02854e =  ~I83451a072082194ecb3f9419edd728b3+ 1'b1 ;
assign Iaca9ef263bf220d786242b88c994fd21 =  ~I52ad85b6a1c822ca8c2459bde8fbd510+ 1'b1 ;
assign I92169291959eb33452b79bfd32618cbc =  ~I1c44d2ef638825862061a8ee1a0a2f95+ 1'b1 ;
assign I126dabc3ebb9c4157adf62b57f217bd0 =  ~I8fa1fd425809cc39cd8e2785773c1d7a+ 1'b1 ;
assign If4433b1ef2eb963cd301946958b69884 =  ~Ifa22335f04d35680eb8cfec8f862f357+ 1'b1 ;
assign I67ac5b9b794787b3c4738c3366689871 =  ~I6aff673c27811b81530453906312aa9c+ 1'b1 ;
assign I4f022d70078c412bdbef158f750d3da3 =  ~If674ac0540f457a21235664c213d4923+ 1'b1 ;
assign I6be6165385f6a77aeedb88f2baaa9cab =  ~Iac223ac498bdcf2cb2514582aeaf76f3+ 1'b1 ;
assign Id1f7fe91547e158e1d39edffb1421ff3 =  ~I7f40931ab78ededfcb52ccaac9b81282+ 1'b1 ;
assign I7a51924134902612db53941390891245 =  ~Iab7c8dad0ca20eb0988fbd99f25591a8+ 1'b1 ;
assign I45128b9e29dd2fdd94a78fc5ffdff2b1 =  ~I3cb5f890a5bd3daaae34c8dfb6ecfc49+ 1'b1 ;
assign I7f1082408c8ebb5be18e8f71ff9510e5 =  ~Id80e145586d7e539a6514dd67ebabf6a+ 1'b1 ;
assign I655ebf19c2f4b3dde716668f9ce12e59 =  ~I01e09bc554768f30dc490041d19b4da2+ 1'b1 ;
assign Ibc9d493a507122d92af42d858cdc4c61 =  ~I0196f7df6f834ae20c4fdd127e66104d+ 1'b1 ;
assign Ib3d3103e5ee4feb160a97c7e26f7102b =  ~I4669c4f256c123a0fcceb55c1e72193a+ 1'b1 ;
assign I6cc56b119e72175df3b7ce64dc3d9305 =  ~I4a02ffa2a79df824f406909aa189a404+ 1'b1 ;
assign I57cf4a9378f1cdd94a1a5608dc57e05f =  ~I3117e5029119e70846dff61d746699e7+ 1'b1 ;
assign I4160ab1aa18e8151c0a5c23b9edeb907 =  ~I1e4e705b3bda1451fc384cd934c0bb52+ 1'b1 ;
assign Ia1f183f2d904d006e46399424e06c614 =  ~Ib5bea8e0072de3de2c8431ea6a35dd51+ 1'b1 ;
assign If979702738671323995e56108bc9376c =  ~I7d9d94022ea95ea01cddc237f3df8cb8+ 1'b1 ;
assign Ibc96fe0a6bf1f95036f97c7d44fab575 =  ~I3f0f9aab07427fa81fc3096c6b6d3d6d+ 1'b1 ;
assign I755a38220a693ba43701d30e7e9508ad =  ~I12a7983041f9c298d533bad58f41d24b+ 1'b1 ;
assign I896fb82baa9647a14f4b5b1ecfa70a15 =  ~I78503880e5c96ec0a03c75266b1226e8+ 1'b1 ;
assign I23d1c973d7a2048353fbb68e4a294c08 =  ~I8adeae445b33f634977957bb1a2259aa+ 1'b1 ;
assign If9fd1e08af14f2fd4ca363383f48580a =  ~I73bd13f381d15e0b0198b60cee44bb42+ 1'b1 ;
assign I8f3782f78d88a5c3bc93709564999b30 =  ~Ic8b651c2b043a4a6e4cd259774322230+ 1'b1 ;
assign I986d61d79ce31f4677f3293339db6ad2 =  ~I76979d7df582f9306e796a03cb540963+ 1'b1 ;
assign Ica4d93d9fad21316002008ade5106a9d =  ~If61d4585986757a525c54589ec93d8c6+ 1'b1 ;
assign If77592d5d8bed32477fd690341e543d0 =  ~I1bc5766a4a3cc2b468ab8ef62eab691c+ 1'b1 ;
assign I25b70c6b830cbfe1b41d8f289c751924 =  ~I21585169e5fceda643bd03fddf8153be+ 1'b1 ;
assign I2a5d65eeffa18dd9af9fe36463dafd7c =  ~Idb2990946f60939136b3bfddbc7b1671+ 1'b1 ;
assign Ibafa6e10bd4edf5d224fdeb2f9adbf98 =  ~Icfbf703890f684bfc96decc429deaa04+ 1'b1 ;
assign Ifc25402bd879bc5c43b4945b60cd4540 =  ~Id5bb42639a1c1c1d67df1c89a14a2bfc+ 1'b1 ;
assign Iec48da6882325d8a33e0e0e845eb18a0 =  ~I55b8ef91d667c1c1d9e58dbc86a2288a+ 1'b1 ;
assign I0fd05e46862fdf8e614afaa3fd478602 =  ~I17ff683da41b469c8c8b82ee32a7378a+ 1'b1 ;
assign I6253a59dca81842d9ab6e58cf204abbf =  ~I51f10296c38872338ec7df35ccd520d8+ 1'b1 ;
assign Ib18d64bc58b354358ee6ac16785880e2 =  ~Ia59ff33765ddf4aeb17f90a70c01d76c+ 1'b1 ;
assign I28689b693a7a5f761a1f252aa3ef3b67 =  ~Ibf97abffb1ec40f2f0e099a814e04ab2+ 1'b1 ;
assign I1a4e6d12f9776d5e61094e0b5edf71d9 =  ~I3efc3271e18a1e350473dcf3375088aa+ 1'b1 ;
assign I8e1ad23b7ac662bb827a83d3709f0adb =  ~I1efd1220ea9100f2fb4f169ceaf462a5+ 1'b1 ;
assign I000ad2287813072cc18dad933758f2ab =  ~I9af399f27c8e2b62b7f3fc6481ef9318+ 1'b1 ;
assign I7bc3698b51b89ac38ba5f4b5428a0c96 =  ~I171bb4ee9be2f92e4d82997108572426+ 1'b1 ;
assign I78aea1705621e2845a331c3e61a8055b =  ~Ib13cd76c20fcaf95f26f4914380c4fcf+ 1'b1 ;
assign I0a31314c3580f5f9e61e79c133e5d794 =  ~Iafb219f1c8c6883e01fbfb4c887c8d6a+ 1'b1 ;
assign I0e274fd7bfc0388fef95a8ceb939ee91 =  ~I94fc9b0bdd2b0a89a9f6351f1fdd4ff5+ 1'b1 ;
assign Id6f39ddcb73d3f4ec081a365d11d1ef4 =  ~Ia9ceb45f33402293c162cef4037ba007+ 1'b1 ;
assign I807770bfa86d160459d6ec3c0f4d6a0b =  ~I0fa4e12e62e8a30b3b8045143b344b4f+ 1'b1 ;
assign I31c89b8a11a3090bfd74b112cbc474bb =  ~Icec1c637d24ca277bb2e488257e92a40+ 1'b1 ;
assign I79b82cb1bfc72bd5a9d313b9e9c9203c =  ~Ie9aca08b988fad20904545fe070defd5+ 1'b1 ;
assign Ib1046ae03c9a77fd2c0b3e9838e9af87 =  ~Ie82304b2c8583f967649475e309e68fa+ 1'b1 ;
assign Ic63723fd43cbbbde51c233a3cca15d3f =  ~I60da0fb8a2c0669d5f9037ae99b23565+ 1'b1 ;
assign I3abbb59abada1aec6941185f95f738bd =  ~Id8c19a3547c17ed513d2d857adc66885+ 1'b1 ;
assign I8d5bd7039a77ce82ce0f6cbba9c2a076 =  ~Id74984743844e9495ea0f528a391f4b8+ 1'b1 ;
assign I527ad0b9382dd7b6e657dc1a32d8e472 =  ~I9edcdd5b927b3f6b3a4c7cacebeb4a82+ 1'b1 ;
assign I8de02f32e14e719f4930d99743c04a20 =  ~Ic89597a95f50382cd3a2730896735d55+ 1'b1 ;
assign I7614dd5e9628c761dd9b2a512cb1da98 =  ~Ibb7d203dfc75bf6211b09ab94877f93d+ 1'b1 ;
assign Icae7efa4742dd0ad943ee1f67b0c9b14 =  ~Id2f2e6837c83973cb2173454433acb88+ 1'b1 ;
assign Ieb1854b79e9a2bc6cf5aa1c319e8e753 =  ~I1259d5918f8d65b4b22ccfef22fe3afa+ 1'b1 ;
assign Iff50b77f300183ca59a67ccbcc9573c4 =  ~Ib84e8c6e7fd9d7762e6e7e508d5ee40a+ 1'b1 ;
assign I4868604f8178663de759d4c63dc6c4bd =  ~Ia032017912715abde99ffdf5ba732c5f+ 1'b1 ;
assign Ife992a151986c58df4cba79b6bc4ac0a =  ~I55c310bfefb635448ef9c25c5d15987e+ 1'b1 ;
assign I9ab973fb74d9fac5d78eb8fc2c7ecf36 =  ~I92c0f229cf7fdb2cc0fe4d84f4d9b11d+ 1'b1 ;
assign I5ee7916e859b86a98538659401685016 =  ~I5570eb486d238fd96f9a59b174f5a22a+ 1'b1 ;
assign I48c284cefb8cfb5a938a8f23ce4d7f03 =  ~If6f01d24acf4a8b38bdbb1b366cd9a47+ 1'b1 ;
assign I5c1fc666b77a689478654dd29519f458 =  ~Iff29fff36064aa4f9d339d4c62956e61+ 1'b1 ;
assign I38bba98b59184c75ba3b27e1dcf52182 =  ~I818d7cae6f1b80ac452dbfc073ccfe7a+ 1'b1 ;
assign I6905b65403c16b0211643227ece536f6 =  ~I77ecfe991c6ec778495d7d5e5e442eca+ 1'b1 ;
assign I3ed34401bba9d5f229bc98480aedd9a5 =  ~Ie7c6a56e8b6f7756bb5a24bdfd6a855e+ 1'b1 ;
assign Ib4d05804277cddc7f00ac17ac14f5325 =  ~I9f9bc8eb8b2978a3dc529c34516fdf75+ 1'b1 ;
assign I41babdca6d3fa462849592d37b0a7998 =  ~Ie3c0e5a4b00a92357a5d37e527d59b61+ 1'b1 ;
assign I58cfec706dc929ebfdeaca6e01b00c0a =  ~I9b9a9486420e7d4aa105c48dd50aa74d+ 1'b1 ;
assign I7efe3c5b2fc69840a79545e0399ce749 =  ~Id12199a504f7aa298fffaaedd1aacc99+ 1'b1 ;
assign I70e3eeb2b3966676d16a6aa4c85753ab =  ~I813691fd8ea36626d32c8d2562163f32+ 1'b1 ;
assign I2a32d545d1e7beecc7531174c7e8dfbc =  ~I5fd3aaddc3eb8afeb82768b45e2d53d7+ 1'b1 ;
assign Ib8fb40e4ba0ba1f5e9f5a99d1271ed06 =  ~I1ac281eab6c7459e835fe992142b7857+ 1'b1 ;
assign Ica792cb9850a61fa4a8bd8a4b6c6ca05 =  ~I49e5078c9161e8bee00fb76bc00b5288+ 1'b1 ;
assign I779e5997c66649d6d54fd7f0514c47bd =  ~Ia697adf14616bf50d6e8178596b9fa7e+ 1'b1 ;
assign I5aa578b0c2831453683fa44af1878cb8 =  ~Iff3128a26dabe63b015dc6afc98a85a9+ 1'b1 ;
assign I735d6229ef1a4ecda0a1f1dbdfb53fc1 =  ~Ifc04708ee5a7cc2b3f1850db778fa42e+ 1'b1 ;
assign I62affd47512c5e8f0979244115624d97 =  ~Ia405859c9dff67905b2e91bcbc06259e+ 1'b1 ;
assign I14fe27afb3df5531b18dc9604e8dbe65 =  ~I2fec8f62b28575e8f3af756db66fa232+ 1'b1 ;
assign Ib1b1626c84dad8ad13c058f921ffd57d =  ~I98e97c02477032ead66dc50f3f274e5a+ 1'b1 ;
assign Idf4a4bdddb88c21c5afe10a02373a6eb =  ~I9f2dc5add3a4d1e6eb3116c741cd2f82+ 1'b1 ;
assign Iadefc2a3d07ed4b2c3c46b2ab5dec252 =  ~Ie122f7d8a48d7ad29d998b6a14b8e70f+ 1'b1 ;
assign I19315957077b037ffc6415dbb06ef789 =  ~Ib5576c996062391f44066d893dd5cb91+ 1'b1 ;
assign I1f9be09334407fc86c83a7c127e17bbe =  ~If931597aab866a74c3a3ffb1cd429583+ 1'b1 ;
assign I28e17a5af7a7286a2643100d6d058dc0 =  ~I79878bd69ed53785b8a5f025a2a00a4f+ 1'b1 ;
assign Icb2297c397bfe56be251ffb6b249a020 =  ~Iefb0a20652954fc2002154ea874c120a+ 1'b1 ;
assign I64a48984527d660002f1f82c376c7a84 =  ~I646ca66e4e9f24b4fb75b38bf293b4cc+ 1'b1 ;
assign I238b5fc70ce9f05b6322a2691b3a0207 =  ~I051f0d4c44123e3637b84a32c9a00a75+ 1'b1 ;
assign I00c16e7ad3821981032a42d5baa767b3 =  ~I1876f9ec3f6f637ee40cdad7cc347f6f+ 1'b1 ;
assign I42fd5b094da200b33036e6cb8c7d0286 =  ~Ic3d6b8dbec6cf92a9b6a17fb2f75dcd4+ 1'b1 ;
assign I98b7e26a0e9ec9ad750ff87cc0641a73 =  ~I7d89f1db7b1015d34363ad781374de58+ 1'b1 ;
assign I3ec904916870171bf837e162d1030052 =  ~Ife217ec4da1f1477bce034cb3545160f+ 1'b1 ;
assign Iedb11b97900b7dd769d31f8a89521975 =  ~Idc5e5e98508c94b87a760f8eb36fad41+ 1'b1 ;
assign Id0dceec6497c9f13ada07138986d4145 =  ~I9e72b0c823f297535f13a1b3072c2776+ 1'b1 ;
assign Ibfe7d9bac29b8838f20cdcfe8ef7da0c =  ~Ia81da7c58d6636ab70e0cf3e263a12c0+ 1'b1 ;
assign I4d6c95605595942a34573d6ed55eb326 =  ~Ibfc69ef08382c79e30cfafd89bfeff69+ 1'b1 ;
assign Id6d8f32958dfa1a98958a84e7f1aed02 =  ~I2d2afa9165b7121dc8289e9e6cdab5de+ 1'b1 ;
assign I971cdf9ddd1bfff5664eec35f22da335 =  ~I065052693fd8ca87614feb60f7ef37c3+ 1'b1 ;
assign Idd8bc1412a0dc5f489ef253a6164ceea =  ~I13344a81551374f665cbc17c7e94296a+ 1'b1 ;
assign Idbeec36de0128e5924e214877c82bf11 =  ~If5a1d2de0715fa87d191ee5f48171676+ 1'b1 ;
assign I50a9cd240979bc56421bf85011ae99ed =  ~I02b256f74ee86b42ff1eba5e3d242737+ 1'b1 ;
assign I6437095f6bad2d4fb2fbe0361f60bba1 =  ~Ic113fc051eefaef846f440e98f2f8913+ 1'b1 ;
assign Ie9b6eb3bbac26635aa00c38110958d46 =  ~Iabeab9bdd0bd82dd145218b563b5dac1+ 1'b1 ;
assign I9f34e81e3ffb85539a6273babc2a732e =  ~If9ce0a09e3a4e816dda002a24319ac0b+ 1'b1 ;
assign Id0a1ab8472d704001e0eba0317b117d6 =  ~Ib5a7d72c36e41754033a64fbe0718784+ 1'b1 ;
assign I9e632217cd0561d8faa28e4b8850d995 =  ~I41df12c7dee8526abf92b8e98965fa06+ 1'b1 ;
assign Iedeb5b7b2fa8acf1ea083102678710ea =  ~I83dfbd224e7465a6fd769e407182829a+ 1'b1 ;
assign I972431d1f5af0bdf4828e4f85591e358 =  ~Ie57bba5092ec318456365b81b36aaa65+ 1'b1 ;
assign I1f41024b715d8312944ccbf70e95bb40 =  ~Ibcf043d24474ab8c1002d15fde2d7da2+ 1'b1 ;
assign Ia6bb5ca05f5d0af452c994dd50004e1d =  ~I2e3385871c6ed8cf9519f273c8a19fda+ 1'b1 ;
assign I9a1d1d1c862808f9a769cbdb3bc634e1 =  ~I664917b9f44515bf556d69ade4ca408c+ 1'b1 ;
assign I9734eb86f4e73ba217739baf5cb1b13c =  ~I28deacdec0fbd0bce49b654c2620ac38+ 1'b1 ;
assign Ifc0fe00f86569956df72d8a960337e8c =  ~Ibdfc4852c620f573f929584e6b816f35+ 1'b1 ;
assign I223341a807a1d555f759632f67815159 =  ~I5a69b2bbb63ab919ea2270503cd326f1+ 1'b1 ;
assign I6c1f5cdf5f2917118941f4af14d67fef =  ~I2eccd8d60a19481fa595566f51c7aa4e+ 1'b1 ;
assign Ie84e88fd1aa2a0b90aa1715fcd27a329 =  ~I49eb4bba42440657fe04b711eedfa67f+ 1'b1 ;
assign I558f70d7039a8bb58d8ea3f72e43dac0 =  ~I9ed8323951af0de78ae89153cbf9e9eb+ 1'b1 ;
assign I9924269ed3de12f1f2a28893c7f95292 =  ~I1d00816529836546b514f54b1275d39e+ 1'b1 ;
assign If1153befd1396be2798cc14535ddeb8a =  ~Icc58b9a24fb9ef7e8fa5f13a2cc0a0cb+ 1'b1 ;
assign I9bc447b20687fb3e7eff45792bd4dc3a =  ~I9339aef608b029175b488e82f5b3f1bb+ 1'b1 ;
assign If590520f01e452db9867a8d6d5dab29b =  ~Ibd2f24860b701ab46e0c436d774e43f9+ 1'b1 ;
assign Id93ee7d283016ab9b0aaa21237237c54 =  ~I37fe66ec8927f27f646b304500400ccf+ 1'b1 ;
assign Ic1cf03baabaed466fe532e4db3a9ea78 =  ~I4bd6a48f494cf633a857b8ccbd67af68+ 1'b1 ;
assign If3031f9aa8f6eba90eac12db7839fefd =  ~Icd7a7566438dc67e77f138ac814844f0+ 1'b1 ;
assign I0dc2708970ca2b6c092273b6626bacd6 =  ~Ic3d4239413333883dd926c7a42c0a87f+ 1'b1 ;
assign Ia58944aebf0b4f0a7d76a1444fced9de =  ~Ib8298d1ead61bc00eb31599b3087d769+ 1'b1 ;
assign Iedd8e69679d10e05f2889f1d71cf0e7b =  ~I23dbe33ce46f94d3dff1e6d391305609+ 1'b1 ;
assign I90f0d471914a2333b9dc14d6d01cf927 =  ~I138286817f424c76e8a4f30540b0530b+ 1'b1 ;
assign Idceeb22013af64b6bb9f0d773e9ffe9a =  ~I30c645a78b900306864a1ab23e923bde+ 1'b1 ;
assign If43574342e60a625fb6bee5a495e88f3 =  ~Id88681d0fe3ea62530166938503db05a+ 1'b1 ;
assign Id285f055275014d9f23d35f91879afa1 =  ~I808008402174fa4edf42783135c0c3a9+ 1'b1 ;
assign I8c803ab08db372802117de4fa4e2a187 =  ~I3ad4d02ea2e52a49b6fa4f1da9b58149+ 1'b1 ;
assign I13ba48a6b360f3cff5f37ce60cb735c6 =  ~I39486eecb7bbfecf26573a7a5876feb9+ 1'b1 ;
assign I4547cd1dad45dfd01e335e8cf20eadd6 =  ~I21e8ea20029fb2cb62103405b81b21b0+ 1'b1 ;
assign I0a305655b815b0cc159ac1c5f4ce30f8 =  ~Id0b67fa451e276889e02779ddb667904+ 1'b1 ;
assign I3633737da6b74284b0ea9a06c3f5875f =  ~Ic328d25a58ec4559b753da3bcff938de+ 1'b1 ;
assign Ia949c1b338d1cba07cf6bb6572c3e322 =  ~I49c44c2f2522e086c2db8a00647ba35c+ 1'b1 ;
assign I9a0185f8400159415bc0ad6c38284041 =  ~Id4152a04385391294f4b8a18df2cb9ee+ 1'b1 ;
assign I3eeffe43e7deed7ee77a7f5a3bce3cd2 =  ~I5b0213a3df61e94fd0b744a8141f7502+ 1'b1 ;
assign I85af0c31ca7002ae569d9f5ce39943f7 =  ~If0ad11ed403cbbed68614b01e2a3793e+ 1'b1 ;
assign I3dfb8d2fad83fbd807fbfc6330c5b857 =  ~Icfa1170bc73534bee13778bc3b88a2f7+ 1'b1 ;
assign Ic12be21bcba5fa49437cc44dd8a7f064 =  ~Ife1bd938a0dd06d8d3cf30ff41a303b2+ 1'b1 ;
assign I713a384d022d3012e3d0019f5c4ac077 =  ~I4a09cb1b99b476fa6fae0bc44c41a041+ 1'b1 ;
assign I80550019479d0323d0dd7e7d0f767d83 =  ~Ie08cf323944813e4b9e2d59a680ffe8d+ 1'b1 ;
assign Ib8a866f080dd997e0b6c93b6c844d1bc =  ~I85fc307fb52d58550eeecd33bc4207a4+ 1'b1 ;
assign Id542de206d736ee3769ea0bd037cb627 =  ~Id00dd13741fe621d0a240bdc92318f55+ 1'b1 ;
assign I77e6cdb09c92492c3303d0213de9c291 =  ~Idc8e891fd432df75a4eb133ce35ecec4+ 1'b1 ;
assign I788c33a9f94b26f4ce0f515891d06f90 =  ~I2a51cada20cbd14f7d5a289599e68b53+ 1'b1 ;
assign Iaf7074c2b570a296fe2ea8a5a7097ca0 =  ~I65a701d1e083e501544bb0fce24f0c4e+ 1'b1 ;
assign I8964c6d3f8e02866a6ad86553ab05d99 =  ~If3020a9109ac83274b5bafac18d176de+ 1'b1 ;
assign I2aa25edaca90c9dae8ed63b48d333c17 =  ~Iaa6bd55038c2ae911e4df08f707c55f5+ 1'b1 ;
assign I51a440917c7ae23339bec6f8a745c103 =  ~Id49065cedf20e13abac8971534bb8b0e+ 1'b1 ;
assign I56ce875e4619d4d8d6ca2fa0ddee91b1 =  ~I0bb64952d77b59803a561e14b950b9b1+ 1'b1 ;
assign I80607da8f92f5a5d2e4798a62a7b1c5c =  ~I01e295a6ab88c6f34b44efcc32a23233+ 1'b1 ;
assign Ic4dcaa520e26bac40b3876f02074f856 =  ~I2acf864d587b7681ca0fb6e2e2bea617+ 1'b1 ;
assign I3b2714d34081a3b6cccc47fa1638e72e =  ~Idfd0410b37713e8808f8bea81e2af881+ 1'b1 ;
assign I2db1d1ee8f546c00e512875ce2e13cee =  ~I02861f333b5adfd4962356cdf5a11f23+ 1'b1 ;
assign If80a6bb104ff3b2020e909103c104063 =  ~I4ddbc3daa65b111cb0d45e13d62cc292+ 1'b1 ;
assign Iadb72cc5444816fbd132256493930bb4 =  ~Id363d158feb8fec19b5f3d73d84f0068+ 1'b1 ;
assign I3a8ec1ad07bfada3d2c6ffca88b8b678 =  ~I8ec9b7a6e65e727abbed336ce240a4cf+ 1'b1 ;
assign I0aa042b86d9f68d22a49b4eb480a9088 =  ~I128fa1e99b7eb9b6905c2cfd26b95ab4+ 1'b1 ;
assign I89a387374771b68d87d7ff2dcc810829 =  ~I93d459b6da42a205c91c48622f0c5032+ 1'b1 ;
assign I2935b3d5c3bba4dddfc7ae03fa77b229 =  ~I1243cc8d5dddf7dd65b40c0b3b958b9e+ 1'b1 ;
assign I4e0c0248f4aa97d263d64dfec36e3aa2 =  ~I238df7e09d42bc93a972da349a00f511+ 1'b1 ;
assign Ia2871d7493b2727d2cb2fbab596b7e6a =  ~Ic658b2afdc7331653fc84d6372d47418+ 1'b1 ;
assign Ie57adae8873946d6c706074b52a49786 =  ~If39be111eb101c9c983fe0baa9a1cb18+ 1'b1 ;
assign If5ac85646e4b339a19af658f01d0a17f =  ~I9d19d5b7d8b256c1707de97a4549c458+ 1'b1 ;
assign I1c092426f34be030b3e020f40517b0e1 =  ~I6c2fffe204091f7f64aea16b0ac98769+ 1'b1 ;
assign Ic719b72ad271bc7c077067518e6bbb98 =  ~Ic4ba4d2e5c12d9f1dd233d64929f1072+ 1'b1 ;
assign Ib87362230682c88d68a0ba70e25f3c20 =  ~Ia9dec5831998d472d11429e5a7e60ed8+ 1'b1 ;
assign Ifcf097a102f8dc1f912022fed893d222 =  ~Ieaaf52c1e663f260292bc1529718d681+ 1'b1 ;
assign I56483ca3fa550dc59bfa347780cfef7b =  ~I37061896a09588a73445deed73d3746c+ 1'b1 ;
assign I4aa9f61be376458185c3235442c8fda0 =  ~I02f25b80945b6f58193fb37add3da2d8+ 1'b1 ;
assign Id91fde1007d47258273299de80721390 =  ~I19045602bb77f12666ebd44f813db2c5+ 1'b1 ;
assign Id58498c34aff2e1216c189b9df88822c =  ~I4abdc8d5318d2922696a8aaee46ffa59+ 1'b1 ;
assign Ib52e0c68caadcf4dd9636a84f5460e53 =  ~Ie139f2048f346d82623c8fc6d40c9acc+ 1'b1 ;
assign Ie19679053b289bb5a0aad570cc81bd14 =  ~I8d99c96e203fafc81d13ce5aee925d75+ 1'b1 ;
assign I8862c5ef45b723c9abf5d0ab6854a900 =  ~I37b0bdeb3cc54d6a97720c4912c67832+ 1'b1 ;
assign I30db951a07af96a8ddf59360141b9a6a =  ~I08257e9e6c74c60448e22fb9855f0825+ 1'b1 ;
assign I4855a0a0c6426d33014ce6a4c96965ce =  ~I32188cca2fc715698fc05b0fc6506434+ 1'b1 ;
assign I362e8db1791718290bd33a79b4fc0855 =  ~I88f1cbab9b8fa3802345f745d024931c+ 1'b1 ;
assign I773f0508440fb71d73fd82a372cc0a00 =  ~Idf548c0e78bd221bf9f612f27002fae0+ 1'b1 ;
assign I792891cecae468d7a87e12f2da62a718 =  ~Iedfd2e04f5740d283388639dde3ecdb5+ 1'b1 ;
assign I33303820ad094d7a0ab53bca722fc609 =  ~I7088c83eacff6f1dfb134f79d469c8f1+ 1'b1 ;
assign Iff98739de575e25104c0dc30f08912a5 =  ~I6f8431671331f4ca7ea19656e0677cd4+ 1'b1 ;
assign I1952614b64ea451e9d0646dcce5dd1cd =  ~I1e31259e267e04920cbbd16bd7aa18bc+ 1'b1 ;
assign I49c1a7d1c20a25496821ad80c7eff790 =  ~If54d9f8088e67e44cfa3026f5a520fd7+ 1'b1 ;
assign Ie2be17a55e79ca76350e033f227800de =  ~I6fd2c0746407b23aec5dff1e083f5fca+ 1'b1 ;
assign I737a5b06f848cacf0c8da4985c73c66b =  ~Ib2147a19b44d361da628a628fbfaa988+ 1'b1 ;
assign Iab160609bb21501aa55b662d2010357b =  ~Ie804d1f4b241a2de3e9d9c7c876d914a+ 1'b1 ;
assign Ief74f1a9d4a43ee5c9def7b83369bb21 =  ~I6cd1e6db57e06d8f5e60a31f48ae4809+ 1'b1 ;
assign Id144423f50751e661db3860a8487d004 =  ~I3e0e8832d5338423284ac4b2a0c5f3f5+ 1'b1 ;
assign I623352a4f6705b21d461d6b32e85c12b =  ~I6ac006d79e95e222cdc66754b67a08ed+ 1'b1 ;
assign I28d1dc8dc594977b5058b5bb9f6bfc66 =  ~I29087dda1a527842aeb3d35d66c853cb+ 1'b1 ;
assign I5371a83bf9d6f334cf8d1c5b082527e9 =  ~Ia67e5920bbac700dfee52cd96b15963e+ 1'b1 ;
assign If1605d6646fd267e701668a7245b3b44 =  ~I1f6ecd894d90547f661e7a3888d048bb+ 1'b1 ;
assign Idf5eb1ac2c5bd92fa08ed935ae298255 =  ~I3112e793c6e79e1f5da2776e69a34e3c+ 1'b1 ;
assign I44ce30330c4d2d6033a0a970dd2bdd68 =  ~I79152f32b45ed5b4a5302f6460707b01+ 1'b1 ;
assign Ic101b8f56ea1e25c6b752583a1b01242 =  ~I3d16e7d6b190639b88a217f19ac63233+ 1'b1 ;
assign Ib7cf44e681881e55d2d353280a6319d6 =  ~Ia1be780c686163cea54b62d6ede72dc6+ 1'b1 ;
assign I35690f724e964248dbb1e80fb1ea49f8 =  ~Ic398c31a2a6ca89d0236534589a5919b+ 1'b1 ;
assign I5affa2759148a6baf5b9f0cd3122348c =  ~Ie91c3202bc957b350d1915000564392f+ 1'b1 ;
assign Iaeea1f06ff0c6e9cfa43ba14420c3adc =  ~I687957f5300b0d4f50d6893cc556bf25+ 1'b1 ;
assign Iac5a23266c3b038b4b54a916dccdf3a8 =  ~I7816b368e8e8b8dd69383b2c9327120d+ 1'b1 ;
assign Icdfb7f52cc27b1cfcde90a100d29af13 =  ~I5f021f4a664205afbe0761af4c8914f1+ 1'b1 ;
assign I71484d7e00efa02a08b54a1405f2902c =  ~I69728004b59b5206a03a8e2087834f7d+ 1'b1 ;
assign I68a9b0607e69e8b3dae64689eb288a33 =  ~Ibbe1d623f8f5f3aa7fc70197acc6df5e+ 1'b1 ;
assign I2598c48aad48072a7f216b2ab56ee532 =  ~I4cb9f74288811592fd97fdff52bd6fe7+ 1'b1 ;
assign I796e3a193b1b66fa9a04ca60aee11ea1 =  ~Ibb471dbccd39d41e951e98348812e343+ 1'b1 ;
assign Ic96be7e69faf0f43b92618131cf0c98a =  ~I7f37d68f8ddcf8b4d5e99fb51eada873+ 1'b1 ;
assign I648afe4114ce435bf1d13e0ad54425cf =  ~I72ded7153883418a712ef967439d2159+ 1'b1 ;
assign If05d7e30b4717e0a1bfd20b90d0539bd =  ~Ie071e08299bff6bbdbe1f84703aaec08+ 1'b1 ;
assign I5fc356af8a62a1d739cb375fb851e90f =  ~I1b79aa38a39ccfc839260af89aa78e7a+ 1'b1 ;
assign I22f4c5403fbe33d18f97cf21786cdd80 =  ~I7384296e4190d83fb9d9a92cf965125b+ 1'b1 ;
assign I9a1b2b9f924099f1e57fa501ba2e33ba =  ~Ie03034ce6233ca24effe53a2c0c8f6f3+ 1'b1 ;
assign If6253af4ebc430e4937269a5f4989b29 =  ~Ic298f77f42fc1d41cce684790036ecfe+ 1'b1 ;
assign I0427d17423548dbb33cf792883b4be8c =  ~I805269f95afbeb6b93182f68868d08eb+ 1'b1 ;
assign Ie539faf01ae85253e399308fef98afd6 =  ~I881328804c45b06767af51e11182b27b+ 1'b1 ;
assign Iae6e7c42f250cd9223f18f8830fb177d =  ~I958993626e6e44e12f7c1e8026914680+ 1'b1 ;
assign Iff47ec1743b59d7f90e9042af7ce44cb =  ~If31528d1fc3a083ebc364e75cdd9c71f+ 1'b1 ;
assign I1cf4a55ebab332defa32d2922b885285 =  ~I4703b8d5a9033027889bfa8685e09e4f+ 1'b1 ;
assign I284913858691ad5724073b73a820047a =  ~I22d8e84d2db4b07111b7fdc6eef34cc8+ 1'b1 ;
assign I35626ca53adbbf0a3a71cc6fcf43bcb1 =  ~I8b7c6df3b5ea575caab7820c95974608+ 1'b1 ;
assign I0d74ef22d31abcec73c7c582310b1e6d =  ~Ia8aa76bccf7eb310a9356e8b7ea1609d+ 1'b1 ;
assign I15f4cf1aa0ad5ce2bda52df338e677e3 =  ~If9de547bf469b8424f1625e990f72b04+ 1'b1 ;
assign I6c5ca5e68c8844bb1617a2288b5bbc37 =  ~I27d51b2015ea9af9bc345adabdb07b6f+ 1'b1 ;
assign I44343a9491069c3c8ea4fbd6255a5a6c =  ~I93dddce2a0dc01ecb3039fac5cf04011+ 1'b1 ;
assign I1d8318b94d86e1fd28323a5e5684a37b =  ~I746da2c1d5a620eb7e749f72f0f04a06+ 1'b1 ;
assign I825e83bd88575868f4fcc9a8b8729663 =  ~I1e15f8d6fdb4ac732768d0cf73af829e+ 1'b1 ;
assign I3184a16c71cff80c8c90b40e45f114b8 =  ~Ib719e667d7ba857f4f7432a245f4a30f+ 1'b1 ;
assign Iae133550f8bad8357a73e7de1372faa3 =  ~I4c6eec4a0c46e4f5d7c9734df48a16bb+ 1'b1 ;
assign Ibccb4a43c410f698e0fff68553326a77 =  ~I95623ec1fd5516040a9492aae0fc2b70+ 1'b1 ;
assign I72dc7aa294a3af89101ea62a4223170e =  ~I69017b49c11de463fe6d881e5c96a1aa+ 1'b1 ;
assign I91eb3e70921e0b141a344bc57dfbc934 =  ~I4fb9ed32471aa614ce6923f6a2279b36+ 1'b1 ;
assign I1986f22f2269cc135c6ed28d35fb0bd1 =  ~I2f0bc217c8a39d71adc1fc45c10b81c3+ 1'b1 ;
assign Ibef24017bc71de9c002aafa7ce9a784c =  ~I0f1c6bb577ea2b8b2ab636e64378544b+ 1'b1 ;
assign Ieae3ed78fa2c45507066f4e20d96e956 =  ~I7a248af9d606c566e03977e985c280e0+ 1'b1 ;
assign I730fd25ffc7778fd4bb02d33cb3870d6 =  ~I0bf9d47bff47277de1e72518e8d88362+ 1'b1 ;
assign I9a32313f2911b797fb0848f7d97e62b9 =  ~I24b6f4f68f291dc50caf03dc902282cf+ 1'b1 ;
assign I6373e2d64fdb5dd77733b3e4bb405121 =  ~I79335b28eea15735f760b7a8b803e93a+ 1'b1 ;
assign Ib437aa67ab7c13b45d7a4d56ce9e79b8 =  ~I0b14b34b06cfa90539c2abca5639abec+ 1'b1 ;
assign I0cb5c7a759f4c75d4a675f9777f15c5f =  ~I26878777354945712f834740b17dabcb+ 1'b1 ;
assign I0ca91c1426ba14a7b47a081cb3becd19 =  ~I6cc5daed4de5950c02c0a57b993e22fc+ 1'b1 ;
assign I0737e0cc7453e328efab2277bb712ea8 =  ~I52c382d5b0c4829127c011fae402ce04+ 1'b1 ;
assign I456af863661122cc303fccb235f3c7a1 =  ~I46ea9871e867034daa2d0501038f15e0+ 1'b1 ;
assign Idc5916c4800e9f647d51c52444ab6fff =  ~Ibb8a202599550e87831647a93a14181a+ 1'b1 ;
assign I57aca70e2b8d126c120736b2606ed333 =  ~Ibb79f2ce0b6028ebb638fc6661444cf1+ 1'b1 ;
assign Ic6650a6d092b749b4498c08d69cf815e =  ~I0d0c07d65eda2eee01df9c330c0d6f4a+ 1'b1 ;
assign Ic2e3b8f91eb218650c7b9c515c7efe97 =  ~Ie6940736944bac9be609b8d58b2cb13c+ 1'b1 ;
assign I93a084aa1e6881ab8dc905dcdcdfd7ee =  ~I472a71363435cb3ec054e00f9123ae64+ 1'b1 ;
assign I8cba172573be52c5a90bd40e6f40a508 =  ~I553223e9166dcbddd1a51d0f92d68f28+ 1'b1 ;
assign I1cccfd1516af59265731121dde878116 =  ~I495309d795905a53b0a3d3daa4f1f9d0+ 1'b1 ;
assign Ia171bbefe2d20b4c058126c33ef28eb8 =  ~I21d358fd7673c4392f4e4b3d3a858b2c+ 1'b1 ;
assign I84bc44a5d53a8f66b985b70c7ec1ae7c =  ~Ia1a60175112362f015c5531f7c48b90b+ 1'b1 ;
assign I321b104ca3c818018d4b03adfe1110b9 =  ~I5644ece811bddcec04c9e3559c86109d+ 1'b1 ;
assign Ia79b8994da536c86634bf6f54a21145d =  ~I37d2f9d3f05cb90e2d45bd578299885c+ 1'b1 ;
assign I4df55ce80eec5fee295b5a0ae92bd6c8 =  ~Ie7d10f3c0f8b0add66d2cdd4435ccc88+ 1'b1 ;
assign I46593a7956590d870fe680228081a6d2 =  ~I3c37396a1cef2f9e42b8ccc126db6eda+ 1'b1 ;
assign I906e9da31de73ae45579607a014e8b54 =  ~I2f82390734079b8d289d48a6682cc624+ 1'b1 ;
assign If5dd1a1b9e3fc0e67a85da3183480aed =  ~I9061728c3163ae684e8c5aec3e807868+ 1'b1 ;
assign Iadfb1571c78c3f0c05e4ef498267df24 =  ~I672d7ecc28a788c2602aff76187aa568+ 1'b1 ;
assign Icebb43b184c2745cc9da9d01b06bc62f =  ~I660b2fe99cd0bcaac34e9540118b54bc+ 1'b1 ;
assign I6e4b0489ec7333abf2245a1b72a8923d =  ~I6aa263fc2a061d2c4059b08309f860f4+ 1'b1 ;
assign I24ac5dd30526c1d3bc7b941103a66804 =  ~If3aef2d755013d195fd44f734365d7dc+ 1'b1 ;
assign I33681b2292c086fe536dae2aec70903a =  ~I3ad2e0bbff17683824f575deff82c6bc+ 1'b1 ;
assign Ia373ca76c3b15a4148532b3822f82ba5 =  ~I5087dc4b32d29bfd7bad49026fa58a5d+ 1'b1 ;
assign I7d08adbaf66cea04be4891db610bca3f =  ~I8a7d893f3ef6d6a93ba552320d901599+ 1'b1 ;
assign Ic09ed51b20f411683a801eaad61657a3 =  ~Ic057537712e09fa794918e5cde87e084+ 1'b1 ;
assign I6a9af8c9009b5de47ebe9ee8b79d3831 =  ~I0cbab5173052c450504e3a7d15ffda52+ 1'b1 ;
assign Ife18e8a16d4437161b75a93e3dff1b5b =  ~I81ee40feb7abd0fec3faee653f778f5f+ 1'b1 ;
assign I0cde86532c8db1a32d9fbe38a40b91b8 =  ~Ia344347a85d4e6afafa2ee3487e65def+ 1'b1 ;
assign I49c8ec4cd33e6caed8ed7dab779e7ebb =  ~I038fce1597157a3d95bd9579cc2dcbc6+ 1'b1 ;
assign Idb86f95570587a0711d796aac7004c25 =  ~I546585b819c289d855cd098818792e90+ 1'b1 ;
assign I2d1373d0b18992fa46a9607a86d21520 =  ~Ibc3a6609765818327e79519f3e348494+ 1'b1 ;
assign I30f26e090ab14551cbac41883ad8a152 =  ~Id1c71a2a34f9e6239559d28fe2780907+ 1'b1 ;
assign Ib1b4e41ab25733d1d6dd54e1fe81a419 =  ~I1cd6cf5f8119d5e6b4ca40694399b1c2+ 1'b1 ;
assign I146c0d5154a6de44c0536de873904ccf =  ~I15e2a1b4356785d73e2ab5d51f1f5ec0+ 1'b1 ;
assign I8eb9d4839a478a4e28b45a549b5682a4 =  ~I803aeb29e66384bfc62744a841bcc83e+ 1'b1 ;
assign I2501ef991a59512c43693ba9d7db8571 =  ~Ib6e220dd4f54410239dd0c791d84a700+ 1'b1 ;
assign I38213f78fd4dc52f9d2c9b7b22136c1c =  ~I8a009007fec23f4d492b0da1b6b404fa+ 1'b1 ;
assign I49ce91ac152279af421bbc6c4d9b8087 =  ~I5f89adcb1ba235a74639eca119fb2655+ 1'b1 ;
assign I6a2b7bb2cb3ca2ab932c211a68dded55 =  ~I8fd2b001ff154e4760ead2df355c80da+ 1'b1 ;
assign Idaae6ba9da8754615a2c34ef859492db =  ~I581569cc2e63bc68a8466b07ca471b25+ 1'b1 ;
assign Icaca9fc70a3ec6c48c0e41f8168e2bb9 =  ~Ia9cfdea21a65b0270de42cef7ebbf822+ 1'b1 ;
assign I4f69b8ff834c7ab3194bc9390ce0f5f6 =  ~Id66a233d2e312aff939549dfa96a8cf0+ 1'b1 ;
assign I037cb596cd48c5533ed22bc32518d992 =  ~Ie479c12c25a1964c3804936d45725bdc+ 1'b1 ;
assign I94a89577951de90edc4f73b281ad7364 =  ~Ie30d8770ab7e6643fcb67463f6999125+ 1'b1 ;
assign Ib7493a1a384aebaa7999ff1fb867fc6b =  ~I4a17ff532c9341e80f7ed0626f728054+ 1'b1 ;
assign I2ceb9e423696539135c5bae5cc2d8d98 =  ~I597bc1ec224007a78c25f7eea24c2c3e+ 1'b1 ;
assign Ia6bbf236436b2ed22bbaae3b8849de6d =  ~If198ec15fcf66e97e69f88f718979c2b+ 1'b1 ;
assign I33cdaee4676d546dd5507df4704ea1f8 =  ~I6aa13ef29cf7e86ec83affca4fa11e42+ 1'b1 ;
assign Ia44daa9ddc3e4d377267333813d4675f =  ~Ide136b08f4b6211bca8cccf494a0baa5+ 1'b1 ;
assign Ie1f8fff3f43426d6bc39e45322a532ca =  ~Ieeab247764c23256749776b0a164314d+ 1'b1 ;
assign I4ee181895efc22862b6e85802a944095 =  ~I210e9ff7f4588185bd712915954543ce+ 1'b1 ;
assign I5c24ea83cabbb6be089ac084732cb9d6 =  ~I59186d5219833d6dd2e813a2910a61f5+ 1'b1 ;
assign Ifee2342449a3b3d0036ce2ecbc9ae189 =  ~I0c8b2bb61a9c3a67ac7e03e40be2b98e+ 1'b1 ;
assign I70a9a9b8f25066612a50e411ad68e6c4 =  ~Ide24c1f9033e7057262da1bc4762b840+ 1'b1 ;
assign I1870059af857c79d444bef948bb536ef =  ~I4677558b9faf190e7960cfa9b8ee00fd+ 1'b1 ;
assign Iafe61ab12e232a1090123a0f16eefaca =  ~Ie38ab94215851e531d2100b6602d5fa5+ 1'b1 ;
assign I10ca809fe9a04eaf5d7784ba69314178 =  ~I3f5119e8fac99376aa38e4765b8b0f99+ 1'b1 ;
assign I7a1bd0a115b3a1f85cb9c54840f5bf9b =  ~Ie8040301d224f78c1fd18bfe9e29e5ba+ 1'b1 ;
assign I986a564393d944d7d202414431c6d165 =  ~Ied989966cebf0d730633606c5182a249+ 1'b1 ;
assign I464042aaa60a41c7e1faf3d16eeb121d =  ~Ib8818bc4ca106ae38cacd5c20083aa08+ 1'b1 ;
assign I34b9a0bf2b6b562fb36291022ddf5179 =  ~Ibf08556fc39044222321912e84a4436b+ 1'b1 ;
assign I17dd8612b5c7f9dcc90f17e584aab2d3 =  ~I985e2740ac0f656da8f9dd973bca99e6+ 1'b1 ;
assign Id77cf7c05844d83e808a694971145261 =  ~I73012d2d9f6f237bc50bbffc199e012b+ 1'b1 ;
assign I276c1155d766437253f12b25066b84e4 =  ~Iefd0d59e58623b14437b17297fdbf4ff+ 1'b1 ;
assign Id75b386d8076893cb73baca69c3eff59 =  ~I68d2443e98f2fd3fa3baf96f98e1f4bc+ 1'b1 ;
assign If62ddbe87274965cfd83189c6666401e =  ~Ia2d1b6833cd8ed02f05281e508e4d716+ 1'b1 ;
assign I4f73a07452638a610b31e3ee52cb5639 =  ~I512e2251bef73108eb0f3e01e79ca3fb+ 1'b1 ;
assign I2a4faf3344d9bf4ee71da0be8994788a =  ~I9bf64811d14ca8b4c633342ad22669a3+ 1'b1 ;
assign I7d7ad0cbb962a47e229fe9d8406e6fe1 =  ~I45a910acd40d5b9417bdfdc50cddf241+ 1'b1 ;
assign I82988dc2dc83ac61380d2a5cb6551768 =  ~Ibbcf5c5f4528b03508b506c43e4511c4+ 1'b1 ;
assign I058c3a9848fd30010e4742d8682081ac =  ~I2b8b54048e164ef2f1c072517fdfe400+ 1'b1 ;
assign I368121c2534820a7147858c06e58b3fc =  ~Ia48d8883fe4f685477da6b4b05ecd387+ 1'b1 ;
assign I03d4541eeb1440aa72ee490c49977e32 =  ~I276395da1f3f1ae246b082408be2cb80+ 1'b1 ;
assign I75fdf5a355949a87b768b1e67db674e4 =  ~I4d0e2e01d9abf9ce839fe650abfaaddd+ 1'b1 ;
assign I088f4a0af0239602d422324549cb9799 =  ~I7e4e7909094f762c54137cbee99255e5+ 1'b1 ;
assign I787fe66b38237caf805ec14970d154c7 =  ~I761255e100d161b25645ca3a5187e82a+ 1'b1 ;
assign Icef176cff3ae503dbbe2af9ecfc4c859 =  ~Icc2ce1fa3cde69256378ec3f4a07b0fc+ 1'b1 ;
assign Ie0a66e4871bfe94f6716279ecc9ef21c =  ~Idd99afa80ca23644675d3edd60e74fe4+ 1'b1 ;
assign I474adf7a975b405c288058139a08be38 =  ~I486bcb4fb0af80c98c2ea21ac64f7a90+ 1'b1 ;
assign Iebeadb39658f41dcf8719ed413e46144 =  ~I759cca2c0003fc2c2af7709c5ebc59f7+ 1'b1 ;
assign Ie018b0d9f05a86207ae09ca2efac54e2 =  ~I1d5ce9f132cd1f46e96b511c77234e21+ 1'b1 ;
assign I51ee69807609fca0f332c8bc31afd632 =  ~I032e26ea05e88c6d325a810b67e82306+ 1'b1 ;
assign Iee1cb471704b2a8718a68ef93fd2e356 =  ~I0f72df5225a1fec2f276fd3c9138e8c3+ 1'b1 ;
assign I1731c0e3be86eec142c3732ee836e4d5 =  ~I0d18cf087b2335f1b9e1a621acd5379f+ 1'b1 ;
assign Id3b8c0ca32331f94fd98c8dae72bb15d =  ~I7684fc23c57105e856050a45640f2bfd+ 1'b1 ;
assign I6a86b0a82441c6c14436a3e0af6b0fb7 =  ~If778767ab80e59e940deeaa8a0dac99a+ 1'b1 ;
assign I8c92ff598084da7a50f7c68da96620b3 =  ~Idaf86833beb8c334f99291db9302ed29+ 1'b1 ;
assign I8bd1862e7bc2e83e9863389d532e6623 =  ~I6610e8d41cea10498d95850440ce388b+ 1'b1 ;
assign I8053269f8bd78a931878c8350693e1d6 =  ~Ibc653e701eb995e828c8180efaa122c9+ 1'b1 ;
assign I2ff66cdd7314276232715ef2361ad184 =  ~I21d36c49c9c766139b4b01df7c00a8f3+ 1'b1 ;
assign Icf541c76bfaf37fe6111de037d205f15 =  ~I0e4ffded936d7ccfc32b410aec617df8+ 1'b1 ;
assign I68319c8b9febef9f564832429c91b85a =  ~I1a5745021323efb5327d0b893962e852+ 1'b1 ;
assign I127772614218dd7c50d3136b4f174d7a =  ~I65547afdcd7fedb7b44bd51358eec4d2+ 1'b1 ;
assign Ib8d1aea4ad24c6ceb44f2cc672e1ff90 =  ~Iada3eb71e94ff6a6f4e5c702e83036ed+ 1'b1 ;
assign I9ca26c8104bf15f48b19dc3256914544 =  ~I077404a911da16d707a326f18717dc7a+ 1'b1 ;
assign Icc76d9ffc3f3d7b410205eeb8232a33b =  ~I6da1e92759c96aab8b9207a9acb244ab+ 1'b1 ;
assign I7fc4551d8a0445f79b87b4ba5f2ffeaa =  ~If7110182720ffa279b1cec1305cf9889+ 1'b1 ;
assign I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8 =  ~If0e20ea1696ff84329b9928d7f9e3381+ 1'b1 ;
assign Ie34c07af9f6adb9e4b636dce3d0682c0 =  ~I4e69ae6e73a856d4e26203fb9acf3565+ 1'b1 ;
assign Ib869a349250a765d2f8660e0dbdcf312 =  ~I64c939aa568669b4567c21be09ad0e94+ 1'b1 ;
assign I1a4fb631fdc7b5454c266589962ff5f0 =  ~Ia88eb16f68265e322509d541eb457993+ 1'b1 ;
assign I9de4e0e86e9edcf948d9eddf0401b94a =  ~I916f75e5a3858a420ab5cd4c43b13921+ 1'b1 ;
assign Iee7b4838986c962969c00a0bbe53ce0b =  ~Id076f99460a8f73a9fd43467216e8f8e+ 1'b1 ;
assign Id81b11a8ca1dd8989e36cef637ae6aab =  ~Ib4d7aeb8544fbdc36575a55b9f67f2dc+ 1'b1 ;
assign Ibe96deab015b799fe7f69bae8432952c =  ~If65d2514892fb7ee64fa4dc37fc0fed3+ 1'b1 ;
assign I986b52155cc1470299321a4933241ed7 =  ~Ibef07e48768252e9b41baf067bb1ff5d+ 1'b1 ;
assign I04be63a04f3942ce749cc9bd7540e055 =  ~Ib8fb61fa9cb8e92bc57c53a567891895+ 1'b1 ;
assign Ia7adea5b0ec86e9fcd427a5468d72b64 =  ~Id8f5f32cd0757b4d6861d17fcbd6e8d0+ 1'b1 ;
assign Ie8990d8abd23f8f9f79d7fe38c57fa8c =  ~I8be241f29e7eb258e9b3501430820b0d+ 1'b1 ;
assign I9d2f90ddddbdbb525d5f070f32546b64 =  ~Ica8a188ea43e2f28e70b8ea4e2431dc3+ 1'b1 ;
assign I905256d73bdb63bf860e15687350795f =  ~I83ceb726e57d52698b57dc39ce585897+ 1'b1 ;
assign I9adcfc18e4471209edbe9a379e996067 =  ~Ic88e7e05d83ff800b4a941ae4b424557+ 1'b1 ;
assign I3d7d048348bf833f744a9f73889b7802 =  ~I7de81aaac1e5776dfb60eed2d12d4f6d+ 1'b1 ;
assign Id619e8d4040014d0e415ff71c5e0591f =  ~I37058036bd9f4331387ee4a9348541e2+ 1'b1 ;
assign Iaf3de2ef283e03dd72002026e1299224 =  ~I570f85838c418d8501c8ccdc38a53f00+ 1'b1 ;
assign I64551529c0028ec145407be7f5dfef71 =  ~I4aa6f0c0f5163b944f11328888af73e0+ 1'b1 ;
assign I5ebe580a943b65fb16ea722ba101fd05 =  ~Ic7fc1f38ad4e9b2cb472ae75bc3c100c+ 1'b1 ;
assign I0921901599c43b27e701758026dd3ee1 =  ~Ibace8d2fba25834c83b1e57195c81086+ 1'b1 ;
assign I6033532f27c26b2d42bb3ea128f80dfa =  ~Iefc1488e3eb60b99ae08d904a15c5242+ 1'b1 ;




reg  [SUM_LEN-1:0]               Ieb085b219090cde5da2190093ce43730;
reg  [SUM_LEN-1:0]               Ib325dab091dfc3a1a269adb3ea9c75cd;
reg  [SUM_LEN-1:0]               Ifc045af19c3f10d92d2b0dfb4fbbde38;
reg  [SUM_LEN-1:0]               Ib79e305e6f44a4a6ebef1db5c70246ea;

localparam I0c5eab3e4dfde17a8c7261f7827e941c = 50;



assign I40a85f3ef46def30cd7707afd2c7fa44 = I5b177dd5c14ad082516b47f550875682;
assign I91679dfab57a372eddc7f9b94a231edb             = I18d11d94a39d5d7687736d266d3e1902;
assign Ib8963a4ab143aba7fadc61d89f937f4e = I477326720157df2503149125a43ee987;
assign Ic2171967791a0329f3e39fc19d0a6bc8             = I6b9ffa985ece553b83f7227e7a85141b;
assign I9565de7442acee8455d1c4f8ab43ab07 = I319012bc6fe93d78de57bcace0caaef5;
assign Ic7e35cf8d5cd230b94c40714f16e2418             = I49fdba80df1c667dd264e5105a530332;
assign I26b11eb80b9a1752998f7ab1379e4124 = I174b6c36f2af82f8047cc76543a3b4ee;
assign I679baea452c3c6d04c53baa88edd8eb3             = Ibf4fc04c9e0aa536a8e4b8a6192d8498;
assign Ibb068f313ff784191769e8da44f023e1 = I8fd5787ebf758919e7cb75d7419441e8;
assign I75a4cf2948bebc58e12bb039ed273ff2             = I899abb7dcba235ff2afb410a87e16973;
assign I2348d423bff186f1841ecaaf44f4f2c6 = I413b1c1985a6c9c6f202e85ff901e3a8;
assign I9d15f76bb68b214057566cba4b511214             = Iab322f0da75316ca9937802a327dd537;
assign I3b28138cac28625778c34d4bb1a4aa55 = Iea3e35ece9fdb3aff3b9ff5369e9a7e0;
assign I8be20605d26d218911e80a883a90d085             = Iba0a4530bce787d70253a92c123f589e;
assign I8928563d2510725797f96917767f9bae = I30c0fcd89e0cc7c5fa348df7b4fa2ccf;
assign I08a8cd6965c23af6650568b654831b20             = I4475d6a1e59d35444a6a2d9647c6761a;
assign I989726d5ee5f23a016e85b0945573f05 = I77b05a8aa92c66a235195a66dc13c0cc;
assign I065a81ba25962785215583e7ece27661             = I217e2e1eb3404ba9ff06d284a18256b6;
assign If88711683bd32856ce45937b841581e3 = I876fdba97e755b74532f7ab191fbac14;
assign I71228fe4188ab1d9796081184a422094             = I2003418e663144ee49f1ed044f6a0062;
assign I015cf78df7e3417d5296eb0ad3019674 = I5590d801fd7fb496019d4c31b7c6d898;
assign Ide9ef5a16d8fe32353c2c2a30e8ee3b0             = I4496255218b6d0f5374328803aeeb412;
assign I31908b38609b532f9f142a97e0442e55 = I25f1ee9cee4d04bd8fec1fe601d016d7;
assign I0865623d3350645e63fa6e6c9b78ac57             = Iecbb3f290db6dad3393b592ca946fa13;
assign Ib98eadb333ebca2f58c40b8f93d87250 = Ifebcf64858d5e2d07ad7894d6182eb11;
assign Ic10356f9069e3651b9c045c906e63512             = I9f88e23f2a17035b31840356a5d0bfde;
assign I4a0f0579aa9b7af7b516780074ca6560 = I163cf58b9a308e0439a8dc7c1526e6b5;
assign I43f41bf07836cee48069e9890c1de2a0             = I3fd4a13843fc09ca68b827a8b09e6c49;
assign Iaebca9b574d490aeab28fbbfb1e8fd9a = I3347717ba9556e69de30ce7533d4f5a4;
assign Ib8dfd9b8badef282ca00a4f793c3c868             = I1530e79da3803bb87787397f19822dbb;
assign I3ad613d80a126f03fb9125fe6da1bc8d = I5f96a68d20e3ebc71dad4b43305baa20;
assign I2fd872df07f50688486c0d602cfc5549             = I613821692bb99a8a6739d3c3ab7211ac;
assign Ic116b21b5744ec42a9f41eff3ddd1707 = Ie117f6ec475f5d6444998af151ce4e69;
assign Iceb7a1d4c23806b8f5824016779ad129             = I5ac600834d567934bd2f0b14a3c38ab9;
assign Id9f7e6885737ee2d3128081915a685b0 = Ia538dadbd6ae3711740595a18c89b65d;
assign I7b561638da1b4a45ff59be81243e4471             = I84fe1a1ecad408b16557957b01cc94b9;
assign Iad36872fbd9ac694d47cc0491f3d021e = I141cda06bae0c5666e3bc61c6fe5ad66;
assign Id50edc56fce48130247fdbc42eeff9ea             = I7d03cdddc264c89446cd80405c34d69a;
assign I0794dcad0f96cf58fda60c561a1144fe = Ifb70a30f8bade95f402e71f95fe6644b;
assign Id13c99b7f7500c8195b54627efbc4232             = I5cf7e3cb90e84c3ac6a66fb6dde220af;
assign I8b4cdd738b1ed431764d4a51be668460 = Ie50aca688b3433fad7565998cb900155;
assign Ia92d2276a8a23521ad1b88df7c27bc2e             = I602c2e5bfa93cb3c87af70dd69b0375d;
assign I79e67c70ee26ab7623355ec5042dcb28 = Ied33f18cbb778d5ba744d249f91c950b;
assign Ia96955d9c0a8a587e0afab37c8415d8c             = Id50fe525d660f0bb0ac3bbe6e68758f1;
assign Ie0a573c73ca9198012dc8ff4f8373973 = Ibe97860165dc5d9a076ebd935385ae51;
assign Ia9b5d9ede006c56a6d83905529c77b7b             = I6a68067b177340dbea2c53f7d8bd5f14;
assign I6a4cd5680e34df5ccfea4a7eb72113ec = Ie46b71f55aef4d00168202431d47dce0;
assign Ie9ab3c88ac62369e3d92d110165a94a8             = I9efdcdeee8883d30159881f8831a2c03;
assign I9885460698fe454e65fea4a6022e5df0 = I92cb615e2c439914e72ce001256518e4;
assign Iea07d1adf9016a29cffd61d183e268d0             = I46290d63552b8cac8d22358cb38c5887;
assign Iee7e507956faf7cd903ac2dd636b7819 = I7d6a6026eb3c4d06e682523424f9628f;
assign I37e6bc7aff363ed0ed1f84b23c5f3e34             = I6435c7b1b3bfc5dae42cb1b3b03aefc5;
assign Icece56258c1ffa7a0257d68ef9ff5ee7 = I06ad520cb02e46d34c45f207d42a9243;
assign I47f17afcd5871fc3ac378316fd3d7ae9             = I63b2f1c2148e595a40bb41968e4b9a65;
assign I6c15ea618986f2043f402959ac23fb1b = Ifa3df8b249467cc1e827c69925ef415f;
assign I57015930f5b09a6c6b030ed01dad2177             = Iafb6296c59c2dd241c880c6d57352617;
assign Ic45cade04982e60abe32a359999a778d = I4ba41864bb1d2130c6971e0b2903027a;
assign I26a7fe395eb583258c1ac58aaaa3234a             = I0b982beca6221db7b3ec2afb3833a60e;
assign I670dbb51097dde1f56eeb7e25ac50369 = Ia67f9b902a21de0414eb8dda52171991;
assign I15a1671def323cd294591564ae6ef8b1             = Iece8968796771c1ef094808823da8962;
assign Ia3fb4901b185e64ccb788dcc1d7cfb1b = Idbbf2ce4a30787c5f07c3b908a73da75;
assign Ifeaa99e03bda8ded058f98387de3d49d             = I05c7cb4a076239b8976a76d418ad6149;
assign I15a23e6922630f6d409706b1c4100d22 = I71d3a999d88e591e102398409b3adebf;
assign If520c1cd27f9d4bc52d0d029f693b660             = I9076162e7b10bffbc9473e35b407e986;
assign I08eb91ffc153d5007de61e2938407d18 = If7f3174da35dd39af7f4792aaa649bf1;
assign I40ef50004a60ae58aedc49eb5e6797c9             = If702042844ed38f5e7103382ef4263eb;
assign I642d63513e039da95a66c1cd4336f84f = I953b975a89adcc88039284970e9b3404;
assign If4132b39ddb92aa02d8d0346fb0e6691             = Ide63b2762649761944db237c8efe69ae;
assign I1e35f6f8ac9e61787a3b263e5e4ac62c = I5a247475beb737d470f03507e55f5b24;
assign If2af8106efc1f7dd02c074af68278b3d             = I1cec628c6d6e22895a0f0c0258851171;
assign I5af04bd644d9c14f56884acd1f6674a7 = I93084ccf5b5e4efaee968b497bb2a775;
assign If8a527cc7f06a9963a80a880d225d34c             = I46b0b74552e89df91c0027f0f093e1f5;
assign Ia9bc04087c3926bdf993858e683dc3f6 = Ibab55499323660588ec82ebd07ab0572;
assign Ic3a431f39c678b7175ed30fde1fa6424             = I68dbff67a1910346ddc0281b445f4439;
assign Ia8c23f2c6c80bc389fd66aee524975cf = If9285bf7611bcc5ea6432215c349e021;
assign I4af080cb4e5cc525db95e5f401019e8c             = Ia42f547c0b02c2de66f2ff383ca1741b;
assign I74ff51ab0824be97bf311b50b4ce5401 = I3566033cf5c9a06977c9182925750707;
assign Ic6386d7d8813731d612e24b715740275             = If456045711d535cea07d9dd5ef9b04c6;
assign I22cf21c1e88c0b8ff5d5b43835b1f61f = I87b10521099179c18652c86d5887c908;
assign Ic512effb493a06ece58a2af155135004             = I9585ff28ce0f3bca71d582b1cb8937d7;
assign I2fc87e59765765e16bae0761ab5741ec = I13a98f98c54b2e412cd88c96f016c41b;
assign I9b6a674dbcbfcf65f1ae0deb8fc3566d             = Iac3dfb28a343cbb391fdf58684e091ef;
assign I6c6297e7aca3c7d8a9f8c3542f8b070c = I6f7a45fe64ffeda9ed120be3a4519aea;
assign Ib4bdc9069d0c08655f5e87f705943eda             = I82650d4bf0a9b51e245665259f40fe60;
assign Ifbc2ba75815cb3aece1d327a5c15dba4 = Iad799775eb657f8973e6dfcf70a9875c;
assign If92db65b39a83e1c699e4cc6d7f9e57b             = Ib21e67aa9696222891a0b33c414b1bbd;
assign Ib1bba2d65c2224f05a444c6170aba187 = I5ec1e530b9007a75a778af4d82ab427b;
assign I0262b30a4efa9f1cfb11d1c3940de9e7             = I1e168bf1a0dd18ff31d3560be00095f1;
assign Id75ce45a6df04b3d173b288b52d82138 = Idd59a5357d4c835379ed180ac0924bf1;
assign Ie8df350430970b5f1229cda772440f85             = I97e6d2bc8c1ad455f7c61de81e8d4826;
assign Icd148cb7a25bc30aafd0271e00356527 = I7a626ec321bf963a5401892a7e3891c7;
assign I8070a3b7d8b1a7ae90c1a2d27aed09aa             = Ie1170db51d408ccc7360ce53c94a9644;
assign I80e8b0fdd6bfadac9c8a788bd9be4b97 = I3342fe0c5d3ee5021892d53eb45bde21;
assign I39bbec42c442d1e8c818f46ad9c096a8             = If58c2c1e1dffe04295f3313595ffe319;
assign I471dd2bc897a40a9463f4984952d4fa6 = Ia858ff5551286beffd4cf82f876d30ac;
assign I9bb81dda8102b829441be46460eb8900             = I9a9fb4da9fdf5bd42cef32c7d8fa65d9;
assign Ic61bade7088606659ef8568dc134f686 = I5402fd208dc7ca81dfd2920a9cfa2715;
assign Ib23edc35fa5bbfe0415fcf0861a22d9b             = I785e4a1f2556289db0bd024e429bbd3e;
assign I298e98803772a458fbeed1de632c0555 = Ic32c6734132776c290155a80025fe366;
assign I9cc16a00912e7dfc05fb505a9db23cd8             = Ib6ca0cbcbaadb956d19a482fc099b175;
assign I605674982abba50698d4d3c2220b0db8 = I5d92fdff96b9cd64f3af2b28b13e9956;
assign Iccefa45795486757515d95e5908b306a             = Id52b94ae6662bb2137d8b9d53280bcdd;
assign I201d44bd3cdf2b34fd2564188190b27b = I221524a69e18854f029cad30e8f94e8a;
assign Ic3a608b850709286ea0ad2f67425d9ac             = Ic3975e4171d618ba53e1569e4fc93440;
assign Ia764576ce7e8ec4fc7120bcb8c038422 = I55e4ad2d71a29ad63b4999d64ac0dc4f;
assign I2213c1a2b831f421707a261f5a58b1b1             = Ib4e0f05afd881adf14a5eab850c75a3b;
assign I66d5eccef31484a090c91507a3d38a85 = I592a495aecc800236c3470ff8e6adbb5;
assign I4636821315d702a677dc93113872e647             = Ifb875d675aa28de930d889ae4d37b48e;
assign I93cee05370c836746d1ddeb0f74456bb = Ifdb5589982db805a0416e1c01276249a;
assign Iaf8a19fde3de660c3fa925593bebbe0c             = If98948e5f60b2c3ba1d7338e24dc0df6;
assign Iaa19be06695f47ff7d10667289dbde36 = I0c47ccef4b55410286248884a7249703;
assign I0052d562fb3182890c8828e52d437b11             = I732bb69d248d700bcfdb287932839da8;
assign I21adefc729265cc5ae67ce279a0a78a2 = Ib68deeb7bec4ca3585d1a4dcbf8793f1;
assign I21668ff77cf75570cae97f575cbcf644             = I403a8ece76036b3ce6277435609548a5;
assign Ibc0592b70bd60e475066554f0c7c4171 = Ia17906696bd0e095d7a5297da2e049ea;
assign Ic279867ebf3055980f3d813d5dc8dec6             = I5a6cf1bdbcb2a342e548fb44c171aaf4;
assign I14f80574ea80b02ce13079854991febd = Ic11a6b77b84c44180eb99220a0c4c9f6;
assign Ifc8c6df8904b97674f2970ebc95b523c             = I83a16a5be8d92896234bb9f2a36a22c9;
assign I09aae1dd6d02bd2a65dc7fa06fd848ca = Ie08ad9bd71329858c1742c8f571a1c36;
assign Id88480a0a350bb5fcf01ed5fff0bbd4c             = I6cad1cb66561eb6f0e3bfe5070b290c2;
assign Idd698fb3a64825b43803642fc91bf674 = I8c0c1a0a35f4f7a688f516c567242d39;
assign If38feb4f76f761dce6145731ad235d7f             = Ia50c447d5838d7979b2e19796be6221b;
assign I73c9bd7e52f6049b733b3a594ad6fae7 = Ib105151d91678f81978495ff94b1e651;
assign Ieb528d666fdb708279184bb59eac25d9             = Ief62ab0263b74086ae23a208da23e9c7;
assign I0fa2b3408156b2b0f656db4947670fe3 = Ie92110d19f4886cdfcfacd0920c06a4e;
assign I631a3300cb6685f47da7781940ec5d27             = I564999dcc2f67c8f82fb5cd16af0ee12;
assign Ifd85deef561f76562208a8798b540b99 = Icf3ad912aaeaa0c5cd1ab0edb898d6e8;
assign Ib54d55a70605119e37e9898b940ff636             = Ifb0e4775ffb73bb2533844db969ab900;
assign I9d6eec32202aeaf66e7815492ac483b2 = I857d3155df0b6dd704514b039c66fa97;
assign I49fb0909ddf66fc0073e6400f1a07844             = Ib109fcaa55c3094cadb0c1f5f40ca752;
assign Id771356ebafcbb0e2bb8b03e49148b99 = I3bc094d67805664859fdcb66f1360e64;
assign Id0eef1adba01447c14a6f005782dd9a2             = I56aeb1bd0b0e9857d9cfd2c6b347fe91;
assign I7f4f192560919410f2526392d10776a1 = Id14074d5230885c38b89b09b130ecf68;
assign I5a9fdec7d7ff99fe33ad6cd8afd9e059             = I02651642fc35059fe9b4141c2fa1f34a;
assign I4e2247be1d2dd1af7467039a05447631 = Ibf312ae4f51fbc44b43848f9df62a45f;
assign I68528be9951f5b8805411711cd11ea59             = I1f1e04979c8a5badc8a103809f76dadb;
assign I5146e2d888c120b7afc430cc8d1dd34c = If6ce2fa9f0b8bc74442ed8262b5089cf;
assign Ia3450e134e4086c35acbdee1e6042396             = I19fe22e1104703ddc9bbc94a5368bbc2;
assign Ib34be78c56c66ff7d85745612cd59f60 = Ibabf61085ca7af8dfc7927b3656a76f7;
assign Ifec374bce7f5507438f550df22d61a01             = I4386a95203c4fe83c6db7e25a288fc4c;
assign Ic6f48b24e0247c43666af5f25f03c1dc = Iebecd2d19f9174d87deedc1a273e7baa;
assign Ie87075ac979410cc11099a356966b8a2             = I2ddabc0b4bc45698fdd877c93bcbe280;
assign If9f312c27d80be62969c60eb9b67586c = I94a9de743d5bedbea3876de954f479bd;
assign If4d3b31b87c0f723241d35ce7e854eba             = I5adddbf99d0d39c5d70ec6a0978f3ef5;
assign Ic7e3298aeb02d5829de1904288687002 = I59c5da6338f431a626c86a065a355c35;
assign Ic53b875b2ddcba11406eb2ca39354757             = Ia24d776498719aa6cfbdb5df69d648e3;
assign Ib45f271c90e7bb32cba9dbaad5334c67 = I8edf1a08ef943f06ee28771c6e140e28;
assign Ie19b39200436b0bfca13502ad36c21b9             = I038ff8eadf1c551dc42d09fbadaea5b9;
assign I727821089976c74cd540ec58ecce2da2 = I1c8024aa9d81704d2dcf63e34853f8cf;
assign I9c981b0614a29386ca5e8ebc06a17f15             = I102dc8709a274d21c09abae1d2ac1272;
assign I4ed27d0c804891ee239ae8259d200712 = Idc1b8aa2f81a7fbd87e4f5821d14bf01;
assign I9938397dc94002481984f5b560fadc58             = I136256458e71d84e850b61a950f279e7;
assign I421ad50f600133f1e7f6a52625181d36 = I02812a8a833bb69eb168a1004b6fafdf;
assign I4c366a57920ff090a98a2cb8b9caa00b             = Icda6fe755f2d840f8e404d84b231e827;
assign I172379505892287217e08c060285018b = Ic44eab478be232721e7a43d14beca32f;
assign Ieafa9d74d4a61d28ac4a913db460bf33             = I1f6cd53f31f27d86d78d5079e84c9716;
assign I8ac36cb7b4e56689efd4a3de1fafa0cc = Id1dafb7e45b860d506e0c2c91b28142e;
assign Idbf9094c94c931f16fba468b9dd59a25             = Ia1f69042d447cb17772b29f634344b53;
assign I002e83f2fb7e5b07710a802aa505b2bc = I9db50007841762c9a10f6b7e9d40f858;
assign I8d8d95ff26f33f69a182b32ccde23905             = I84648f139f0fd470a62f0638aeee9e97;
assign I26fe780ca6becdc9f86a7be04c6257d2 = I36ba87b69b5b9dd919319230f697dfad;
assign I8bbe1a2ace8f51aa22cca5d9fc66f136             = I6ebc0ad14d76d3a80a4929ba8b5e7848;
assign I3a8d18e570ec3aefcdc29d7bc783dfde = Ie7d9730b191781c78391141d95d4f8bd;
assign If0a3b88a66a816b25f17ced5d0e8f775             = I26cba2d4920ff7fc40b1723c29ed8391;
assign I4ddf83c90adcc1bec65f265e898568fd = Ib774f380e3d7cfd1f5f064e93d8134b4;
assign If7e146da4f3bd255b8457fd6902005f6             = I27980b3a1936a92a1751588f91a5f542;
assign I0c06a37e120e59f19578c68801a4b6ec = I13b0c9578f7b6b3b7e6704d7b44079c4;
assign I89a3f8d5f760d1a650f85814cbfdc017             = I5464cf638e0ca778d4e113b216084180;
assign Ic290ad8aeb51c16106f9311b06134a2d = Ia01c82761aeb124cd92fb15ee367ee8b;
assign I3e0e682047f7cc36142e668828cbff1e             = I1804dfc05236c728f563342eb011f4f8;
assign Ic4c7c898ca601e4d44076ec5bb475979 = I2db290170ddae8dc52ce07edaf48b365;
assign I596ad7e132f272cb196b74faa8c75aa4             = Id219264de5f6b67cff866b2bafc660b5;
assign I380cd867541300f76fc359d72f49bdbc = Ied764ee7730ad129b6f62837ef50774a;
assign I5267fa34449e6eebe891017fc32d0749             = I03e4f803d4b82aa774662e02b188b0a6;
assign I350f20848080cffa45a31e2f1e553a3a = Idc5dd6caa4ed17a63746d30d381a944e;
assign I2dc64c3b06588542b027f997437bee63             = I32e079707d9ce4b31aea8fd2c998c27c;
assign I912b9be8432d4eb792d79566a8280703 = I719a892ad54e63b217c7271741b29cc5;
assign I753f92da60980736440aba814a156f1e             = I488f60405ded7af04c941bdbf55290f8;
assign Ifaed59e29ee3ee9166192bbbf04bc682 = Ia0c192e590d8c914555b434ce5a634a8;
assign I733605337bf6972630c089d32fd7f98f             = I26d314b69785bdb0ca8cd52c258c3b35;
assign I7eaa9f70586b12e371db5964758ee7c2 = If2b40d249c531e10cc22d1335f350441;
assign Iba70e737d52e6812a67c159520e5192f             = Ia490437ab050e63e611dfb4d9366017c;
assign I9a8946bbda4bfe72fab3c2f59533b3ae = Ibe7e5c2cb9c50eca34a3859d13e83a92;
assign I7d77ac9b64b2e8cae21c6e36947e3ca2             = Ia6cc50c8b7f83dd80d7058eea40338e9;
assign I29fd8dea7c3c39722614210cb7f65851 = If0970d9f7b053fce3ced3521b4885588;
assign Icd0622a90782b9c451950e7ab0399567             = I3652208cee3ca6dcdef63b7df53e4329;
assign I54bed2059ffd24ac2fa91b038c0256ae = I777ee54ff20d0544af18ad8a870d6915;
assign I1487170cb1f3370ad45efc801cefc8ab             = Ia9a4760f6a2bf8f8f660e2b0c31dd823;
assign Ic3608e6a6c45ee04ccd8198c88c69003 = I4edd64d1f1da865b1eb886e22726a033;
assign Ic3ff7ce12c836bf0693252b9a7a7cfe8             = I5ec267a535ad08c629940d70c61894a5;
assign I37da881d3575c055944719409ddb66f1 = I4dbabfd592b74aef93b819163130ef5e;
assign Ib23d889edb5a6d9f27de977d3b1a2616             = I17fadd913ac1008fcbefff48ad366d8f;
assign I2b6999fd13f9e57ea33c0b4602594c66 = Ifb064c69c7110c014593149ae69c75fb;
assign I8f2986bc015fcc64ac5e5395ac6dd851             = I275728fecbd15ba77f57860bb329da16;
assign Idee62819bc831a9ba7c73dea46f3da9a = I2c741a5fed7d88e9bdd6b7459feac649;
assign I7d5041a6796c00188f74936d283defe6             = I8d0bc446761559f2188e78200eb0a895;
assign I48c95e9ee4d7dd54b6bf21a9a5b20635 = I8a9e516aa824260998d10db758642bb0;
assign I7a2e79d42779ad235bca6ce3757cf588             = If9fc4683c2f0545e1f077541fd25da66;
assign I26b2a20b53a3ef8531d6798c4b272422 = I8bb5522183b65583fda83067990b3e94;
assign Icd1da43a4d95230e79dbd35a7ae41066             = I1c8e7559160d5a1fe1fa0002cc414d1c;
assign Ib814d21cc76c4f3135a4aa813dcb748d = Ib0001d7298ad1f3b1c7603173a70d8b5;
assign I5a0f27df5158309f32f0df31e8ae3ae3             = I059014ede8b9092d817c0aaa1c7ed388;
assign I44dcb4df87d1cf32ee2c9bea836223ea = Ibc9a860879ccc58c815b9f6caa23320a;
assign I4255ac1af4367c321567c4e46b06ab25             = I6294fc2c9181871210e0cfbb9834c3c7;
assign I96ea91e1bf398f6b2973e815a6a10aaa = I17c9d8f658dd6b2916b645d103f4702a;
assign I72369dedfe36cb22269033cc305b730c             = Id24dd0ede5504678fbd809ffbacd0dcb;
assign I75458b8dd7bf267526c36af5cbfcaad1 = Iba283e99a57d0a3b78ad2e309c316b65;
assign Ie65a0634454381e24bb3223a333e3ad0             = I496994e784eb114337ac9e78ec0c4d3f;
assign I230ed2d0ad383ba3a6b5b69ce09ab4b6 = Ic98c8641d2022080297c54ff2539e75d;
assign Idcb1d8bbdeaed6768c2a418c3048e6ee             = I44c28351f261765c28a066a581c27c13;
assign I6c09d773366bca735c15703f7c2c5a11 = Ia9c273b32d0701c7f185ab2de9e57829;
assign If3e5161254eb9056914c46263b865c10             = I84419e016619a3a33224eeaba85e68b3;
assign I146e4737d01377560ffeb78fce84973d = Ibf5c141c5cc0a6a20c05b52bf8282476;
assign Ic1faed76fca5a9ceb7db26c2f43623d9             = I67d114d975d5d65f575bbb8c819fa22b;
assign Iaa4c0cb6fd4dcc74d6ffd2bde42b7947 = I2518ccf385b3b677d95983bc550282e8;
assign I1d1a7c5928982c278d068ebd262254da             = I6a452adc2501774b55e5fe73c642ea26;
assign I49d021b0957d65a6c2608de826c2676e = I86fefad34d3c864dd0e725133f303b4f;
assign I47b1695a74e4d27389b97543415dcc67             = I33792929f4428ddf0629231288e459ec;
assign I72393e4bfc85c2b9ee24a4395b3568eb = I180d4f3b23b518271d7cb8189fbeadc5;
assign I5c05da8a222ad5effb9815cbf3ec25f3             = Id0013f18ab77416e08d994c360b13473;
assign Ic9f855b66d25668256912f2e434b4854 = Ic7ebdc317c978eb275eca41d5b9106a5;
assign I6493b3c087d4685a6b3f98c73dc2ff49             = I5683f67c7d462c01c55b8be9b6d1fca6;
assign I27fe4e83261eb6a1789a8f7d77a0caf1 = I84057a3b319ab3d6a2ed8f2310f970fc;
assign I2c72248cbe49ec0a0febac2437b8a6dc             = I4a5e3cf3066a4c2f7f5f8dbe824ff88f;
assign I45c158cf7145668cb8524f7fa06f9302 = Ifab075b1437495268b6a3be4cb022e71;
assign I6fd1b4395af175eff85b3bfeef4c329b             = I93879adfa4333a80be696d846e34d799;
assign I16d2a9270452f0d8b6eda06ea939fc6a = I89c5af1a6176cefa1f77ee69996473cb;
assign I2508854bcbab37bd09c9465c377c06aa             = I199e944b303446e2cdafb6f34d0d12c7;
assign I1ab974ad9718ea8350d76bbc1510d2d1 = I17a6511072c7fb4846be5844decf17d6;
assign Iba7608ee0a01af103e022bcaf564bf6b             = I91d282de42df72b1c439fede384d6336;
assign I31467f39d6b5c20d4e155d19afa34e95 = I9d18ff3465afd8cae63abba68487542e;
assign Ia9642d79bb50567348083b4435c7d66d             = I8a06d2c278af9d552fa36a61128b8a9b;
assign Ia8762fb956b52535ad6921e9191288d0 = I1e77fe6aeaba852aba34ed37dd53add6;
assign Ice9079fb6e08d629f8c0c9ce332c8f11             = I5a36e45af7599ec00703dfc81f9d1176;
assign Ia018c4c165c5af9a329a63aa365ac038 = Id38852415486e6989b89a0d85ad6771b;
assign I39ff4663007dbc89b403f3b08a69bb6c             = Iae09429ca8733186fdb3c50f36895746;
assign Id85085de57a0152aad8cf5e27a195052 = I89af7644c48a80d7d22f50b008d35841;
assign Ib01cfd833a63500e03333f263805db3d             = Ie5f74b33d06ddb8b32b57c8c82392001;
assign I461b443279e5bf47de450846e3da7d8e = Icfc03646b36b971b9fa57d04a26dbfc4;
assign I0f034a8f077b0ab231727b6298e366d8             = I7d3cdb71cdab3a85122130207d872476;
assign I71d07a22b66aed8c24fe4dd203869fa1 = I05e739fc87e962848f265e2c73338cac;
assign I17d9e19854cef197fd3267618617efc3             = I68ae9f2a14b161c940f6685073eca97e;
assign I173b85306dc75e596cfe67f7c518f36b = I624958486d181501c7a8ec2642cb503c;
assign Iacf9640cbf486411d6ceb8fe1a2fd5c9             = I778f907b5eacdfac02b0bc4547af4ea3;
assign Id57948138d3091aa350db0d906b06b34 = Idd775d9fe6fa8dbdbfb07d4071b9caa5;
assign Idc629414f6d0236ce0714cfaae23f065             = Ibcea5bf1e21fa764ac9f2d2702c8f79a;
assign If6b37dd338e28ffd7fb888bc56f716d1 = I17086dc5193aa55e5c6f56ecd365cc00;
assign Id92a37c091100e9df08e24498ecb4022             = I93a3e1a8e414d4775f19c0c9f16d07a8;
assign Idd412a66c4a434eaaf337b6b4ab6b0a5 = I7e12ad8a8ef857e02f4563b2f3a7f0ca;
assign If6657f90c84ca5e2ba08ec705f34be03             = I8772034840834e51187950d320f9eb40;
assign I5829341b8f12f906ffc53c9d716e6556 = Ibb35bace971548c9fc98d773d1aff712;
assign Ic51bb9184dfd103703cd0c6ad6edff4b             = I3d0aa00b61d4684ad46f49329197c901;
assign I449b6fdea575e92fa4603f141ff359e8 = I68b585571699a57bc6ba5e8955467119;
assign I4378d139db4b710e3587aa72df22b70d             = I146866a6d46604c47d87afa3c88308c6;
assign Ic6581fe8d97a45b71a1ca8d9ec97f97b = If76f04fe0baf171d7df2c0cd849aea2b;
assign Ie88285ce2b9c71de02ebd62e8f44ca72             = I84cf7aa78617faed2f1762bb1961cc0e;
assign I4af6879c6d4d2b96562b1c2ada8f92b0 = I5134b762ac428bed07ce102d8927a418;
assign I88f1b5c12759a5efb2d2ded8483c9ed2             = Ib1f43a0b9c86d236b2ed71c35c296b9c;
assign I7a176a15ab2c5396639be387bc43896c = Id277f5f05551eeb5dec1701056330da1;
assign I6fc8044eb226a14ff1a786ddc96d2414             = I88aaa7538f9007ce204319ec639d1c7e;
assign I38c29f53b042f039a908cca7d09cc2bf = Ie886c5effc85f1fe0b6411db4a2cde77;
assign I14cf5d43fc9864820a8a25efcc5c6d86             = Ie3a171564602e9936d7960e83bb0fb3a;
assign I1e5c60072bcfdc56b1928040edf9ecb2 = I3c10d579f80bd0106506ad047d75f188;
assign I1d9b9ff357667a362f0442f19986f451             = I732b452fd9521b3a13ff1f965c443325;
assign I03998667df412d12539d57112b6b6f76 = Id18c5a1d4eaa73a94e699e5f9e3c3d35;
assign Id88568dd34fbee42c9cb8cc15ac5c31d             = I16cd75fd747b600e90763d8ce9c08210;
assign I2ae5c6ae2de0db31a656018e19d086b9 = I9ece87047aec25abc02a5eea72f0e647;
assign Ifaff9dd032cf96487be819c59b03000a             = Ic6a7d6bfb12f40ae8823db716cfe017a;
assign I1e27f59e10400144106861daca51e721 = I12f2f886517647044cc251861721bbb9;
assign I0374ada4fe50717f2158468b7ad205d4             = Iea38a3c260d0caae4ae042264a0f4787;
assign Iba8577f8233fe013584171e588868e69 = I27e1d2e0e980216b27b90ea48c061025;
assign Iee6f2484a381bd42e441ff072ec582e4             = Id6240152bd22a9655b18bdfd91812e03;
assign I1d0a95c7cced8ede694d02936af63047 = I41eff06fe1dea8be4613945de596d3ca;
assign Ifae345c79662c3df3dff0fe68ad68746             = I07eeb34c9dfb9baadb9f263b6f095ecc;
assign I8b072ed41d990e6afa6fb5d22990f4df = I94e4041b482064334fd0ed92b91bde89;
assign I1eedecb1d8ff505c75be7787199afada             = Iedb57db3cbaca9f9a469d91ed81466a8;
assign Iab0f19858a1a01fe09fa3c99d92a79fb = Ida3d808d100e0bba290f96ed9e744e65;
assign Ie48be9e6b6fd63baa104d0a6a4561a1a             = I2972b771a4e99ddfa2178349a805b16f;
assign Id88441b410f55c15465eff4cfa216691 = I4c66570630a650fa7b9bec543f685487;
assign I8eef6ca0a61a21882ea28b3d63735228             = I6a61cdadaf987763080e6ce4d1605ee6;
assign I894540936535dd20ff1ea5c47546e5fe = Ib1a40247057324b0bd810c844bf11f51;
assign I99fb9030e8361e57818c07511479a9b8             = I12e430f1ccaa6099ba9ff803c85d9532;
assign Ibb40a1e09cc59e00ce8ba1460e0712d4 = Iddc5b5b4501f9f13bcaf22081e5a70f4;
assign Ief67e897e57b96e2ec200e82bbc7caeb             = I2cc3c84149c81572357c01219248aa3b;
assign I5349c1efb5233e8cc6c472ecae80ccc3 = Ia71cf07b645c58cffe33be1a9a960eb2;
assign Ia445bdc7def7d8c1eec31ab892c25c41             = I6d4b18dbba5c2b058f93a8d46bed38ec;
assign Id90c5bcfdae1c4abdfa194477917dfbb = Ifba3e46933049cb093d2c1809f3a8a3e;
assign Iad166146f7df5e8068fc6efe4d3e4141             = I32ca5d01c39fe736d6ed57d70fcbd555;
assign I1dafa9e7b2a353dee90a0b0f9685a826 = I4acf6d84471cd237f65c9b2391b7a20c;
assign I4ac79b67a8904b95f7912d24af420585             = I8807f2f633d64cb064fbc149ebd30412;
assign Ia75e6368415ff53bdbfe81ac2bdfb290 = I17b3a9df6752da6cc987e902e6bbad48;
assign I60ec7459bbe99fce295406bee1f2af46             = I822d3b3516499e58ee7777b99259a206;
assign I91217ca822fb03fdad03b8d005edadc9 = I168afc1863f909dbcb6a9230db9f3e00;
assign I6fab46b1766878b26b53f352fee98223             = Ie706bf8dd49322fc1d5d83e40fb20f04;
assign Iccc6e66d1f26c4a5874ba02980dad6a7 = I989dda9add29306d7b3c0f376822763a;
assign I36ca732e811d67cd742d24fd4cae887b             = I9975f2ca851119d7ec85cfdefda150f0;
assign I15e9479f1c9aae3c1f12f0f301ee275b = I7f7b30f2acbb8e31f50b58096b738254;
assign I355725a804e0df68b4acf96ca98f2448             = I2e0639bf4e48a7b1486beebcc9ad7c0c;
assign I14692ccb24148a020dda28c6f61e3611 = I615053b36a1851a06125e2ed5ec7f880;
assign I357137b41bb91e0659b1ac6ead9b5c12             = I6131789039de7dc431c3b9b59ecb7654;
assign Id237c89ded30e926343fb68d786a76d0 = I9890f7fc708c7b8cf460849b4a30025b;
assign Ie3a336de822ac7baf8486b1618ef1126             = Ia20482fd064712397fe2f9f77f4d854b;
assign Ib56bd244f7a9876fab3d51a21ef163c7 = Ibc929201e2eeb3e61cc8f0acbade497a;
assign I354fdd241d5d07f0d8380fe8924e0a8c             = If052875ec5a78a68428a1ff09df623df;
assign Ic1db9806badd4e959a0f0a769e15b6c0 = Ia098bbeda8b755ece6b88eac83d03e55;
assign I634484f00590216c0f74f975c9c83400             = I2e27abc9297a3fa647f50859af7cb094;
assign I3649823bb60a4740b6a7f94dd26e45a1 = I87f34821cd0b58f8855b25c75f2dd32d;
assign Ia89da2f1890524ad3519ab403dd0686c             = I5d5e3b64ed1ca16d65d8eadb8100fa06;
assign I8d7596d25b93595ffa1ef7d273c98c14 = Iab2f643f81921ed8464e1bbd9fa8c68e;
assign Ib1357cb20f471f1670ac2448f964f8eb             = Ie91a08b49b9bf23270dd3fa331e64968;
assign If607fe1cc3901fc74590a81a26ccb4a8 = Ib0dfbbbca2d3d264065f73b4241caed5;
assign Id38b705f5d2863a020a475ffffc8afd6             = Ib599712a1e8fadbdf7e3712bca6c0b74;
assign Ibe2cd0729747659786b76f044f3caa6e = Id20e72ac258d1d1b6cdca1e6c9e3596d;
assign I38c3e3e136acb79c8a0ff850bcc55f16             = I1791c009b0838ef10233015f80a5c4af;
assign I38e96074261512c31ebd15c6de4b440b = I5ebc3047985651f4b9a957d502a97e95;
assign Iedbe9d0e48bd36064f59faea51afddb9             = I3dead2d8d18ea8503a578469625f3aa3;
assign Ie72e9c0aa298ff1809a47908ff86b6c4 = I53222c82827cab7c770e057ae91bc10e;
assign I6359856a1843d8c8b65dc478bccb3acd             = I2fc47140b9df2544d7ae9c82cd38ebd6;
assign Id6e349e3f114f328958052a680a95411 = I339786aa60d4c71d12c65db27ac420fe;
assign Id6e5d67e7bb7c4b999459374ea80459a             = Ice09150d69c67cd2d08d6e63b8a9bbc7;
assign I6dff6c5c76c92ba9626512b35a573ac8 = I7a387a1f887c32e9d0f8e89912a8618c;
assign Iad44c932cfa5c249c5e59f8c706173a8             = Id67765c4a6b11f6ee0a4524ebb2d1ca7;
assign I5145ca1a0b7eb68adb93316264ed0084 = Ifa09fc1b009d073d5a9973b430c63469;
assign Ic3871325d57b310c95ca02fcaca529eb             = Ia17bbf4b7f063de0bf0701276b7b0c20;
assign Icff67cd5e9472e77380eb812deb625b6 = Ia9c8cc5e3becf3d48feedec8fa2c93a4;
assign Ica1997c6c569c1d1f45224fbaa4e6b59             = I9f9075a7745d475331f0b25bad830421;
assign I88adcddd217c9b2363fe254b0be469e2 = I4f134c0669b5a6a8c7e03be7eee30c6c;
assign If9c12f8662333fb54a45cfa1bc5da487             = I4d832ef88af4d4244516b0bdfd2b461c;
assign If149258ed84a848bc38011bef172b6ea = I1c4b29e48d0effac4839037ae5688334;
assign Ieaf14683f40374c4531326d228cb43c3             = Ib2038174dd555b1d058778fa904aee65;
assign Ie70f8bcc335351e60eecd70b90d4432c = I3ade020bbdf8f954821f737439513043;
assign I05341013abd4206eb66fcddfd63bfe26             = I959dff5d57b4c2adb85c3602d5874c90;
assign I5277100478097db96b41fe0988046442 = Iefe4099ff7e457f6b9fefc83e176c1a0;
assign I78212ae965ab2dcb2eed0b060d6b253f             = I30dd112c5a6793cf37bfaaf8dfdebcaf;
assign I0aced2534542d8d2c488c7082ca214ca = I487496233a32f657171b3789590d0522;
assign I29ab844f80c105d247c5c15faa35863c             = I4d4a0930420b4d7da8b6e91b2b25bc51;
assign Ifad6157e5199a5b5dbd2465f4cae5b3a = I39d3bce4060032a81e6b6a1c1805cfe8;
assign I7ef544597a185b1de63b4ffc4a1d44c2             = I7ae1d318fd0df386e0c8bcf0f0a94e4b;
assign I2bf55a177a00da61ccd463a450de2bb0 = I9963d0b24763ed8038b1f3922b8f9548;
assign I27fd0073dbcdee599fbe85cf48806efc             = I06cc62e12d5a261d672b5428dbc9767b;
assign I521e3e69d81a6034183d2ba861ec7726 = I5e69e930a318dcb0594a823b3129d650;
assign I5fc3c26d6c5aa893dfd5caa0f677233a             = I9798b16b4658501d739d46182d7ab169;
assign Ife32264cdbf7445987f5f39d6361d1e4 = Ia50526cd3a3174bebc5a7a0889fda661;
assign I15da71a21f5842cb65b543d9bc3e267b             = I90bc85b7a6e56250bf13407ddd32bf11;
assign Ied102cd26c4fc50aa354b16a35d3490b = Ie7470dd75b54d14038de19e4d3043ba9;
assign Ib3b1db2d8b669988c887ed780e439b26             = I88990d32bd34da606660f1c078b36ce0;
assign I5900a9bf6a83b1965f0dd9749d90e317 = Ifbc6aa14cd448bbe416897a3671ba857;
assign I5d70bc64cf7b3d3ef4180e082e533237             = Ib32ce57f2840a45fce8e66f71b37719d;
assign I1b4d2bc08a78865fb281a44e84088fa5 = I7547c56b32513ad45d775b4502596d9d;
assign I6354a0e638340378124e4df7f3d145b8             = Ib0179c2048d6c9d1865d171b48c521ff;
assign I70724327149d97d4d4f3f71a1500427e = If10f33385e236eaba56cbab8c2883399;
assign I438522d92cce6f7010246424746ca255             = Icc8ffcc0641f0f9405590338e6b5e517;
assign If91997f00102c66a7630ffb2d041d949 = I17d7f36fdade16dbcf621fe302bd7e57;
assign Iab953a8974a1eb619dc0f074c003b5f9             = I5d6cb688ef094e1f119d8536f0f56766;
assign I25da82603d45fc12f685407e8dc2f6f1 = Ie9f37dba0791359bc426a73639ce33ad;
assign Iccf255fb3422c558465e45226068a16d             = Ia5aa7c66d2818982a661e4d048876d1c;
assign Id2fdc5b6c996c567743aaf021a5e6371 = Ifc34f5d6b7a7d0533439794958959856;
assign I35b2c7e9cdc53a98913e1c16a3a47b37             = I449e514b6afb3e8e337691fc64f7431c;
assign I8d57ad30940b8351a829b8ca99921a10 = I87211ac14d832ad3205d47fb83cf256a;
assign Ie33a780b0221084898c9fc5b237b244a             = Ibbd5f0906646560a903abcf6848ee80e;
assign I2ccb382adcd7799634c86273c8a39199 = I17cf58ef5326978c62c03c56090a299f;
assign I9590eb28a81c730b83b92ef7653e71a1             = Iee607ab8132caf0f678324d20394f533;
assign Ie521ecd231d7bfedc8de182c5050f6de = Id79636d195efff260c430978f0bcee9c;
assign Ib8bf21f32c0e8b9cfa42a53807bfe3a3             = Icc90fd3c992755ac7e4aec1370600e06;
assign I855892c34f1706745dda4ffc3e5e5a98 = I8015717cd36aabbf2cf4aa3a5c234690;
assign If6f3d91c3c7a43622b9a522492cd83d3             = I81e0ea92e07ed7d29b4ab769443b55d3;
assign Ib945fab3df6e5a7494b7fe463384ff4b = I9518532a8617fc8290eb6a5e981dea94;
assign I1c2674b2e6b269ed539827412c5199a5             = Ie7554e9d2bb6287b440973a9effefb50;
assign Id4fa22c6f8634ae38892953bd6ab55b5 = Ib862ac63c230ccde7fae0e62f9d047fe;
assign I10f14b6433498e3b9e9bf021b60115e8             = I3fd483389e4ddb927e7be7636441f0f1;
assign I3d8295457058e1d34bb136753b69aaae = I013d84bfd582acc7accf07ec522961fa;
assign I0236c912c6d684bf4862b725be9d5951             = I3d7a6bd63d9f66b068c08cf9046474f7;
assign Ib8df0659486e8ecfb5c52bc2db3a8436 = I7cb58e4c486e683faa4acad4756815d5;
assign I92496f68b44a94565af28a2c28d6fbae             = Ifdb5bd8e8237676fd8d2816bfa53f0c0;
assign Ice8927db6ef88a90daf77ea5be2a34bb = I67d57e38df8cb35ca686ac2eb44e233e;
assign I964e17c41a134c080e9c43412a514f3f             = If2865b698bf9c511fcf6724856074335;
assign Ifde5beb333f350ce581a137dae22b99b = Ic0c13c9a929c8c46e8702cef74de8955;
assign Id023a6298e65da1f4da3831f5136afc2             = I077ad1ef2fe0a7e791fdb45026788641;
assign I9fe47549e560319ae8decf04a9db5240 = If66524125bfde5aa48ac70c4e448b38f;
assign I6a3f405bb4a0c4448d9b9d3dd95d036c             = I4c67ed6284da547b599a4602a3cc51dd;
assign Idcda31b4dea85b3acd88cad806aef569 = Icddb43f9b760a4597a0bb637fb405616;
assign I0b56aa7a1b7549c91dddd3a06ecbaacf             = I3d0babc64a3400a1ee57fff14920d1e3;
assign I54da9f6048b299dd7e94962912b86407 = Ie41ca18c7d11a47e274f9c33f75393ec;
assign I2ba1acca919bddcc22a41a28d43a4e3e             = Ica1731833fd3d6a881b3a17a5916f7e7;
assign Ib1da5f847077624a37594c2db1b444fc = Idbf4ad11ab2a27044193448c8739fec6;
assign I7208256bb198bfce1be71390b01bc028             = Id5705e57bc5c050342e82a302b73902e;
assign I80c640a2bc35e9012dfdda839dc5ed1a = I04864c28351edb33b61a103add6fb875;
assign I9015033ab0caf3fa41dae4de43f24a82             = I4606e0ec878c615753206459716b5d25;
assign Ic81ffedc7f65fc4d390acd0a30d5e427 = I431fc2e9533012c8571d8158d4777dea;
assign I5149125aaaad943d891df6a3c2be93a0             = I5ac4f231a175a60f63db8d4d71cfabaf;
assign Ied3448df1f31122d619b1a4cb316f200 = Ic3ec6375998b05a3e48f6c5fe7b3910b;
assign Ib528bb7a64cce4f694081d151fa6fa86             = I26a3cd9ec3a564df04ad20559039598f;
assign I017d4243cafbd5d4d615393de3a29aa8 = Ie95662d4faf6b5a4cd5ecfa41697b983;
assign I735db8b0ee0ec98e4cce0030b11508da             = I26801bb91e66797982b66ce815da85a8;
assign Icb2adb3572c2ac780b4fb413c6ebb375 = If3b77c41fabcdb283f2c6fdacaa5e9a4;
assign Iaf08bcaaeb15bb0c971432f7f8b16d0a             = I3b617a013c15e8b623ad517e08df3a00;
assign I711042dda213300a90c51b09057b64b4 = I6c765e677f42fe600b848698c8a78349;
assign Ie1681d905517daafcc7584725cd6014c             = I65f5f9a3f7f68f4b2fd7695ce6bf4629;
assign I59b7772e832e814877d4f9e7726f5143 = Ieca2767ac27170058499d83016447aa7;
assign Ice73589836da9028def6efb24a04dbbd             = I7d405b59e360b17d7f2eb1805b796fa9;
assign Ida6ee8eeec2fa7a6bc1eeb8b5c3fbffd = I403303228c0df825f67436f4a7e64061;
assign Ie22b94121b58f17af14c75bfb27f96dd             = I033ad5c570f42830b265d7bf6a102757;
assign Ic7fb6a8351310bd93953232556a692ab = I0ac421af6e311b6005c3e02e93ff94ce;
assign Iaa40bd3abf668a21e0f87c7bda7b3f69             = Ia00376ef5aca6a428280f2dbf25ab1cb;
assign Ib2ff62fd117b50bc0c190b8111b85f4b = I849ee5d34760be03d4285185136aa52e;
assign Ib1a2b31d49ae476e2f1fb9acba2d5af0             = I252b17144e39018fda208bd18b555c09;
assign I4d46847f77bb17019eaba7ead1549a87 = Ifb422c30663eb4824caa72326b238df6;
assign Iadeedf3870f0b1eae98d0f7dbbeff04a             = Idb756c313694457c14b02431f3f076c7;
assign I1d6145f5c5d5049a1ba3f3ef8a09924e = Ia98de3691917dfb63bebdc3f8655c8be;
assign Iaee6d725a8b2653eeac6d5acb91f8f36             = I0c1545b312d755b14ee27b399a1d3079;
assign Ie5e08b5111cd2baacecc68000f84a9ef = I67f87fbb746dd937fffc534c596f36c4;
assign Ide604e9bbe35cb55892a4602e18b2527             = I903842d13327b74a952be0aa6c7ab0e8;
assign I3d61c9137cc0cdc892bc50c659fa8c47 = I23afd747ecece714e32fbb896b5c022a;
assign I6e37582849c2c98fd15ad92d22c222da             = Ic461c1b7bd09b59297193d388c525ece;
assign I15411a1495f104308964c62a1ac7fe6a = Ib9db80f43718305a8a8774d8d80c86c9;
assign I919d36a7f6ad42c4bbc23222beb73106             = Ia14490057ef27f5df5f1b23ca6440a65;
assign I99f350aa0b468f89e8ac4b3da627a81a = Ie6212a29c7c6b035cfff4c869f945b68;
assign I42f9b1f8ef24ad56c10086852678b456             = I2d3c1e36bd952fdbe4fac5f3af07e666;
assign Ie23efd54df7880569e2d45a8572c02ba = I41ab6fb6ec6ef7ffff70e50f25f217b6;
assign I70ae07db9b44d530be220f06401d3d3d             = I7fcea0a5f9987b2414ab443bd07c05ad;
assign I29de3d73d38639aacb693c8080f4a168 = I0bce960fcc58938e6a1e01b912eabbf2;
assign I4afdeba4fc2a12a6cbe3567a519367fc             = If0f5bf08d96033f6281121230c1e47c9;
assign I09fe5010524903c8b34892f6c308d670 = Ief72606c77113ae37845e4aa4a2ae5e7;
assign I770dff588ee1f52f58bea1921cb23383             = I19412627d5c573ceaa981cd7f1027e83;
assign Id1af840781c6093921ea2feef85b6bb7 = I5ede62333e0f7ddc5446b653ba9a2382;
assign I140078292f7209eccacd53a8bab18016             = I7c72a1709b233f745fb0323d04bfeb1a;
assign Iab8c6e113a90faf59bb550681b0dc7f7 = I3b775b06b5d78fcd7373c966a62f44ad;
assign I648d2a279dd1f587b1e45eeb35f2fa90             = I2639cefc25ac6f4982e4eeccf8fa810e;
assign I2110f3928229bc70d8ec9ec7f1c92520 = Ie34534dfd435b3d1cf35e82ca71e83ba;
assign I856fa68463aa5ef1ae53442699d38b33             = I76340f05f74b295583bd9353884979be;
assign I0befd079483b2da8d410fa137f71d801 = I0ec27b590ee6dcdd9c1086105e3b6c23;
assign I6f3be51d69b2b64a04e55b8946d5dd56             = I00974459262f29ec2b5472472e49faf6;
assign Icd1a2b8c1a50f9a1bab48ebfbb87ca73 = I452e51cca9acec44e36e4efd21b43034;
assign I66528f43f614f0edb715564eba3c77c1             = I075efbd3c4d87df8d733f0b3db008b1f;
assign I4422278d28ff2a983cc3a4ad8f2d655f = I946246be5b4745508b7d4b578f83aaa2;
assign I0d9f8c99194d9d6e187b4ad02fcce8b4             = If8bd6a5d380075f1ee7f7a4542531dbe;
assign I3fc4400a93546df2e2aad374a4d8c7e4 = Ib2fe0f68044c11f879e512a200f8099e;
assign I74a4b9365391fd20c34588002ad40547             = Ib81b730d107434503c988ab9f00e1605;
assign I6c6a02b572e98d30ea5a0406be5cfd11 = If2372a5956f21f97eeb9c76281b6675e;
assign I194a64bef92ecf6714141eaa5d41c9d4             = Ib05cffa1bb31054450391bf9e17f8ef9;
assign I91c29953d4b53657da39b53d8c909fd8 = Ie596289582a73e37f78f4ca4cab21e3c;
assign I7d9ad929660cd212387d893266b681da             = I627097c06e3be5a4385171f3ec7ae5c9;
assign I10441dc2915fcece28b38aa6b4156f5c = I7b80b4902fe98c10dd72c9eb082346e5;
assign I62d8efd4227cb3dc88aa08b6585fafc8             = I76e2c6001e1ae97670539bd471fc74e8;
assign Id26aa7283f70b13f1eb0b97ab1222da7 = I3051f561a5e1131ebf167cb6ccb5adf4;
assign I49f2a06ceb3a59773c65b19f54ff362b             = I8b4433056d26f4aa60f18418b0114930;
assign I98b4bf6c27d9420941d252a98806344c = I388528eaf83566cc56b23485a9c05962;
assign If004de0cac6e5f7701a1fce48c6936d5             = I99601176686afd8fb85a85ec43849e6f;
assign I7814b43f7573d005d6b9350b311f93df = I3ed6426fbdba8aaf1c948cca7442b3a6;
assign I028ce03be0618b816e0ecdf43d4cd6e6             = Iad8276d5be3d9c6fc085465f05ac2aed;
assign Ia378bb83b0f76d4bf7de347a8bfd20cb = I7b32c2b108e24750e2a24785668af3ea;
assign Id332e7f482524adeac7f7cdafcf5ca46             = I5e5dfce3ceb4fbbfce344bd471901736;
assign Ie814322ac906e4bc9baa42fef66e9b8e = Ib81431cfb3b281555fa7e5b4582a2524;
assign Iabbd1668e0014df518ede5216232834c             = I22ace766690e445ff36176eac2473368;
assign Ic3f5c7e9a546509687973efde6a8a8f7 = Ie5373b01a92f2ff85be8077cfef2175a;
assign Idcb37cfc357cc088c775409fb9225b51             = I896c57162e4384f021d822789b4c01a3;
assign I5a7668981b781cea8cd3de0aa6687bc1 = I284b23051c85300c2a1e3afe8f25e99e;
assign I2ff3edcdb6158f1e3c9a555aeefc0850             = I3d0367a799090b3c9048235436a39063;
assign I4951067363d095f73676e08c2be255fa = I71d7f72d83b7410de31e09ea96adb95c;
assign I6b24690f394792edb0d82b3b9e110851             = Ic0f25799f0dc7cc33de95e47ebcc083a;
assign Ia02db0467aa519e8920344525ed30dfb = I4af3e2bf2ebc913ac902b48da672c5b6;
assign I63e45abd4d27219bddcef06108b72021             = I7186b368e297d0db1f746c6241eae65d;
assign I303114e80311c7f6552446bbcb0fe6a9 = I8ec99197a7d823f5745d382c10161430;
assign I226383d68f89db716cfd8d08b837865a             = I21d63f6fe5c72798aa4636527c02613d;
assign I7a5c09537045dcd633095a86a6c530ed = Ia3559d98eb372b7307f30ad1f7c4c7cd;
assign Ic72f41f9bbf470aee3c9b9b8787b31c3             = I15e0219f2da6f52177e76580198d0e6c;
assign I6aac30f1ecc270161a81bccffab85efa = I0e8679271ba733bb87c44b6b9f0b6ed2;
assign Ic3d00a27f15f8983a120395082854d6b             = I4cac308bee8801c4f9716673e39da4ab;
assign I79b86b24bfa472a80487e7ea64f9dd82 = Ia7c9c24f8e993526e76c6915e56908c4;
assign I19bba6a58ad3ef959b33701f82761984             = I6f4f7b4e45a495fe139955e0605ff208;
assign I208d1c07cebe2f45b25b562dd9109f7e = Ib895fec0b3756932b85962c1d129a03e;
assign I2bdf5d319ba9089a4da34b108f5c5ae5             = I79ae5f2981b7dd91141b0a22f012f4b1;
assign I86a3b6dc06c6c99cb1fa88023d920423 = I8f1a8a22637d37c3692e808d5eb3d543;
assign I96008f47b9f134c9c4274cfcfb28e550             = Id4b4d757e50bc2721e8725ae10d88c9e;
assign I9c0e0297c0e5042f1ed791d9d97a6f37 = Ifad8c7bacf72583f91be27fbe5b7a1e1;
assign I34be4b353cf75603301372840c2f91c2             = I4513152c34d5d00ddcc4f099481f659d;
assign I3af891fd5da91085a79886d82e6bdf48 = I384e50fa8daa639124f083dda56fac00;
assign Iec71fe7fcebccf1ae0d10a5d187fcc44             = I7bd4e77993fdd5a0833f1cdc7a382b56;
assign Ia1c63f27861c8e594f01ffb31a29ba0a = I76aab345d13c6678fe37a4a7133cfd7d;
assign Ia91800792941ec7cc60415c3f844e4ed             = I13b0d404e7a96cd53147b574b242ef41;
assign I62b87c6aa6ba054ab5e80842ea738020 = Ic76e72b434b47c10ebac3fac4ea50bde;
assign I71412803cc5229025487255aec62ec4f             = I4acc3bfa99b152c6ef6d11608f639b70;
assign I429241122829d9e51a3db90b33a44ac3 = I835b902949c2c4c09b757d4d35574a76;
assign Ibd89458312687610aa166a9538968851             = Ia1ec7ba972ec6f0049c4cf00b9d42125;
assign I162416616ce392c679d22b115c192356 = I5f1609647f1e71cef4ba2d605c6c8445;
assign I1c3c4ce44610e04c5eef2fcbc2ea5114             = I4fb5494e6f04e29d76bb8d3bc8bf6cd9;
assign I62edec03adbb7bbda313abc2220a6a5f = Ib4f368fa3d3ec11d9ffb2ae9a2ae6310;
assign Id7c507d96098ee7a955af8a48ee5d72a             = Iaffb0ef4e18bb7b582275b43684fcf3d;
assign Ic3e192f5abb5526a54ea249e736702b7 = Ia1b617e3d141263b51e58c5ef0bd7a89;
assign If1607e907e626902ee26d15020a64c21             = Ia5e3649f8e32a81606ee34353c54350a;
assign I1ae99cfc5ded208c2dbadbabf36fd629 = If343015b4815b01dae88bbb6f2017b3d;
assign I3ed5d0fca86f35b3d4b4a89c6147d0cd             = Ic675cf7eac5ece436feb5a8acd642f6b;
assign I1ef8bfbeda31b3dbbff053cd36de4859 = Ic98f33c6a4613534bcc9b6bc4b4f2d17;
assign I599d01cfe6e54d8e45d64446c446818d             = I71357943bbe307c9ae9099d4bcbff882;
assign I6d76fd8af44893ab0f82a282aca12377 = Idd0f3cfc5599481c954a2bfe69f044e5;
assign Ie15e4c1bcdb0e18085d4b320ac6a925c             = Ib2684f54caebb1a1c079a2a4f2cf0dab;
assign I86247340bd399afebac1ffe403a3331e = Ie74c72742807ae4243748fd27d80d626;
assign I14834fc8e6489775359bcecf5a37ff4d             = If19836577f9a254b365f0dcfe0ae55ce;
assign Id932053ac235b3035e2f3d5986b7d398 = Ied8bd4b6fd0e4fbcced6d20eb7435f55;
assign Ic87c3d7762a18772972552162e1d1a8c             = I2f47a00b58779b836c08b472d305b031;
assign I4b43b5eb71dffb4bcb9ee541a537b427 = I6cbc06919b9c695d99621db6f8d768cb;
assign I157fdf8775206858c08682db3039b084             = I8b2593fd0e35c37f68097187a41596e2;
assign Ib481c772e0ef5d172f6b079dc8df1ae1 = I641539560711ff1824bd90baa0f21f96;
assign I8f0a90e761111a613d2488285534a500             = Ibbcdc1c30d3333cbec65d264890cf3e5;
assign I2e046a6e848cf2da29e103872a10c26d = Ie624c4dad5036a25ca314b94cf3c4b95;
assign I5485d9edcafc6202f6e5f0969979802f             = Iec6e9640b0494777c013c97613855ce7;
assign I2a64ca51e05db642281525ccc7cf9a06 = I8510240df7dc41f85ad58a39868a1fd7;
assign Icbaf92a8e9875bcb19a1d074779a9ea5             = Ic10f396b52dda0dcfbf2a847cfed617c;
assign I4275f1683058cfab72e02f2631d2ee96 = Ibe3d3e6bc58efc2e9d9eb1f96cdfe424;
assign I20c2057240417146df144b518b43d052             = I94ebfb633f3272b8f40303ce768f0ade;
assign I592fab4d3d2c1bb3956b89eabc06dc56 = I72939e49bf2d9c6a84e404419fc644a1;
assign Ia30539545e66c4cfc16828140149180a             = Ie975a6fd78adbad8b8a56bd6a3802e4f;
assign I6520a98d1357fc57d687f9ea9a60508b = I95f0acd4f955058041c035789c3a4d99;
assign I71e101962e766a4d1484b3235359a4b5             = Ib852991e38422ba6de5e18a879ddc3f9;
assign I8a022ff37fcd6f34531af4dc7f31a223 = Ibf4b3caa5655cfb6663f9b7e2383bbbf;
assign I7fe364f9f537cbef782e7007848a1c10             = Ife665c9aa6794cccffd04923f4359047;
assign Ia95cd411b17d1c5aaf9e5b583e9398a6 = Ia0116a3cebf94318ed5b287960957ad6;
assign Ib0126fb335e32793c400a97c5a4a337c             = I076cbc669ff4fb135ffc85910c888241;
assign I526597e8561c75326b96e85743420a1e = Iaaaf373f7e6f55214915b93da9bd71d3;
assign I2993acb61f1abe529f8a60c94a438550             = I50245c953aab8c513b17b894afb36a6c;
assign If2c489abf57879ea491d9a95ce7e1cc1 = I0ceb14ac0187d804f9692e0c55b8e941;
assign Ic3b4752136ac08e343933ccc3a4ec47c             = I33ac557ef59d79e8b1b359e499a00119;
assign I1dfa9cd65fb0f7c62439bc0d9539e45d = Iea424dd9d8916c4951b8746408b8a521;
assign Ic1efa395cc1fd2c5a1d1559fb169a5a0             = I173fd30c1a5367b61e3fda352365f557;
assign I5799e21b9e2fdc554f8ec65b98120544 = I049d1c09c15def12ba7bae95fc1c3d55;
assign I52dcf5bace9cadcf8a895aaa6a8c1da8             = Id6f5041043fa4fd352e74016c4e7de48;
assign Id109dde61c0ee952c9053905ee54ccd8 = Ic14760b65c6fe150c3c48e64389a41d8;
assign I6b1d01c3cb8fb51e43cdb788b89816be             = I6d863254c7f0b52f803b2af4b184f99d;
assign Iafef3ac31f22ba4f5ef06b13165e97eb = Ibab1d13cd6a4f7b0c79c9f845339e53f;
assign I33b99994abbb5ecf8eed4de39033e4f8             = I1eeb9c94908cc9ddeb8e3904a145ec6e;
assign Ifc59d693d6dc2fa6848f37a134fbb316 = I2919272e9ae3996a3e1d602ff72ba86d;
assign I39e6d3fb468aa40ea73535e81556ea65             = I6211e241282624fc50fb4ca1842ff9db;
assign Ie83012a17bd2730837939cf0454395c3 = I1db4ea6916125702e7fb09d0f742e60a;
assign I5b55c285f7e3e78447fee68532ab9f7f             = Iba09e22ece1eb1639d2bb940d3273fe0;
assign I1f37257664651a57575f7ae53ab4e180 = Ide06ba186ddb179b489ba6e3e209e3e8;
assign I13a9eec6175e695ab8bc4516cf57d6ec             = I2fe99e4fb8c660d83508bff50ab4929b;
assign Ibdf8f7dadf142fe8a166328bb5461308 = I6f420c64640dfb0c001f57df7e3b4504;
assign Id0344146d1a53d418add6d2b185377dd             = Ia73db0428763da3c0feffc94a8a8f4f1;
assign I0ce12cc00bd66d743ab82e89887190dc = Id75c23e80cdf25d883806ed20d4ae783;
assign I20590d8fb97ec0b2164ffe17826136a7             = I6542fbca90e189048b15deaa3af5d836;
assign I70145dd478e7f0c74c0299cdc0ab8ad5 = I4d4901ff372f6820ca9c8c29cefa664a;
assign I05370777439b01811fe7f750d2f724f4             = Ieacf022fc976bf397946d6481468d6a4;
assign I03d54826d217e4209d0e0f82beda4100 = Ice0234f25de4ab1f03a3cb01a2d61dbf;
assign I8cab9fba615b94fd4bb6934325be8ab8             = I1cef7e6e0555e076b68bbc57de8f289f;
assign I0aad448f6b0692670432efdd1b92d115 = I1b78785ebe2e7f77a3125a6334c4dc54;
assign Iee73a7c685a4cee03f33d3ef379b1c8a             = Iadaaac832a1422494d4206edee770d63;
assign Ia5a7e36b324b3a34be321ef63db22f50 = I9eb87e62d23bc87d7cd82c0f329f247f;
assign I32fcb28a27356bc6f403528836ea4c1f             = I905b0ec8983ba423798bbe8282728af8;
assign I01399ecad74618d26fea1ef278a3125f = Ied6c684cdd280b41ffab93a026d27282;
assign Ib74a56900c1f8b159ad381f61acee801             = Ic646b82fb6e3d0afb3a58c4e0d68f06c;
assign Ia56986ae4171b36a362b170920663c44 = I1ca188bcdebbf41d84f7a5220bd1d195;
assign Ieb38fa62119a5a77c060d6634e051298             = Ie57f41c62e23092974664f967a27566d;
assign I7785a1b6345c7a2086b3d2a032970fa8 = I9322a2a61900943075bbc23c72a3f65d;
assign I86e495dc894d2aace15c1aff89798bf7             = I34524ca1dddbeadcc060954238175e7f;
assign I778c7251ca1b16e1ea1a4720ec7ba2de = Ie79c93f1703121713fb9401617f349a8;
assign I740dc91716e3906ad078e2c7cc3c925a             = Iaf2a93993f99814321951a6bffd8bdd4;
assign I1fcb2b0e5beab6a80ce06aeca85610b6 = If9a5d830e3ade0fd96b98f5949f165f0;
assign I081b38dbb37d4c14a6a9fd3fefa13daa             = I97e4f7a9a8a42be813c6e4128936df3f;
assign I3f8184c2f7e604f0581e5c02f5b9563b = Ie7a68c2b368a295f95571bc4a109b9f1;
assign I633a74e4dfa841c9fd13dbb6564c8493             = I682a67100f862bac0155a870cae0528c;
assign I25be48f72f47043fb6e8b7f774db1912 = I0152dc6e6a7acd72a2144623e63998ef;
assign I0b7b4c0a8503c751229edfe0237cc903             = Id5296b03b99bbf52d3ec04dddf3e84b1;
assign If75d53ea58491447eb2344e993b4881e = I9b560d9baf8a7422b0dd84720e924ced;
assign I43b380be6df7df0d354223d0a0d6d6b6             = Ibb089d47014f9002f2ea6b431156d9af;
assign I4951621739ec145bcf3004b0f72e26db = Icf25f076eec2bf81c899c66f6cfbebc0;
assign I514d2dc697e9b39ba027c418a6df6cb9             = I83496522139d35aa028dc9cb8a78d442;
assign I959793f388e50197e4e31dae019d64f2 = I7332e088bbff69db19c62685e033d26a;
assign I3ea4c33a9419820ed54460eb64134dff             = Ifd4ca5a83fa0c09b043ad54d25971410;
assign I8bccd3ff9583b2e33bf26d779f1c6233 = I1b6abc8fbab3849b285e9f88a4fe867b;
assign I80f3c8559da8e97bc5397bb8b621a0bd             = I6efbc715be55b616551a7d4650a446dd;
assign I177f26189ade299e79c1406cc8171ae0 = Ic14f948884da19a272a4760ffaab9ea9;
assign Iaf4ae293c576af16f5f43a8b86c1aa3d             = I572bf74835f5acdf5a17de2063c293fc;
assign I93f3cd21e4819405b800ade59c9ccdd4 = Ice5f7168aeb940d48093cc9df7cba36b;
assign Ib42816335dd8475dcc78662c4c0786c1             = I5f8194ef67d22bcd38f415fe8d9a6ce7;
assign Ie655403fd0fb16aaa04783a2ff742064 = Ic5c837a0556d1cb66edbf0294d08283a;
assign I782726e317a2aada9e755bcbc4b0d3fa             = I3d3f2dff1f64ce14071e5f315bb8a57f;
assign I1c3163e355c43d0a134c88fa671c41f3 = I3600031716c2b4e21c9f577d34e033dc;
assign I1eede74f12d37331b399eb7136bc621f             = I8e3880fe0374bc068ed14eeff9f6d009;
assign Ie378961bdb2de01ac733e765bba5eaa4 = I859d795a7d141eb777c1f3c038203794;
assign I343c9efe71164c01e9c7d599e032864a             = I51d8f49653c7468b2923390dc5932a2a;
assign Ife404037f29f17b3edcc4d1334298781 = Ib9c194ec16f435a9357cb344cf25bdcc;
assign Idb72c046c5996fbbd80b706666ffbd92             = Ibeb380f8f935c8e061fe00734675662a;
assign I4109fd0e3086c344f926c4a83b378296 = I69d82ab774d52c219509e993e7cc4deb;
assign I141fb1cbe09f9abe282cffd4de815d25             = I641f4280286c9343b7ce001a8b43fa21;
assign I5d9e11667955d8128b76d9144463e59c = I51ff4bda38746682e3cd4c68118c3216;
assign I11eb26cf0f0b3a334e8f7317bf8d9eb0             = I796970d7c73d8fbd7d25793d0dbf9872;
assign I70c06d2f51ef27666c8c39e0a13ff5cb = I2eac5b39c6f485c9ae0bd341f894633d;
assign Iad354d876cb9fc72fc0143e6f7da9357             = Ied0b1d10ae09c523d1cd1cd3e5b184c6;
assign Iacd270f7fbb94c91757a4f8780616e1e = I12a18a1f8d4416e9bc8abee6ac3dacfc;
assign I92d9fec22d36b1baac8bd78abfc1bbd5             = I7d0d39d94d929741158c39f69e8169e4;
assign Ia95e1a8c5bce4673824d56d6fab81f4b = I45bdd0cfe107da0d57cad1333bf95e3b;
assign I262f2390e77ec486ccd3a6ed05816e2d             = I2349636f6ea8796c7b798aa555641a9e;
assign I49137af52922e3872901905fd7c70601 = I768720af835b02a8dab376ef23d17a15;
assign I461195b7ae78743e09ee50486ad6ebe5             = Ia3739201eb91605fc115bf320d4c24f0;
assign I548d9239de9b536e1b581327961b53df = I1c074a53e6c0f2467bcdd7c952f51670;
assign I26cb63ba20245b2c332b09e25c4409aa             = Ic74cc511acc98510da011e126edaf3a3;
assign Ifad4cf6d79d76caa33927ba4a6b94b45 = Id3de87169c440f95d406693ef77cacd6;
assign Ibac5e7b6d4bf5cd6926358318f0c418f             = I89b1312c0696711956ddcf787e37f3c9;
assign Ie78dd544469009d2b182d2b76694df6a = Iedc463e359dd3003d9f7e50f3e858e93;
assign I0d53bb5344cabe5fa5ce3ecf7122a260             = Ib2ef1187c1743da2cd83eb9231a7ddf1;
assign I69122b791a8f717c501f2842240a51f6 = I23955b54e486f0f0d21a2809a9472b86;
assign I94f1724740defe5bb7e40041d0e266a0             = I21710bdb6874ab83e2b2a2cffb026ab8;
assign Ib89ed0cfe4ba481ae28b835d4248babf = I24075f37c6bbd90c83370de1a2e58af2;
assign I6ae2523095237282533e0b5f1c26b488             = I2ec8afd22c84596550412a5d2c7129af;
assign I6ec25bbba8c41ebdf4efa95fc1d8e1b0 = I37c49c5a2af240496f5a5706b0d42ea6;
assign Idd7691d31f8d0c09ee988116d574ec59             = I57056cc2fd4bd1ea6e980cf90c22e871;
assign I92953d645060c118de19fafee18e34a1 = I44daa5992b00e7af19adbee70bf01f2b;
assign Ia0d940e16c8cbd4f7544f5a5cd7d83b2             = I233becd31032d63e65371119edb2cf79;
assign Id89c23eca2ed6103c87dc296082605ab = I457ae11ad90c8478751eb4b42764e158;
assign I23eb1dc4d1c992f804dd04a2d823c778             = I0142623400f5994f581a4797fd9d327c;
assign I070e631601f2529f8f18ad0be6a70316 = Ida3dd5e990ce3c237e9628a9a090901e;
assign Ia630e59cbce82a570ae3890a6c0221e5             = Id3e298c9f2709d8dc01c18626ea846e8;
assign Ie1e3e5fbe2e2ae4cb3218616bcaa0ae1 = Ifbadefd3a7ab50719a703400ddd742c6;
assign Id1bacd13718f7c29c26b63c239d04dd8             = I1044e090bdf84a1bd30438137d6ed056;
assign I6b2795593e93e47b2733c1e0003a7806 = Ia94c439131e1df5c95fc8ad3cfdba473;
assign Iecc02842a2d2b9b9e8187f2d39e62e05             = Iff0f43c1fb40bdb3271a3a38d89f4d6d;
assign I467646a701c26d253f43251aceac9527 = Id88a7edf897eea1b4a137141789a04f5;
assign I157bd468200e63385583b9045758d81e             = Ibc71a0c3641097c144513810bc9a0a7c;
assign I280a8abed1540ebaf599c094a0a75797 = I70dd1350d65155ee7b562f4c79024a3d;
assign I09e9a3cd4c12d204f760758e873a177b             = I6ef3b025eb065f833efe6daaab699efb;
assign If75560cad0cb26bd315f3711d1e9711d = Idc445d3f5b3b62562b0ac83e5f17e92a;
assign I32701d9e4b96853c53f0ab651a6a4ba2             = If76152e9435e7300b19095a9b070e0f4;
assign Id0d79e0b7361bae1b007c8a7d606f6fb = I723a6fee3b2496f23c48b3584f8bf9ce;
assign I5551342f1751fc64f32744a46b9649be             = I5fa63303ab85db9c8cd268528eb604ca;
assign Iac7bb2fe5935b53852a63923c53f13a1 = Ied638fee34f8baed4154b0b72e43a21e;
assign I7a0eada108891aba06cecab5071232c9             = I69d6adcd3d35a24b393e97ed6a99c061;
assign I4554a553586d9966e7d4e8d99a5c799d = Ief03713f5cf37200373a20d42c7fc9eb;
assign I4df3d4dac24877b14e6d361bafc1a800             = I8980eca0e5973840121576b6eaaab736;
assign I84a85d995e807610f153e72ea3df3ae0 = I3ac0799861144b599995318bdade2114;
assign I765a8825e42180a6c63f7b33703bb483             = Iadbb5c4f7b7c02e151d5118a7ede1f0b;
assign Ic68f898ba0d0073df41bbfae0944c9de = I648b62fa0bc2185c1756ee531e8e34de;
assign Iff7c29299f005c1cd5a16b64601e727e             = Ifff90bff22a3bcc33261004136d2e655;
assign Iab98e00ea4dca63c81eb8f78a133b1bd = I1b43f29e0ddb72467befd6f3a9c1c829;
assign I3c128efc9f80c9b8334bf7b61de71b43             = I8d13628f322640414a4b556ee48d3bdd;
assign I67aca5b07f66a9f3e8a5550020802c63 = Ic07c650e6e49892a41cfaf3a37471426;
assign Ied00d87af99ae55144fdde41ebfc1357             = If7d187cc56b1014b1582c5f5b94759f1;
assign Id4b0e0110bcd34cf8f0a9a92108b88c2 = I4082b3564c1949a19ed35bd5a88e1ef4;
assign If2539da6722562bbf31786fd0036666a             = Ia01d5a33078abf4b2d6c625af01c25f6;
assign I29ee6514004941d4280cf4a93e7baf5d = Ife631f9a3c4c64a3d92aa9586ae75f3c;
assign I17a5446e942bcc1dc2c96930e0a87a70             = I4c74240688b5635b5323ce3a8ac666fb;
assign I3bb0ea6e5c41271be14ed45d4b8ece5b = Id0f4dbb72da33748d8baf723c5a32567;
assign Ia5eba52d169755c507b9e0094e467fab             = I943e9afa0dc80fb50b5869cf34726823;
assign I0a1dc75c36d5fb043c80dde4e8c5e577 = I44ccc3ae897109dd51f9afeef93daca4;
assign Ib9ceb8315f0cd848f861bab677c2c694             = I44d8779f30245bc7f1475e6feb762cec;
assign I89e39167f230c52eaf64e8c5ce8fc38d = I73bbf90b625d56f663ad10f9d21d8e76;
assign I8e96c69e7d872be23229353808c34953             = I479e7456c445ad604ebc134872a0fbfa;
assign Id6e88b1c05e5f4e7188f4b646f428b55 = Iaac1d82f0846fce1bd88ebf8e60300ac;
assign I719b67f84e07e90dfd29a8cd5d94cf39             = I484f372e3a2e74e0791b06aa666b781e;
assign Id9b024743e4060a62c6dde2646b5c998 = I002820a37fa7c6c504c487df4368e2cf;
assign I3e4754acc31d99bc71525789bdee0c1a             = I64b07241996c48963595f28e35a75be5;
assign I2bc4cf6682dca441749b95f63592dd8e = Ib0bb71b1f8829347b3a9a7543f9dd964;
assign I0899e8fec1a7209cd94757c0b2f87c9a             = Idf678798bf4e1cd316a49a2b413cb29f;
assign I05d8735777c75ecc9f1e5d2f972f5c21 = I1dd4671765f8826c2fe20c592c5e32c8;
assign Ied029d0bdea3bf134744c99426fa72dc             = I35fd5e5e93f992ef5ff6b11f9d69609c;
assign Iaa201a0537ab3cbcb5bc065871e0153b = I3175159add7b814df637c2db8feb43f6;
assign I5aba6218461e8d571be03a3ef041ebaa             = Ie72397edc1c597c0a8213b67a030a482;
assign Ib76deffcb8cd38d5643df9447f3b060b = I48cd09f035f668536cd288a23010b07b;
assign I2c835dfb3596b8bf057a7cc21122c81f             = Iae50178e99a07cee0eea6f7cfdcedf1f;
assign I6483a59c7f2bc77b445b202f0448eb2a = I76992221b1edff5684c482df7ac4693d;
assign If6e745bb85abba7282dae1f6f701225e             = Idd7082c7a65d7f8e0ea88142312a631e;
assign Ic1ffdfe961dc8458b1d4cb36642a386a = Ib13436ad16a37d656d6b1ee95b9aee20;
assign I918c46173eebc5b2a95e041cfd91d958             = I4b580dc4cfac9e9315d03b60e2a915d9;
assign I0fb493a1f8f2810ddf67a6cbcb2c782c = I47b0847946b0e00961233ac0101fa2a7;
assign Ic8be2c94235fb40f78da33179ce4873a             = I77cdc9841414221c3f6c3cf35397059f;
assign I2c555af9585a50d2cd6a27c223c8722c = If2042aede3390bd208a281f0380c95a4;
assign Ia3104c69fb4f7abfb5efa3874169a7ad             = Ie59619c3e78e616e1febd2db2fa940ae;
assign I5f93af2953a9f1aea5cf55a037f7af6e = I119b2e5c2fea5338244c4019884af26f;
assign Ib71b3d357c98dcdfae5c777ca3082275             = I5bc8079a5896f59bc6137b59c4b7e750;
assign I25b3e2b9f55ea811784ba8ad8c5f516d = I3751f191f5009322acb7c9be4f8d7129;
assign Iadfc60386481092ae85cc148a2c40abb             = I239bf978d991f702ad23bc6b4b8be1dc;
assign I93fb55e460d75b8d36c19833849bc1d2 = I14fa7aebb608d4a3d67176ba27d34d9a;
assign Ie21a2c9b22e7bf8425fb5c0f33e5f4f7             = I450351fbb31246b49cfb2d622b9e90b4;
assign Ic51082943371a401c48202b4e655e84c = I7b813d83b13bb7bc13940cf5714c06ba;
assign I7c3291f0250d13ca94802b0b071a95c6             = Ia7c17a0979f3bbb9e9e821bf69a239b7;
assign Ib53122ae54dc4ac5b090ba8aa3ab9959 = I0eaa22f5eca8f33dd254fe241017a098;
assign If79d1d378f7c6fd29fc3335ec5f5c51d             = Ic22975c34b92a39bc8940076e80d3c0b;
assign I459abcd025ce92565cbbfaada735a325 = I2bd34b2fd12f12bc301fd0d5d69c0fb6;
assign I086bf19f620c8a8f6888e775cb1ed7f4             = Ia7be8cf38ecee4568a939cb2ef727619;
assign If8abbbaf2986196395e63aa49b1022bb = Ie517386cb5832e406fefc5e85eb2e7d1;
assign I4a8abfa0896ce414d9b98093ef84455f             = I3e475cb1733d494f5f7c4b26a07d5852;
assign I830ffb778558295001c003f114b66198 = I3fd0fa3b774d30a267d61e9427d09f3f;
assign Ic7147944f8835e26b9838fdbdc18ca41             = Ib2c0df16678f6aac19f7af4ad4e53ef8;
assign I56e732494aa029b716ac04289d951e27 = I4ee312036de8c08300c358edcff1e1e9;
assign I7e393e6c1d1bc44daaab120d55f5dd59             = I8bd2ef39eeb7089409db02e3806956ac;
assign Id077045b00947ff1b4de86777d84a48f = I1d98943b01a6a2d8c4db18b98dd62f5c;
assign I356d747600182675699a2d2634d4c5ce             = Ie3669e34cd19462f524932b3d232b546;
assign I7ce7ba4f90dea6eb91d61cb456134df3 = Ib715b1e0061b84ce614a30d961a83e7e;
assign I802c554d5b04af6b949677819a4966ed             = I1ecea23a4e56948365dcb04c5bf6d6d6;
assign Iaee8dd8470306340982baafd8c9e28b5 = Idc07dc30c0a957e474546ac7a60df38f;
assign I4f8792c18bd07b23e82bbc44b4ca947f             = Iac222e9e39e300d7161ed05153cd9ca0;
assign I35088305c303ace3b0bd194f5efa557f = Ifc640243288c9b37b7eb9e00351b23f0;
assign I3459d98131faef5a5040a03847890b55             = I292683f8453be58f65370a286c1a4505;
assign If28f074339d099d0c8f0e582c11f57e8 = Ie83fa8157a7cce44c2e25f46ce897dbb;
assign I512cc8f6519aa08aee18225b56d47c9f             = I1dff7459553fccefc94a6020cc248a49;
assign I55b6efd25a905ab958ff62e0334d0116 = I570c036d0237c53bb069c52d621e539e;
assign I4a41999cea9357a85c73a0af509eeac9             = I9acec7aa4b420b7c820028b669a8bfb4;
assign I859a2864cbe2fffc01b411e7b0a2c3d0 = Ief8c2838abac83370fd7ec25c06d509b;
assign Iceefb06cb3715e1b41e6f7d89420e5ba             = I714b7d8b39c4135183b605dd97ff15d6;
assign I3ede6ae83cec11aecdb308142c26f6d6 = Iad90879acba3fc2101829549264960f3;
assign Iaa5b2807e5cc2403c5787eeb3d10ca6b             = Ie5856c36d9a310f890ecc5220590fc3e;
assign Icb7fa4f4271f536afd96934a45bbf0ff = I951dedd7af44c3865a8f36888432d0c9;
assign Iace01234164c8a9f7c98eeb83268745b             = I062b1d8d3b6fe6d8e158ede1f0af9eed;
assign I4dfd9e0bf539f3077f2d5a8bd3b5e469 = Ia7606050c683ecefc510ba92ac539a9c;
assign I22c8ccd4a9018ad1c129aa058bf579d8             = I0fbd5b5eef6da9adaf918390f6bdbc27;
assign I795091257b4f78363310623b731b347e = Id3b089fb6edd5bcfdbca142fddd5ff89;
assign I87d6a5d30c3e4202cf51f33c7a770c51             = I73fb14b30841cf67e96ba329fdfa3e35;
assign I6ff1f76a6ad568b5fa0cb300a67ceea9 = I561d79eb079915c0b1732cbddb119c2d;
assign I56948bc48c0220893d68004615a6ebaa             = I6d6cfca51988c5ac32471fe8f4399bbc;
assign I5864383518b7c9a70f69b0fd1a64d4aa = I2eb08ebaa07a1004638cdd61a7209b7d;
assign I698b1dbc9d8664d1c86c7a763d97b3b7             = Id7940e4951c96c3de9f45119043fbffd;
assign I30959187f5ac883ab77af90ccfce5704 = I46e1047bca2b38e62b4de80d1d2249de;
assign I68b575fcbc5321d4d26a22bcdbb506f6             = Iea71361c5f846419eaa18ae4b9463ee8;
assign I0d2bcd2e24e64ad5703a580ddc415f3a = I41796b587316c600bf583edc62649bd8;
assign Ib6aded6c73a8cc3cb964b0ae895b859e             = Ib67ac5fdd6e068ee799965b51aa893ba;
assign I4d1ef379c32f93cdd18e2415ba83a5ea = I0a569f6536789efb7ad2377c11842830;
assign I6ca8a1fa2c72b1c61d11dc7d1ba5f37b             = I0bd84509dde112f3657bd5a12a8df72c;
assign I921c8abbe15effa3769c5c3f81427274 = I8bb75bf828d5ef337fa6a965808e4638;
assign Iec1368f034655d61354ab5b5e94d7d89             = I2caf86026460a024f752fa71b44f743f;
assign I40cce0292c07026fb144dc28ba228485 = I47cbb92d2284aef7b9e56e88f0ba6f7e;
assign I08ece7cd684e593e02321612b7a88cee             = Id81d9c9ffa81c2653dea2e872ab2f71c;
assign Ia1401fc86b9d014a28f1c5bfa7aefc2d = Ib99e1b93fb7fbda260d93eea3d24c3e9;
assign Icdcd83341f6b5c404f91ec7e97d0550c             = I0b4d1a08307d452870c3e762bd038568;
assign Id3899a9a35b467c103ed0dfef20dd4a1 = Iee6e52d75c093a24eb4e5e0b45feb256;
assign I82f266e5792cdb6e7ebd264e246161f5             = Id75cc40233cc8648e21a750d882d5ed4;
assign Icff78887751d68045a0bc21e69047c79 = I19b73c5c93a71e90f620572f23f0e6d2;
assign Ie1b7257c99831ec5864f65958ecf14fb             = I3ea9815ba887e373a0a477654f136856;
assign I9a2e36db1aa972536df63a24462eba98 = I11ba339c8250d07b497c88a39a6df1ac;
assign I1e43c0aeeb8a2461d208eba24967af30             = I8b26e270c3ca5563da39e7092ef830dc;
assign Id74033401d8494d013fcfd1f69537592 = I8a4c1f23212ff846400651b100add502;
assign I11c1fc94a3bd6dffa17e1571cc6ae97c             = Ib03f94d7e5ff830d5063cd514e7f7998;
assign Ib64741c15a5f128b008851c36d55c0ca = Ief18a19d451f05f6051e3cc8de16d73c;
assign Ica6707efd6d44ba6bbb87c0593a3d828             = I00b05bb0b225b27562d6629725ac2126;
assign Ie75e57f87e9c8cc7d29519f0419f1b22 = I7009c18515dd43d8dd2e5d1ee6779641;
assign I939368b76d98b43826c68c7f468a5632             = I1f273682cac5644f1fcc30ffa20f8cd8;
assign I95bc08d218c4a924f810b69c7e2b923f = I173aa69cf52114e223ac1410d90b4bfe;
assign Ia6eb85b127cf9c1a437611556296b967             = I483725645504999df82a4d0660873c1d;
assign I6dd9a12bbad2fd4aded0354fbb09c6cb = Iada5bc4a51dc1bf57bb9cca11326bdff;
assign I93bb43c1b89d4c70a57bdc019d64fd22             = I689dc18b56442b8db01bd7ca4c44d615;
assign Ie78ca77c4a9cfac31f52cc1f49e5c6d1 = Ib6fbe376477afa58bfcc17a8564f78b2;
assign Iae449b74e50e0907feae9e60f2329426             = I805d665f394ff24f230bebfa6d252122;
assign I771cf2bb35d06a6009955936e2530f07 = Id48fe0672aa98f987162931527e9f9bc;
assign Ibfacfe5b83819afe7fbd4bffa2d6d4e2             = Icfba3f165f1cdf2e6070239100e9ac3d;
assign I2d9d14b5c585e74db793171f304e5d61 = Ia4e89e99acb95f4183474b94798ca35d;
assign Ieba89aa901e61218074af53a2484a74b             = I93c51f71db0e3df7f6e2978fd93fbb54;
assign I1e7165374d01b2b7abb1e1883daa4463 = Ic1927bb3335f6a28c0816eba12d3975e;
assign Ie0ee5445c56a5f9b41640b57422206de             = Ib7410e44d23eea21613074695b64bd2b;
assign I783fdf0d5058b09d9d0d5c87d9926c50 = I5b8a1e1a6b904b0f6822c224ee0486e3;
assign Iacbb4daf5ce5c7eb1a2afe30d0cb5382             = I93cc273684a376d76a2e3468b3dc8bd7;
assign I1c66ca0e94ab96e8420e97641a5a707b = I8be4711146486fea913843e497065b50;
assign If08370fd0e8af818c6db20f43e74034d             = Id133dc3fa65840136b1157fe97a1e962;
assign If5f2d3751eb3af97e20c680475976bb6 = If4c36727ab1c29bf78f72e8acfc00d7c;
assign I8b3b875c6c07bd97ba598a5139156fa4             = Ib792104b6cf946d632f7591f2cd5e104;
assign I96f91ace9649929071ca3e6e87eda861 = I9b096ce09467c10f448496fda13987d2;
assign I680be647bf2a62e0ee9b5d379dc87b4f             = Ia44bcc8308360d3e6fa351bc108df3fa;
assign I27968f9d2e9dc75bfa55b1e5ad6f8c8e = I57b7b48f13436b19a8d6a47e014eb41f;
assign Icbfbb37bad6344005dd233b3605a784f             = Ib29a26c41a3ba089efd30c3256106a7c;
assign Id53e488ea1a69e9d1e50dc276c14bb43 = I5446c1c323774715371c73bd1be66697;
assign I83330fef69470d2f5def8e6d7d9c50d2             = I8999f385aaf15b67e4c12e56c7dba7cc;
assign I8440ba68619a5a3aad3510ad6ecaaea6 = I6426943b4ab66f17c2b7b399ccc7a6a9;
assign I7b33ddad346077928620344542b9481e             = I202980f6263e3b312c38061224992740;
assign I9e00e6e111b313b2efd5c9d32eae6a8e = I595665d8128bb87ab62741d7ac520a4b;
assign I8d0a1ae4c47edf1f2b99d1175aaa7197             = I1fd9ed3763ff0ce0a671360f83bc3613;
assign I1836b01cfa5570153a8e4387baee29d6 = Ic920452d5997a8477724fa78c86c0fba;
assign Ie5757e7b1647ab7d43cdbcf98cbb77fc             = I4b58194aa6a5b5c825f14bb926a0ae9f;
assign Icad06a6e006badf38d87cd3c4fd0981a = I3a8e9e7d2cd6751e8500a5567cef5acc;
assign I0539d598bbe3d50940329a282c801328             = I706daad77f6a6eddf5576c238fa4714d;
assign I8c061e6f5fb7e2be23d69254f0d0f59c = Ib0dadebad37d9ea9d01350054872863c;
assign I8acc93b34974c1e708b0e1591f7b2d3d             = Ibceceead1cdcf8805e9a9f93b3b783ca;
assign I5411a76d49de45984ac852d98159ef5d = Iddcffa815489773b3688fd68dba18bd8;
assign I11d967a5c5d14c88b5587d4cfed1d05f             = Ia5956c899daaaa0b2b0c16f524feaf98;
assign I826369ad5207f64f64ff58abdb9f321e = Ife0952b85f14a960007b67646b0cd969;
assign I6da2b3a481ee71b85f3087b36b399288             = I7f353333180ccbf6a271c9745430b199;
assign I4c266cd72fd1cd92f21511071a51c361 = I4d54dd2ee2f32909098d3cc2b6689220;
assign I280e20c20c0b4f26278b3de9b2ff84e4             = I958f0106e3ffe429d0450f4b6e9ada3d;
assign I76aac239cb31a0bdcebd7a3e3829f274 = I797c9cb725f88c07be28f017871d17f8;
assign I544f6263f16cd5e0b7cf28c511a8f6e3             = Idf02454b4aacb6ff03288bb19a4771b1;
assign Ief0092617ed13bebb791c57c0da0b12e = Ie165d0729542c81ca89f45d15e0afd3d;
assign Ie11da10808c4ca84f399535df6261307             = I42f39cecfe5c3d77b3fffb624cdb2c0b;
assign If1a6e0ead8f7aec9046bf22a1f59cf68 = Id00642563679fa9a6696f8e7bbdf6576;
assign I27458d76b3ac6520fb379405c6b2956f             = Id7b0871cafd2630ba4dfc3e058613908;
assign I26ee3d378528d4a8469eee34a7b5652e = I258c45897919cec5c6acaddee7f3a41b;
assign I508bbade361787127e1a2e8687ec884c             = I18c1c4d71799c5da8172f6cc63d2d37f;
assign Ic8f3b5e177f927b64f1213625abc76c2 = I1e11f0088959aa40b4ad1a047b59caf4;
assign Ic19486b6ab0373b9c0ad8f7597782d8f             = I7d53f3ce487b0a2446d5205868c29175;
assign Ia813a2600edc508e2eb59a9856e8fc4f = Idce46f6d03376bea1ba361e8c59f8bd1;
assign Ib8e68a77ad8b9e7cf415bee17645c3f9             = I37fb9120bfe27a0e7449583dda735479;
assign Id04ad2fc64d6c346ae479abcbf3df41a = If17c0096ce34b88007247bf4c429d5c4;
assign Ie84be0ae8311d906eff08f7f5b214943             = Ie7e15e6743a750cbf1b272da694b47dd;
assign I2827f1757a4ffc394869610f710291c4 = Ifda1c55899cd3506853cc82b450b3936;
assign I2525111a2fb5f10d64bbd16e148653b8             = I66a1e62b25bce18e36d78c382b40b1df;
assign Ic8c6fbb1e7408869e5d11d0aea83203b = Ic69094123b75ae36e3e54f179a9f2cb5;
assign I691c84d81c60a462e28e2b2bae3ea845             = I9b81ec12daf51cb61f7dc0b9ad01cc1d;
assign Ibe0134da146c0c96af213013c5215943 = Id182a776b03f48fb139c28194ae7ab6b;
assign I4904ab14b19fa1b6befc218bc7be3842             = I9d76cb6c99a69086774f7fd471dadf53;
assign I46a2e76ccab8ae201f78845054028074 = I65171c9ee8449407484e5c82d13c6751;
assign I0ff382edfc8051459657ffa3899f5f73             = I4c59798356c8e05f8b2cdb4e202fc4bb;
assign I1ee771cad3766a589cd62746062401c4 = I92eb6f60c14ee9eecb01718b01ea980f;
assign I8f94dbafaac589ac9f14b56d4556ff96             = I395b43b11730131a5f4331b2ce82717d;
assign Ic37d0375083a9415f7c0e9650ef0ecb7 = Ib5d1a7cdbcba0b654c12063d4f1768e1;
assign I7b7cbcd1c6d2a2eeaaff474536a69eed             = Ib3f07793c2e2cf7b6ac988be01a55829;
assign I73167dd9e24b49f6af3f7493cc2f9c0f = I07abbbd75d91018ac53f53e64cffafb9;
assign I58dc9cce6384160c0a85c6efb3319cdb             = I05ad19dc723fe482f93cb524c8c86cf6;
assign I156970479a68c248bffd30be0097ff8f = I4cdc955fa9afc75c2c977de4ec540e1e;
assign Icde3e6dbcf985682041f30903ad95572             = I1db8d47c1852578aa6325919279419b1;
assign I851f4bdd95d1297f7ff05f01830c93fe = Ie79ce8adeef2c3c24a3386f054d0cf5b;
assign I644ee0055a55f54ab3544bb532e39c61             = I98ec1bdbb599febfcdc06dbf807ab781;
assign If6f8ef7f0cc4860dfb264b645ab0898f = Ifc2963762403a00c4f3662b2863c991e;
assign Ic90b98708faa8c8b75d4bd9a52c292f7             = I86f73b27c90bbd800b521fb8953d5506;
assign I5b983a4c1b35218893ed1bb0aaae26c8 = I5e8ed024e2f2548bb375a2ecf1918a5f;
assign Id2a7f0781d18dccc7c4e0b383b7cddfa             = Id117870de7302febd51da982ab8b524e;
assign Ifd281eb29091bcaf3a2929983366e637 = I256050251d23250854ff337bef28e460;
assign I734e601f5f9d568a44a48834559e04db             = I6cff1d82f4c1bf7789e39b964dd9e6fe;
assign I5ef5030a4e29e5e3c981d2616cae1ccd = I20ffba20af04b99954bf719589e90d1a;
assign I749e987266a20840bb8a4b1a2a2fc5b0             = I5d9786c9b4566669e7981654c3c10da7;
assign I3051150debf8f223b936ea5f169623f8 = I7353ebf3a1cde89d2bb3fa667f7f5485;
assign I9d2864024148337277523ef7fa2e1600             = I83dd9071e7e35d7165d556a67d2d1658;
assign I9b76f1b49c0faf3f89256a1fe04c4597 = I97e82e5f6775d1e31537b891597223bd;
assign I754563caea429d3d0e22df5d193b84eb             = Id62c5db9d4a4e5eb91ca4b6876d36a9d;
assign I62626dac5bf648ffad6e6e3cd836ab9c = Id25deba967318f049de8163e67262f4b;
assign If8bc141d98ebe1be7fa81cde5c65868e             = Ibeb5414f37bbb8176c1a9ac51957dba0;
assign Ic527dbbf40cb847b5e5400f177a635da = If876ca6a14ffb4323503ed46666bc25f;
assign I11094e852295755925c3c61f1df81643             = If40561e9d6ab97e7dc2c6eca6d0725d8;
assign I44683db6537a0ae1bfdca8b6448c3772 = I5109afc4dc91780e05704ea5e1399e3e;
assign Ic419255414995e7168afb97b051fa64f             = I630618151200231dda94b3fb59a24829;
assign I5a03f223dea2bc87a454b29c3fe6058b = I621b20d29d3a9a9f41065bc3c3bbd2d8;
assign I202f88fdc946494d55fc8831c2e8a34c             = I45948c2ccae2bd2c2fcfe9c75787e2b4;
assign I8a7824d737ac024ffd25428f6599c070 = I76fd9005abd511c3c5bf6c77de8bf2f3;
assign Ib60d4ac0fcadcdfce5a14fb92f58423f             = I73048e349b470dbb16b2b3e69aebcb3f;
assign Ia7e5724b4f05b0b6bdedaf264e797855 = I925f6b549a25cdc8f85152eb21ea3b58;
assign I8645e1326c66f5efef4b9c923599d1a3             = Ic3a706eeb522f64147d4946983a9fcb4;
assign Ic8d1cb210627d8d6e717625ad3dd0fbe = Ib42d37576e3aff3d205f1f8822cc58b5;
assign I2afeb2a7b199c0c6738938f156ae4274             = Id8934e8818877e81d701105823366043;
assign I313adb9858a6a31cce5af3d108459bb8 = I3ce10718a2211184999663c3c2493cc1;
assign I7992ea31927b4f0e268462a3b0f18c5d             = Id5fd5653bfa014fa0e956ef4b1d83291;
assign I36dd39ffe6e62b2518e12bb8e544ac20 = I06b48093d4c9b0327c3efc6fa4ca7daf;
assign I484545c4d2c869d79eb17f51e11070a3             = I41821f6b5a613fde6539e41a6a0c7b65;
assign I94337aa2c4ca0ec7a962962780f21f11 = Ie8e29053f122a9247b0dec291c6ef4f3;
assign I280fa9d114e227cd649bf0e55e845651             = Ie8d437ed136f7f5971638d1f62ffdf15;
assign Ib2443922534953e49e1af5343c028fc6 = I9b49e1acb81ef5b088b808d2e4ce9954;
assign I0426ef66185128dd1ef4dbb68dcda585             = Iaf46eedc430b55905d73486ac0752c8f;
assign I08d6c121fbd306f3908a88ce10779ac5 = I364ed3f83c49626bc3b939e53524d9c7;
assign I7a2e554d07bbea291f2cfc18694fca3a             = I32671ef3896bd0b586f13c092dd04b9e;
assign I1b947b03d2db27afe8faf78f580c90aa = I8188dd7cb03854c6f709de06ff785d91;
assign Iace8b3b3a4c16763132b5aaa6b24212d             = Ie8bfdf207d647c9f161bdf265a8472b4;
assign I05b4915602c4c635f9e91ff69432ebf2 = Ie7cfdd25541414ff3f8d6e5d7677fbe5;
assign Ib2f5f5fc77ea8b529f2471c54388f2d1             = Id44fe933294cafff88d133a0ddc1a832;
assign Ifdd87b92e70f345ca64fa4e96d732210 = I6386a4dd26e7c36165dc265b3a2c93cf;
assign Iddd954df5bae9b4240e0512f746669a9             = I20c1f8e56a14db0665160ecbb277fb1a;
assign I67335037a5b54e1b5bb316cd3519e790 = Ia659126b51468cfef48c97a135a71500;
assign Ie5f8620371236cb11c9e88c16b509ee8             = I7627f96e870f6a3e8abd7ac494bc178c;
assign Ic0feb7035ff8f8962a79aa20f4129bbe = I866b30a63b3b5fb708934a1cbb0e1d9a;
assign Idf600b93ee1018ecf969ed7944b6bc7b             = Ia2d3997dce108f85ed64e88780e99efa;
assign If11c3d720e491cfc18684f3a23f6b93b = I2b7822d5d77aaed61eee87570564df76;
assign I7f90f96c0260560ad5e6dc7448b2670a             = I6a25dc88186816258f1237123ee4968f;
assign I5d4a36427e26532bca590796e4107dcc = Ia20709f08cfff3a51d4af1e81d640400;
assign I29e940970d87e8e09b26ab1b0b8f2286             = Ia9d61848b5384a8cc63321201174f3d3;
assign Ib0eb8c6ddbbcd4825e8fc5b1c55495b3 = If1c0a3726041f70e508d68cbf6e40e04;
assign If4d75f83299a21802b6fbe136913489f             = I53ed79856aae53b180f28b47822e89b6;
assign I0d5ab203120026f15a1d563bb65fa1ab = I019e399a1cef87745e025a7d74e94db0;
assign Ibba4e82d1510ddc16eb4ef64893cec02             = I76503bcb779e039edc9acfc03a2d1ee6;
assign I35ca485dc9ef601029877a4ee46ed942 = I0dccb8eaad52ce4d780696a8485420f1;
assign I108c269ceec4adcff9afeda01101b838             = I18ae85d6725cf0ab3b69bedeef651425;
assign I8c1c4b4851ed06bce6af5b392c75c6b8 = I1ff042bdb52aac5d69791e96e2f9706c;
assign I488f6d9676aa85a55d030bf12e8997a7             = Iaa3bbfc6704e70a55b8e1083c326820f;
assign I00fc4e266ce9e790501c78809bfae38e = Ice1ce5b4c30841dd92268559ebadafcf;
assign I5395ee57418c31e11cf847f0f514ec19             = I8c1c3ee4b57d56ab362672dfeb4e0ae9;
assign I35fa53ff8ca5fab19b6de45beda84ff2 = I3d149293f106ae8680c7f4702daa0bd6;
assign Ie9b9221b2122087cd5f309570b6d31ca             = Ic8e0765b1cf95f2578a7ec656d027f6e;
assign If3c4067202f592fabf77cd76db5575dd = Id17ada8dae3f9810d1892d34f2288859;
assign I4eadce87f47df6d8f0e4acd057de5a09             = I39eaefaae486119c8741c5e9b7f85bd3;
assign I64276a920c9ccf7576c15618812fd152 = Iaa2cbf59f6f61198b4fcf5a741cd5bc8;
assign I99d761b75ade1fb2e8afbb1a77752609             = I6ac8d8000e434fcca222525ac00f9849;
assign I478a999d16ad8a5266769d1b8caa79db = I3eeeb1949945032d6c1759875426b733;
assign Iff125392fa39afebae1637a19c4e23ec             = I114cfd3fe8f5db92b879e0dce592af3b;
assign I29f2854aec43820204ceb8f3eceed6c9 = If2dfcbf493b761fb5d7c622e739b23f3;
assign I9c633aa620cca127b0ff8cf882178e76             = I8db1c7f6b5c7c04f71e7fcc18f7b9941;
assign Idf664119a34b4692c0cfaa4c742480f4 = I3f5053e519a928640ae49cf4e5b39d1e;
assign I4e08021c0235fafb60200aab97827a8f             = I89e516738a408ccbd495e4f5aeeb38a6;
assign Iae32c64d9bf268ccacaec2d40efe70f4 = I01c94743a11042e75638ba6618356203;
assign Iac4e3d20178049f9c59abf374752dccc             = I0c02b9318bc4f50969f8d486e587a627;
assign If30e09a7c080fd91758eacb33912b8d6 = Ic2b000c3b2ca3beff2d427caab04701a;
assign I3e59b2419c7dd1553b792d536208514e             = I79224b17e2d1f87175f3118287351e0e;
assign If000ebe4f2ddbec4afb6c0e41abb2f9c = I1c2ee281cd47a8414851c5e1c758ea65;
assign I86255756ddd1f88b74e070b19f8c3bfa             = I41ee2f859df1db26618ab9c2c0a57be5;
assign I714abef2427918d8967e5fff40fd48d7 = Ia3ef2f70c5abaa852586a33c505aee0d;
assign I91a6408a11fab36a8ba3dbd3f895a803             = I15a667ea371ed0fd464f42fb9ef61766;
assign I6229267ae259aa8193a90596f8c1d432 = I0a0340a0e52145f3597accfe4a4e8624;
assign I618d33f26badabfa578908903a613bce             = I25c2d3dd7fedd28f0be0e3d8dccddff8;
assign Iaa26fea88e8b3f2ce1d402b48c7a9eff = I3c3c22bf63e55a81ae91b1dd1ef615a0;
assign I8d7c1fe2e33bbd45379b0325a3c5e989             = If22b31d70158d864ca6b0201ffc2b7c3;
assign Idc0f6e44fa41f76f3ddff9628d25c005 = Ib02268d5048c7c8e83118070e927453f;
assign I56bf74b5890ec67090f499afdc0a9c88             = I7950b8505327240095538f60d81834d1;
assign I7c14c6e871660c6c830de981c07f6b2d = I30be0b18e4415ca50f2d8149efaaafe6;
assign I739267bcc50c54b8a685cb3c6afc5cc1             = Ib75297152c09323c7a6f674c93edc01f;
assign Idc5ee83aa6a50531e6de2d9abaa26843 = I3bb4d24caaa0882a75125e466070f0b1;
assign I822d7973afe090b2764335f1b72dfd0e             = Ie813deeac800a6b251209a1c8e2adb12;
assign Ie0ff06499371f17cb8c56c9f0c7ee666 = Iaf36ce8598a29573979c683a5e2cf9fd;
assign Ibddfda6413e3dd2f483c3174ea836b6a             = Iada283b3152a5316b6c7077292ac0a29;
assign I59976ed14d4be22603d2d164399389f9 = I82f0e5a32d1bcd761a74f1f9ce8c88ba;
assign Ie421da1dc5aaea57c50d0c7d9c5a2717             = Ic14e12a907c5d6b7ad2615905a64886d;
assign I9e94cdbd4a445883fb45fb3ed1b05d7b = I659322a9fd0d5eac514437b02e0491b3;
assign Iebf769a6bdaf214c1006c55c608d4eda             = Ife78b0889c9c7129a3000cca66ae4aa2;
assign I581b4fe258cb92d51ffc1482da718625 = I44ead0ab5ccc53226fccc03024643771;
assign I12c1035353e553b3b6a13bb174ce6020             = Id926d49513e089a52b17978a9ab84372;
assign I19f794db275b2266dd9a91b3b0174329 = Idc2a9c6dd8d2aa912548c918c8a488f4;
assign Ibaf2f1f8bda2f6b932dc30f8369c0e1f             = I4dfbf2a2c01ce39fea9b756f9b106fc2;
assign I7d4b8ac371172cf90b31890df5693875 = I08f22261d5713c0636d77c7938f592d6;
assign I88a61cf72347d695489909d0819332ab             = Iad7cce628396ce9ffac3ba9dde7ac494;
assign I1f02219120214ac3e5f5279031facc56 = I04c734eb876aa722e84d6b9edd297978;
assign I39289e6385a9bc378a9b8dd440249a7f             = Ib71f9f92515c200bd16591c656d69ee7;
assign I569a8645fa9f5476d122bccc7f40fd75 = Iaded125f7fd5c833e7206dd7071069be;
assign Ia6d61947d36fc128c689808c82db80f6             = I8e39b301e04135b8ab88d54e7c1e22f7;
assign Ie620ab2c461442bf7c7ddd962dd65839 = I98febac90cccb5fc1f3d966b6e38c4d3;
assign Ief5cbddfbfb98fce4812a676849b9a98             = Idadba73fb37b81563818e82af3d89a58;
assign I3dc4a3e2c52f2f74aaf1e640543fcecb = I0038305f94aaefe2cd1a243580d95932;
assign I3ca2b9b77ed8d78a10aff42a07a53b07             = Ic19accaf42ef2b61fb52ab3621622ef2;
assign I749c798e403cefc3782b3a63de02e227 = I0d41bef808860bde56d48792764612d5;
assign Ic5467e42aa377c6ffd8f70673808774f             = I94f508ac67f07b73b3ff1d5aa5955eea;
assign I3ce1a50aa7de5d1dae422eed03c450b2 = I373be7c3f9511a2906584e33e5048abf;
assign Ie9b042f686381739b9ff219041f1e0ce             = Ieb8588293562c9c25897044b9e5ed6a4;
assign Id9474b1f0f1ab396654b7048eea873c2 = I2c8f4a147b363d9c5ef0e080d9a9ed40;
assign I694d471fd353eb54aae08a2afa7b645a             = I671d71d9ca760cc759b96bbacd361f90;
assign Ib7d69d239aac1a9de86e2f2f1337c5f6 = I9171019227f35760d02d0c8ce786f4d3;
assign I15fafe2baba4d2f28037023a81ce0a81             = I3f793de7fcfd045af3970e4ec219128b;
assign I40a799391b45437a24bf9c7cbc2ec409 = I669d34b955d2991ebbb31c149ad1b6f8;
assign I1c85a2d1df6749a194072eb731506bfe             = Id49f950b3679093b10f8b64ae89c5558;
assign Id81eae2229fec7726aa687d711d1b998 = Ie0b5f51835ebdb508a596eeebf0e4847;
assign I0c4268c01aed70ce4fc71531bf4bb862             = Ib70c7567e552969a2757c1f48a2468ef;
assign I7bab2b945804593835eb8b63143a3345 = Ie644d131c4f2c603e8e64c5581fdf822;
assign I7d4924388dc5373ad7936dca76797473             = I6dbd0c3ac9f2b3887d87e316b8b40b55;
assign I4e7f07fa261e44488cb5b0903d2e8c5d = Ib70e99c3acc76286a6811bcacc9284de;
assign Ifa43d74fa91b7b9884969f575ef9ca8e             = I8c309d7fe6aaa8c996e39b8f3dfafef6;
assign I5d69471b78cf5aba461a12cfe6d7d11e = I263aad78110a1136eb7012c6983b2a8d;
assign I3ee10f6a7785a236db317515fdd23a2d             = Iefdfd7b1924f8b6049b02576f9948027;
assign Iba0af171e17c12093f5dbde019fff4da = Iddb75e0197b9a76b36a59ac2a7ccdf3a;
assign Ia34e42f8de91fa4861b0c6cac5dcfc29             = I2c14ee79492962576e12ff1698ac0fe1;
assign I580c7b678e4f2c08a4d521c335392c07 = I8e873fb2321eea82bb590a92411e2e2c;
assign I46894c6526983bf1ce4b503159131b41             = I56e90395afb09c7d775111d19856da1d;
assign I8016fc36bc9614afef570a084942081e = I6cde57127c5bd2732e71ecb7738fad6d;
assign Icb82c9ff4cb58159a1c3115c6fdd5f8c             = I90f0c524f6b98c28d18db952ac40c83e;
assign I744066a189658aad33b32468934ca485 = Iae6ed7748692f2edf1aa9d73380075f0;
assign I3ec5819176ad4b0895a9118d90ab22b5             = Id50649fc4e9de24fdd9f06499a733b87;
assign Ic2a5d82d3e19ff84f46d2d71b3d544eb = I08c03198b9599b2f4590e3022e398f7c;
assign Ib7c5850b4f7cc77be2048d114a2128d9             = Ifc988e99b4c4c1ba2d5cf3a76695900d;
assign I935a700d902a104974a961beca5ac99a = Ia62832d325f86160285c4d1a790a32cb;
assign I4fbdc4ee57a3be42b62d9bd43078d6ef             = I53c579c64f0d911fe3fbc43dc3e981de;
assign I902f91dfb3bada8a106f46923239c93a = I2f23d4cdb6f5f827513aa60266936e4f;
assign Ib3367565e4456da15e7c2315dccdb5e4             = Id729d27d6424495fdb4deb2ffc038f01;
assign I4d4f46a02cffbf72298704e8a0504fe2 = I4b99891bed4f5c149cd4a5b4f1dde0f0;
assign I4accbad1b451ed2b622e15ef9ae16d13             = I8816c4edb8c7f5fd6e7a3c81013116ce;
assign Ie8fd35237928694738b464d52847c2b6 = Ia4f3cff223e24815ee1d86bf41756f06;
assign I32bb50faa2b246b2d3b462a79be597c5             = I88ba486c5bca54f6c120a654b81e0a90;
assign Ib73fc8722db87e7be4b14ce361b79719 = Ice82cfe55a5f226746e59e5c8beb46be;
assign I33bddb0adcc2af7b12a83bf843036385             = Ie1ba6d92c19ebbc5c994d9da3881f6c9;
assign Ifde9664e13fe94aca97da5824ef0c08e = I09031235f61238b0e32ff52641aab70e;
assign I2c926fd9d306e9ae13364e07c4b0395b             = I023278cb7d70d4608259e10c89e97117;
assign I3d25580e525216c23557ffa5ed998bab = I9d7614d286377329eb3999213889b707;
assign I8e517c401d62dbb10dcc96ab536f6afb             = Ib8c744194310bd59e983e392b828e9b4;
assign Ia3d21a8d9a8c24b112965d6eb966de8c = I56592e1452c4b559af19465b30230ec0;
assign Idc6d40a49f05c5422758cee50f787eb1             = Iaa2aba39e0454008fbeff8f9aa87a481;
assign I7d7923beddaf4b873ae819914599f02f = I384d5377ee6b8f7eb2db23a2e444ddbc;
assign Ia6308e16fae5428f4ab6560f5b21479a             = I61a43aad15d7a9943f74617f434af306;
assign Idc6a066b872fa91ce73e9aa21d668e83 = I477a920e2326828bf026b0a6b6a18e2b;
assign I448f126fd3932d5065abbe7bb2d92c56             = Ibd8114af3027bd3364395e7b94484272;
assign I5ea37c7893e55ef146fb831d8c09e87f = I5196382b75d16892d550f17893de15ec;
assign I960768a84aec9d5b8bc7c1c523024a25             = I49167fd9caea095581855b45b1f85d49;
assign Ic38315ea78c667a1f77a5fe34ac62412 = I213ce488e5345fa405a9c5df297d6f74;
assign Ide1d7dc22a4b271ef764df14ac22366a             = Ic502f151ee9ee01786e216d90a29403b;
assign I2b954aae3ff5e2a0ce92a55107a86a46 = I5ad7eb9d3ce7c712515254f892d1670d;
assign Id9364a29fd79b52d0442e18dc0227854             = I25f89c7f7f11c7e2811913d6254dbc8c;
assign I958138e39e14c8fc1de83d02091b8f6e = I914dedc1d5e5e21c9b8d07ec0ecc01f9;
assign I2b2bd845428c49346ef8e94e95b618f8             = I3f939889c013f740cc63c981d2ff85b2;
assign Idfd5a9e4c4cbd4ba9828220a7d021d28 = Iefac1e428116a797c2c0803410ac5601;
assign I7ace6778ac86b3e05939a3fcc716136f             = Ib0d2fc4f353a82d37bec9aa19a80475e;
assign Ied5041c527b4f04647dc80932b9ce7c4 = Ib534288c2cf976b6ec85db743bc2a823;
assign Id113cab2dd1949d32e3c1c15273185c8             = I2f19b77e5bb1b22b3cf5b1ace31ee6af;
assign If6488c8e84e69a99816842a90c9578c2 = I90023493600924a76d2192080cf6194e;
assign I103f1449c78c47396d6a54dc1c810934             = I283f82fd4a9700daca6ff1d16f747a09;
assign Ic65f12c4a71f8c3af75f426128b333f9 = I8b419d5827e5b1af9649d602401c189a;
assign I044e01e8d2df46e03f00a0af2beb0bf5             = I8dc5483fb01a06ad8650e5fd4df30f49;
assign Ica6cd8bf97c702ae2541f682cc418a80 = I485f9d1104a965d5d035feef912a2ca8;
assign I816704585ad393f685731104ad3ec64f             = I7e3f6b4bff19a0644c12fa4ef3667d84;
assign I73054b5829fd26eb2b09dc585f2c62f8 = I474f6bd977f4197742d0bddb3bece684;
assign I53121a39de0bcba91a4d0438be2ae958             = Idf2371d30bec7ad5dea346a4a48a6e75;
assign I221be7886d94efc9e1ec553acd79dba4 = Ie989550c9101de382056dd60d5da0e01;
assign I45a7ddcda2662e36b7617dfe64514346             = Ifd5a3069363cfc42e5a436856eeee708;
assign I33557b5dddc36fe3625bf64e016c1c7e = I9b76f0121a3f7e887e7121db50024ab4;
assign Ie317e5ea2ca4ba2060d0f491290af96f             = I1a4e12577ac5e87d40bdcb54fe55818b;
assign Ica7d3d482ec7dde7081b68988f76c9b4 = Ic3fb524ab434e80b3289c9241b65d224;
assign I58703e8b6d04f8c69ac38f5fcfdc4efc             = I1f1b6c20910c4f14999da6c9fdb4c349;
assign Ibf9561c2c5242296a3b607627e7e7989 = I259010e323e1e8dcd9dd719091131f6c;
assign Idada779a1ac7b844867571d77054b657             = I1b0a200eea98f075f059d2a26b00f833;
assign Id0d621bef47b5c5735a4a999611a1c4a = I30d615203b697787ead37394953925cc;
assign I5ea02b5349cd4d99ccbcb6b26f0cfdd7             = Ie0dded072843efc1613cfe7136af37da;
assign I33cee0fcc65354655c9e57b3d43c11f2 = Ic9146d8b3dd0c612073b70b8a8791e8c;
assign I30b0b1d54912c1a41a02a25ab238bb54             = Ia6d6a867ebe63a8926d9affa4c15e376;
assign I8baad814c6bbc783645f574455b0f2d3 = I3e0b41bee4c76eb5f3340ad23bfa01ad;
assign Iee6da3120d73373627b25ab7c0dedd28             = Iddfc447b0c96056ae6e6434799ea00e9;
assign Ib23a7e23bc223c7f3e83661811493229 = I389ac86954fd70464c9550e3fed4ed33;
assign Ieeba01b18a244ab8c0ac263c138fabcc             = I36d03daaaaa37229d462f4bf5e521f73;
assign I55e8b1c375d49a1a1f044a4a60073d60 = If4cb744ee52b6ae793431cd038069b57;
assign I6404d0df952b5bf8292c753e4c6f35d8             = I91e49319831eeee5dc75eac77ed8f8a3;
assign I023853b98208afd9bcb1ff63abb91b2e = Ic3cb34aae74c5f1a870b3635f8a40764;
assign I913d818403024510c55b65b56a38dd89             = I4e9f03752b041491ae2bc40fbd2b8d43;
assign Icd656c959fe941e863db11f02d3c514e = I877e8d94236c3d8b0a31858a98fba5d6;
assign Iadf927d18644a232ad1f1eba7db82934             = I9a71e50dac7ad707a4b0946ebc1fe6d4;
assign I06cea262d84c35f3e6a1b6690b82cbf8 = I77371f0e55b4684d1af196ed52d3d997;
assign Ie4c9797a955778694dd8615219cb51e7             = I8220d15825d6bac07d773ff0db2f9795;
assign I1d7bbe81db5320829eb5b29252fc6cf2 = I83c7d177eec2dad0a924557cdc91ba77;
assign I5510b88bfd65811b3200adf4ef975b48             = I6b2dc98acc78a1151dd6670ed981d839;
assign Iafad27be14640dbdcff055b7e34f6467 = Ib1073489d63ea33d7f3892f4ff875358;
assign I7774313f1ae5a2de98855aad572b3676             = Ie371be4323965591a5786063ba028ce1;
assign Idfd58540bb8d1465514c3c843d303825 = Ieefbb5d6f4ac1e586832c5c0f513c5a2;
assign I46ee30b46020d91707689f3468f00e26             = Ic4985251ed9f9120d2232ec96949831b;
assign I7c98a5f1ea935e4de159795b5dd795ed = I5a21996f5724a2a49fcf8e928c01b062;
assign I28a5ed4c239e64c76bb6e566b50cfd23             = I6015d64c067415fe216d90a5be409e33;
assign I84b1e71a64cd4d96c44444e337dde784 = Iea1297491d1dfe98f395d8c73808a893;
assign I529f92b82248efe2cf64f7da0ec8283c             = If6f304fe091216273270713c6b6e8a6d;
assign I609aef4d51d5d190deea41f71ef0403c = Ie9236599cea94cfb603c6b977fdbb44a;
assign I7846bc2cc11e08d05f7c853c4920d555             = I779ee6daefe3c5c96548dc5e0ba83bd3;
assign I68a99adfa01586d1ad7bdeb282f11d87 = If8fe5af7e5c3c97b5a713f6bcf919f1f;
assign I7607af5d98e8070e3d15cee23cdf877e             = Ieef21b505cc215387f8930888062b767;
assign I1f68aed9a1379bbbd2c531fc0df392fe = Id46108963921efa50aff64d4dd7d1701;
assign I79a705ee1e414fe4a5fb14e9b3ce9597             = Icbabacaecbbac74901402e5e5874328b;
assign Ib1cbee37b3fad49ab5805647ccf95b7b = Ife25829fb3c5023b7d69bbaadf9cf77e;
assign Ica3a41ace27f7d94377981079952f4f7             = I6ec13a161f7f1a0f57e9ba4998474954;
assign Ibbe9c1e2c9f2c0b00e4be25205a824d6 = I3375fff5ee0d4b4b12c5a70fbdee59fe;
assign Ib730fdb59198f23d1e590f6d6039e96a             = I71f9823e92c51be2e9a050d01e63902d;
assign I6c7e0e56cd76e03261638e924f90377e = I68c35d63dc95baff41b4dc27a86d2342;
assign I31243de90dc2a1656ca9d5e03bdd78da             = Ia0037030d79400734732f061fd81edf6;
assign I676d7f8a89fbbef4b067d07264ae427c = I8da50e5093acefb6f809aed64564a53e;
assign I04f90a907f10a7fa1ae3591b48094d5c             = Id796584e3e7af67536a27f7299b71916;
assign Ifcaf093fbbec17632ca0050583df41c4 = If988b82b86db1f4ff6d3695f7b0197e4;
assign Icfe1a689e33b2b9aa9dba692d6d610b9             = Iec938bc1bbad930fade05d74c10989a3;
assign Ia358ae5a96e63f3bb5c6bb34f263c387 = Ia9f5ce4603af279bbd9b486b67016482;
assign I56b3a97dc3037f0bb2eed93a9482c813             = I2a7a7c5eabd1623c1c3d4bd93bf18617;
assign Ib1e4443484bfc289563a8b7d9b1c86b6 = I0c5539373b3868d0664a92157b4b4226;
assign I282d2eb4e74e034694e33273b9cb19d5             = I71cfc7fd85636c5554b9fe9f9ba8e3aa;
assign Ib3baee13e51f9fb8c39d04211497e274 = I03b0694777d0160a83cbc82ac1397736;
assign I31d25b1b49e65216e90b39aa27acd6be             = I4c8ae97548bc3dbf3e3621f80c3e0835;
assign Ic24de5d8c9148fab7b9dcac9d8996740 = I10fca5f2cbf5e2bc3433c0dda579a051;
assign I85d95015a9ce27a18ccbf73bbbcdbd70             = Iaa93c760705c984a0eea90d41a6c049b;
assign I46489795c1a8e178f1b2d40711655c44 = Iaa1e981134f5a5c02983c49562683bc5;
assign Iff7950f24f0a6b0073942c37fff49d37             = I2acc73851f8a803e69c0f1865e00f46e;
assign If39c47fd6b6913ec7946018145d31945 = I6eea5fde8e2517554ad6ba25018572dc;
assign I6072331f838d82329a07a4ffa340c7b6             = I928333e9cc75d49fa6f7094e49631123;
assign Ie336a92376f51b145c60f935b8fd0f8c = I85c2bffb93569d9fe1b1bcb10b98bcac;
assign I1f6540c5f037d861dee2c0091cba01ec             = Idf02dd4b7e8a6958913e6180fec1feee;
assign Ia6f981e46e3d7ead096d73154e97dca9 = I9eaf4e9ebe07717503ff69b51f0e1905;
assign I56ea52c50a188ec47e48740839a031c9             = Ib30cc7931858974728d92eb68890449f;
assign If7593819b136ad3db74d793e5a0f18c3 = I23c8b64e433af0bd00cef44e38df99f8;
assign Ie1f41720e296ced1b74cb325b666d88f             = Ia504dbcee6e5894fed83371bf70b2d44;
assign I0b480fa6fe571ea7d25d13f8f1ba26da = I7bfb4c5d9e22d1bd8811844d9c74dff8;
assign Ib3a0307176d424a4733720416d71069d             = I32b4e50b8acefe1c108d777da565f4ed;
assign I66ab48b076a0e2006d1f4741e15f3c36 = Id00274c88b93867a80606343add1cdab;
assign I9632bb500b7faaaaeb649d74c21cbe8c             = If9fd1d8c0c13042a6f2d258478b63925;
assign I9e397fd8cfd4ee1b9cd3cccbd4c03005 = I7741e239c16828889d488cc87647c154;
assign I8522c402e654d007abffcb0e904af5e6             = Iccb437017198e4421ab51d74aed779f0;
assign I177684367c872f5a3df89c0d2bb95434 = Ic828cdd5dfde844df4c150921af2a443;
assign I2605f078c1a9006c93855a9a2b0cf6b9             = Id10bf2bf52a8f1be9eeafcefd6dd5dcb;
assign Icdb37cf629ec16db879e288eba5ef9a9 = I61e829cbf7d6c0ef8ddc11677981e2cf;
assign Idd0217a35c3adc8abc7bb581a5df7a2d             = Ie590c921147b7252d2605f7712dfe437;
assign I225d035b7f8d13e9895ca60f3da8bf90 = I7050adb9d06f767549b7f35c4679e391;
assign Ib57ef2f577cca54713c16717cbbd1ce9             = I178ed883c28bbf3e1ab05cb95f62b343;
assign Ia3572b856ec1a14e316444c2f15ac9a5 = Idc5fb0f3a04ab32948e249e088a11b11;
assign I2e11a697d7f17ac30302eadb500de72d             = I01971a175615a422d264805252f91f3b;
assign I2c927c7ee3628a78f48c6099d2036959 = I9e8ae2aed048068b01b3bd46f30baae8;
assign Ic05b46168884322644db4e331d37d759             = Ie770c4567f35b40c46ccbda059e6d3a8;
assign I578551b6331fffa97a6d05652e406e3f = If43dd31198c8a0da6fabd194cf13bb70;
assign I2f34af0036985cd94ade9cc905bec065             = I25975702f0b9c0baf586fe471676dfea;
assign I6f301798efb2c67ea363df40f2fe340f = Ic0732810fd355d59a3168be896a0f9ac;
assign I56fc99a22960232b305d6e683c66fcc7             = Id2ef737d910326394b68eaa0833bfccb;
assign I744d142b9316b9f8937563c1023882e6 = I7dab71adbe62687846fc027d2789451d;
assign I53c88dc237bb2cd02d50fd7f0a168a48             = I577cd1f9ad512ec10f5008165f2e4a74;
assign Id7fa5f9fb6059439297f246cb228cc02 = Ib16548d471f0a4f4625852ea04335dcc;
assign I21de4f6194dec9e3c401934db92c25e7             = I1de8f87eb39276e073f5804b1df3b67a;
assign I18e9dd5583f3ac91451a4e75f0d5d474 = Iff2f1716cbd73b406d8f07c22dc79fc8;
assign I2a9c673cdd7ded79e09ada38c0f47e6f             = I7f8e7928e6caeac14f787d7e0b6a47df;
assign I64afac5bd1ea7a2ab696e630cc3ad162 = If1295608bd218ed60922a0b95bf1d098;
assign I7450d4ab3ef0227e93a02bfd620d047b             = Ia7048aa3f949b0b2e54ab900efe01131;
assign I0b3bfd6ce482cfb20d461862a0bf8f61 = Ib051eb1091a85f85a1e50007f1b27cab;
assign Ide86f019e9573706c25bd8b4552396a8             = I1fcbb73d165eab038c745fac370fd68f;
assign I16119df9372ce61c0c8600ddba36e607 = Ibdad0ab78e4404c852e60a2b04c3a5f6;
assign I07b417cdcc99eaea3413f563e26ddc73             = Ia822cd52015d599bc45ae7338b4e88e1;
assign I0957a6c9a87bc89dd9748491807837af = I5fdd8e1550feaecd81b82069fe73ed7e;
assign I8eba6f14f42701d22859fbea94bd1871             = I56b85e2d5a7259eb50fa983b92d8b160;
assign I12f8c91d67e31e11033d5b3b266c659b = Ib4ae1cedd09d72c235765a6cd7e91366;
assign I49b64469d298012dbb131d879bff38d6             = I1d23632f8e8f66a30b4ef6c76aae3ece;
assign I690b96154d7717bf62eeb740b10ce6d5 = Idf04e08c120ed116af14a62659675b44;
assign I2b16e5b4e279bb29c3c675b72083e5fe             = Ib578de11f0407cfeb0dac68bd5fbf7a0;
assign I25b3993479d7cc172ba6a480628b9188 = If6a5dc79c0f6ce348956286737a369d8;
assign I5d5701435c96f1078e741921b56e3c65             = I08879fb80c58de5fb2bf547ce013c67f;
assign I7f3a220cdbf5bf1737690e1719f888e5 = I6d4fc81ced37c159303c243af04d345e;
assign I761983331fb6e3c6c437b3f1660f0b6b             = I8f7c4c602b7de5d9a401d3933a7e50a8;
assign I8d068dee7478a9f899c8145ef6d824a5 = Iba1c0ebd9cefeb0dd7f690bdbbbfec58;
assign If7f373506cac70f8ba1222db135c27e8             = I2ab4cc1ef6b743cda8765a22e28fd7a7;
assign I2286af8d6007a7da5c745d75f407b5d9 = I3472ee8c06644490252e606b62bf9bd5;
assign I5ce8b2f633011e89356243a1a71edeb6             = Idc58a89f7d8ee884b198b6e4752ec58f;
assign I214f77e05ac2ce4b94d4c5e53675717d = Ieb7614ad1b1bfed3e2b0089a72fe214a;
assign I70c92e8ada46476d15ef4b3c620d2601             = If9c0f4c64c7648e509077df16c14b7a1;
assign I8fc900d4110bc862ad7287255dddf2f0 = Ia8e304ca12c82e41cb8e4de7be199394;
assign I644e83f0a7d432fba38ffb2d99088eca             = I8cc434418203702ad5a21eb4f0340dc5;
assign If609e068414eed49fbe97f86e2546768 = Ia2c5fe53cb5b318fa63d09881609655f;
assign I73203143fe37933c16fff873c1abf512             = Iee9d96f800fc848f3c4b6b6901a72623;
assign I69177c754e87bc42401bccf54b770358 = Ic124975d36a292816146a2fe61ab3ab9;
assign I039f05d5be891a37e04556f1eae674d2             = I989036e56c9c7386279e83ae83ad4f7d;
assign I3b121702ca62507c2afda1ed93183499 = I3eab1582cc42db0ac7739386cce2a712;
assign I8ad3627f171eadcc960a688ac0afcbc0             = Icf23ca0439c76198fe647a0b785d9503;
assign Id979aeb39d36400b85386a8e96ca5a35 = I589062eca318b25dfe5735da455b6fe1;
assign Ib193b07804d6d5f111b06bda487bfa5f             = I406bddf2c4a4b6e6aedb86d72f14994f;
assign I61ca2dba668792ee6a83850e2f118eb0 = I05721e06a1acdcc0571907c7d853f18c;
assign I51e98035b35a35fdc52f5bab8f19c152             = I5331e97930599788b1df06992c5e4a5c;
assign I7e7f1d73e81031a38992b4f9a3f90717 = I1e93f0470d2818249f1c28ef2a399a0e;
assign Idcada1bfb3c0d1f2a09aab58a2071a57             = I98577e71126ac9bdbe4359101d4d48d7;
assign I029dbf330bab56469b88cbd602e8e16b = I453dd7d7c0a2f003f0b67e909630d641;
assign I94c4e11670b4233fa072517a8f19c901             = I696f551b6f96d0f7d27eb685bd374229;
assign I47ddb6cfe64c5addb3900e193094ac8f = I6387919f2426c283e2d70e471cda54a6;
assign I09b5273bb15d48a7fd78559930fa6d1c             = I1aa256ab19406597846ff353b65224cb;
assign Ibdf7e609b7e42c57450d9d9fdd610881 = If3db87afb3ea184c9e4020c5e45cb161;
assign I885433b0ab16c6d87abe45af13c9e529             = I00f1b24291a0e8496e13fe076e377cb8;
assign Ia096e8920afb814330e53778c955f8b0 = I7979161aa1e2262ebea862004c387697;
assign I5ed85845c39337c37791f16e718069b4             = Ie6f40dc356120aeb6cfa7a3fb5fae8cc;
assign I365fd3d16d984516e33a7b68338d0384 = Iaddc1f2e822fd2fe9d9046d759a82cb4;
assign I1cd93172cf5996bc870063aa642188a2             = I67e23e6286edc4e01a7ebdace62ce56d;
assign I5e86c33e58b50627d7e69a4200525e05 = Ia14bc1fcd5bbdcb60b8e68298f7d716a;
assign I198c055930cb89d0390c336eda8fed4f             = Id2c7c6d20146edcca65120c025e25a0a;
assign I52ef2681091d643e4ed026581feeb3f2 = I04aacd95d9e44657f616e01c9053f0fb;
assign I15943aa74e9fbbaebdc0d54eb6a3bffa             = Ida1e2d8b0e45e14c4c669c8b9d6947f5;
assign I0e30717ed1e983e1c5af25037d5cfca3 = Ia8974083bfd064f2c27dcd421490fcfd;
assign Ifb00ae47340bc99669c71da34cccc59e             = I1fd443d00410d0577eef9f1f26e64700;
assign I640e720e6aaa2f8e14b5dacd51cc6e66 = I268b60cb371b3d46dc3f8b0009f541b1;
assign I688a2c72e69b217d2673e8da75146a83             = I9ea760f08ba7b84fcaad929a3669450d;
assign I81f4ac1f01d8170f427ee5ef89e8bd78 = Ibeb8c72b90b50c6897224ca1a792fa56;
assign Ia1a0d8d7dfd6e877f15cce773f85f5b7             = Ia522420603dbde92a49da297554ede5e;
assign I8319f97640191977a9b89e7639aee739 = Ie232799bd6c4ec99e24c78f3ad798265;
assign Id4451722e8e2393d627dcd0175dc9903             = I9be575cacaafcc13a0306545be56a04d;
assign I21add24f8eed563787b8567fe43947f8 = If2cd93b57cd1c2b91ee7a73a97dd19f2;
assign I3b6fde4ed14cd68af1468ae1d4cc1a22             = Ieb9a03ad2c7c7df356477e8b4224ebd9;
assign I1a772b29d533c44422332cf291d27253 = I0987c561670b7b2b6683303c1be39561;
assign I57d0920119f8901bd4dea2d5f8fb5d90             = If7f263cb2fb7fd35682d44c42639bab6;
assign I8ec002e0ccc2cee9a210b987bf1cccc7 = I3b30b4ab00a49e10a75587aa324d6132;
assign I80a89644e278e96b1cd1c4b7f764dc34             = I5046227e18f800785f8ddfb4a89b1bea;
assign Ia13212b613a21e983b097fe0adbe59ec = Id81305359a07db527e49fda05cd2784f;
assign I5d3df1e7563630311f56143ee6d97a8e             = I73feb8438775bf3faffed6895b6a4638;
assign Ieeddfaf876af8120f779286b4f60f767 = I8b2a79aa4ac88e6b4ca8188a7852022e;
assign Ib57795a63d642a73456324bab41384b6             = I6a423d4e11a97d84120a475db8fabca1;
assign If1912201b852f91e8aa0c73439ca7022 = I6b5645cdde4b35a16fe3e91d90caaa4e;
assign I2370042234b0e93bb66e44b97fca3e43             = I2098616787bd728bc4af6be5ee094bae;
assign I0995a527d1b13090cf68b771d591c041 = Ibc48fabc172f27ebce18d0a9b5120dc5;
assign Ia86740e870d8063f0266b68ad6d7481d             = Id9ef21a12edf48e574256ea34fcde992;
assign I04bb94f5e9927cb7efa70e68658862d3 = Id8292eca087c1a17dc8b5a572a76f21f;
assign I90a7ea789d3bf7f9126c786474a56da0             = I31ab57596896201ff52990b0641b9511;
assign I7594f22f889c391838f987765ad478e7 = I6ef260ef75e47b011a46ba2080ac3684;
assign Ia4b671f3360f3ce55db0dc0e4d78ddbe             = Ib3dd33a163b0c8153edb4fcc90a453f2;
assign I93a25759f720769b941088884bb6db59 = I34e6e9d2153e4a70ee36ab85e72d5318;
assign Id96e744d9b10dcddd1ae0115ea57a76a             = I28496a34b2ee033767fd64f631426b23;
assign Id518694e3b3a268e7168c17250bfab52 = Idf1ecab26889c4adcb835fda6b1cb368;
assign I4d226dd2f0bfcdbea6a2e6a6613c1b64             = I0a4ef7fac369df46d1a4b094d7687645;
assign Ieaf2b41941b840b3ade630e721e6367a = Iddb19725b093506e5e521d8d68dcb8e1;
assign I5029424c9d9fe923eeb858b1e62cd758             = Ie7944f3e2adfac325808f8711c0eedcd;
assign I01a2be56c727d7ca0c5059e8d34919cb = If8572800d5d80cc92dd917b60447b63b;
assign I992e7c551b4aa818606c3465d33eb798             = I58cecb5376f675339028440f0671b0b7;
assign I605682c90ff448b91a2e1a82a3cb0c08 = I3566f2779e860008b1a5d305366a07c9;
assign I97f2b15ce0a74e68d5a4438111adcb0a             = I62f85c1602819e586d9656ba42d263c3;
assign I0a075b833950927c58d8f55264947f00 = Ia9f1e580e8f441394d719d52a7bad688;
assign Ia0886ce792e062e22d0c224158cdfb7d             = I79585885950084095d2ce4a31aa73e4c;
assign I3b699342f0100a2d56c7013da055fdd6 = I0b573d3a86a3111451da661e46384876;
assign I1e805c70d50c2765b4a03ad2982dc421             = Ic3af09106eada35f1d786ed60e314ea5;
assign Ic223e47525ca27261b7db8c1afddadc9 = Icb0841ecf142687c3aa23e68f01c927c;
assign Id9b9a8fe43992ec0793845715dd2226c             = I81e374d671edb31d060875cdfdcd61c7;
assign Ibb5c74ed3a37c5e244e537e8b8d403fb = Ibfcfd3151af0d82bfce293ada44059b3;
assign Ia6a7f9beaceb08d81012f0e72171252f             = I1e22ea5ecaf87499b7106246a824a547;
assign I5915ba867f798193c35a4af58e8cabf6 = I220e32641265b46527ca61111f7ebf1b;
assign I0a9a09b0ab43d2a0f1d1d01e13f0333c             = I0e46eb0f32c91384b07c7b1ba84caf98;
assign I73ce6acb5ca8a57906440578f4ae15aa = I0ff479e61d1a0cede88ebffb073c60be;
assign Iba58175a7fd5c5da650222193caff0b3             = I562b5f77aedd91f0cb3df00387c7956a;
assign I9cea4e30593a1275f4450adb25b5c5cb = I8e87530a131b5a73cad6df68b9e4967f;
assign I5dd29fd1a73df5662d2b636e7285bad9             = Id819e47f502c18dca8d1e804d346c1ea;
assign I3dacee8649adfc1a8b2092f5af3cada6 = Iee17ece482d04964d3c21a092ec955a4;
assign I7c19a79f441ecbb73685db5a505e7479             = Ie0586f4b015fd32777d24c2d9856b27f;
assign I00537a49036c970d6df97b3917de104e = Icd6f8f5df6b4ca4c81855e974db76526;
assign I7401a0501ba69c5559fbf00c77e58dc5             = Ic28248b41552d2537d0478c23e33e0f3;
assign If6ce1f97c23f1d1bf23c283ce37682ce = I2bdf4736022e5da7294a0e851006a124;
assign I89537301987d6da0dbe6cff3caab3ff4             = I3463cbe0d16b14aa670fda6a0d34e255;
assign Ieae92b67815d507df906e1be71d6346b = I1c7e41b9cb1bdb6f649c88c0ed3f4100;
assign I9aaa036a6158d11c235bdc8406d79f4c             = I0aac7a09d9253385d34e87bfbb216a79;
assign I1af89e1ec1210d4d3dafc0927b62afe5 = I7ce064a756dad56d37684d5d7d168047;
assign Idd9f7ea657ea9cdcb45a7e4b573b9d50             = I305967a657db8531d1ae309fa3e3b98f;
assign Ic264e7826b90e379048b094875eeb921 = Ic62fc602da3d16fe13d03a49a21269d0;
assign I89013d61c1ea8da8b1c6071cc21c316f             = I0524108ee49eec5fa7861bed35e4ea3c;
assign Iea6d4bb1137e579b1605a16c578cbd7d = I5364deb983adc2ae505ed2b8c57f876d;
assign I1f00849ea055a7893df386aed162a7b6             = Iced1e0b874918a1c66e28752e340a51b;
assign I706d85c9d83bcfc5a2204a67e5c1f84e = Ied2ea62cfb21602645babc36e27b8218;
assign I53f275395dd6be17961a5edc3e8da7f2             = I670e910f74fafccaa9f1a8279fd6ebb6;
assign I6e832b004d0dddf4c3edb682669acf7a = I2ff317d57f59747c4524ef4278d51092;
assign I6ac24c46319a787daa5c545de8c6eeea             = I02fe6b32b2405fb94afd5d7abbaf0195;
assign Id0f69c70b38b7483a19e32d5982bb4b5 = I6e92a48aaab94074a555efa9bd1e7243;
assign If4d5b48882e9e628cf51ad2ac2f38c22             = I5f5304e4b132f816c87248d3ca954164;
assign I9cb245dceba82553db23cb15854f59f1 = I79b85da6e5ce0b02ebd1619115c98e24;
assign Icab010d78cd66b02e089c74f04bf4e75             = I0ecebe47e1a9ede33c3995945a6ee760;
assign I978d0157f7403d2f35fa648271f4fbd9 = Ie68b31360c12a83c6095254b6f14603c;
assign I84c88b631bed5311cb6e99e58941149e             = If425109071b5310e097d2174625b6383;
assign I70e5f31e8c4f1aa9a9aa21c28ba20d08 = I00d3f14b20e1ea7d726533386e0eba27;
assign I5c942076b173cf527e1be2ddb8560e84             = Ic0f324c7ba05a7cfae9d70b62e30f94b;
assign I3cf2040a93a0184f619ce941c4f910d0 = I579c7926e7b78f4ffc606adc10522f53;
assign Ibed2a63af723a7abf96dacf1951e5266             = I35631cbe926290974c90ddeb9b07f231;
assign I3278841178f87a4d0ccdf8316c3fb689 = I837183265ee22d080e81fea468ab0887;
assign I242a30bdc8699d8ff550b25dd53d6c59             = Iceae425f37f3b1194a2ef5cd46d1b6eb;
assign I73d0e5f3635c5a2c3f1824c578c07658 = I8e1ddd7e4185c28caa71d30bc28138f3;
assign I376a48b7e0195a5aacc76a0ad8bd14b2             = I4faa2187d970078870078c3eff180b4a;
assign Id1b7ef639fcb74c8fa47fd7ef0cbe96c = I9539fcc40d26b13015a864718b116d5b;
assign I21b062856ced09cb9131c01b5e166f32             = Iec2860f518edf688a9b1b2736ae00835;
assign I1c83edeea3cd4c32bae64594a2f8b256 = I02849282dd1bd663fd39baccf41762f9;
assign I6b3cd79aa87235ff174c0299b855dd3d             = I20e7b48527e4456874d59e50c723c6a5;
assign I0b930276a1887380da03c22aa8fb9adb = I5d6e576b0fa7e3219aaf9ccc345085b8;
assign I814b62120953991f9da055f118967e05             = Idd60af0dbb02680e11c1b1734f23b895;
assign I63ec886123f0ff76bfa46c2d6b2c5760 = Ic0191941cb968bbd7644c21767423d2e;
assign I3f33901c407a87e10d86c13c83dd52eb             = I79cfbb5d5e920bc8cece60565ee0c5c2;
assign I32bf44d4f4df42cb664e75ccef06fb34 = Iab0bff1633e2f3ea0bfbc291f3ab5d29;
assign I241622b0367dde514f96ece55c8c3964             = Id765a3f659dcdf01cfe23cafdf066f92;
assign Iadc0319541fc978cd0efbdf5b3af7078 = I8850ab26807dcd55fefadf6310729ca7;
assign If9efe7a1c359ec03014a52870ac13aec             = If370aaa56b4ba3eee873c99a86577c3d;
assign I9f4036502b40315cfa7d8bb9b83b5806 = Ice59d2af73d0b0f2ae91a2ef0c2b7f04;
assign Ibc73d07e0c97a6fcae791e04106cb082             = I4508376202467dc1bebc69757bd5f95a;
assign I91dd649eab4a8eb0f8d97553560d3b7e = Ic4efba3932e598784f5b9ad6ad04772d;
assign I2f3ab9654e515a54e22e73d6c130ccc3             = Ibf115f80ad72df8599073c05ac58e028;
assign Iee09e9c54961c380ff7e1758c84d663e = I9ad2f6fd2d7f68011fc926ec9abd5c34;
assign Idf6875955525d80dc660ce956f4a84e7             = I27960a9d3923d053d466955c660a91ca;
assign Iaec27722c40c7cb0c0baaee4d30adc72 = I5f0751fceaa008feba5c6867ced453dc;
assign If94a1abfb972f63629d07e64dc23863c             = I7c52711e3b71823dd47861341d22adc3;
assign I5fe79d8695d426ba54609af4b38bf2dd = Ifdabf743a8cb46b7053000ff48ea0c60;
assign I0c0060fe260afa3cdc72f35ffb6938ff             = I547ea6a130740e4b0bb85f6c9d3a6549;
assign I8a2b1e09c6f852b0aa4e599e7ef42187 = Ie562ebb336e476a81f20a652d4cb20f1;
assign I6627bcdbaa8afb115123777abd45435b             = I0ec19c18ef7da4793427a00a652a9a35;
assign Ie1f415cbb2d3e1d46f2e0e4201fe7ba0 = Iefdb8bd28839af9413a3906cbfe715e6;
assign I70d32affde22f9dcb2d77430fca39069             = I640d147f241267ccc89f9ab132d724f8;
assign I46a75678565a43e0da6b6dc55686c4c8 = Ib9d58222da98f29fa302b4896594fe26;
assign I76060709de3ea188748849f043c59ac0             = I3507152877484394769c12879ce0aed0;
assign I200bec7d713bc7f05dc3931f20523763 = I9f6751c15237c20b0cf2175575195ea7;
assign I07b9b1f4fa01b16cc69356057d3b6154             = I382f86490f568ead2dcf51e8bc6989f8;
assign I978b7018cd38c7c4f0b6199cc46d258c = I081e2595b18f306a74d070203447ecf6;
assign Iabf572c97b48c6a7dcc19e56676e3a82             = I953178c54a672474dda2f48c70ec21a7;
assign I9d298dcd244445c8a047a1ac056fb6a6 = I3b84dad6d0dd8730312b3e20c6d5a2a8;
assign I5814a85c45fd0f7be21ed325235fe4b7             = I13b43982093e885ae7bb04a2b61e4eaa;
assign Ib5de0226d215418202f2cff36b573daa = I6ea50be10bc990a1206cdc9e28e0c4c2;
assign I2288a6ad3b748b716249f4adc42d52c4             = I3d7491ac28a4adafbc138d17f08c9111;
assign I58e42ededb36d8aaf022e7b42a8fb36c = Ifc1da524e7670772834d521a6fc4c96f;
assign I60cbd4369e7ba9b6532f279e5c59084c             = I3e0ca15752add87cc01981e7d89d53f2;
assign I8017904689642a7e3d82c34839403614 = Ie2d946edaddd3c87f328e861f3e72c0a;
assign I95361d5f524ccb9feb42811af5c482e2             = Id1b152deea3ee894ed5a4c6ff10a6fda;
assign I773d6a848aa20abe6d1ebf8f7d6dad85 = I43c2fab87f70ea883321ab82de85f133;
assign I022df337bcc05ac5648b8ae2e42f3a76             = I7df9cc0e3ad69985fe9a3c8f2dec1de3;
assign I8bafb2d0a6bf186c179ee07ed51a2e33 = I24645082ef16129eed1c574f5fc601ca;
assign I2ead0e9941e2280309ab53535b1e1ac1             = I52910c0c2d26095c965d32b85e850d92;
assign I63d8a99e826b0d6a5051fb454f15f44a = Idb1efe99b5d7fd567a7f82cfd52f7eb8;
assign I3e5139f24e3d082eb31b0e61ea9fa1aa             = I93fd4b4f7d01ec59834f3054fc2eddfd;
assign I0b831c8e1d7187024eb93f980cb04f61 = I1af02ed6cf00d4cb0704b5e44c83bfa3;
assign I60d9a7f95fb8623753002ecaf9a4efcc             = I481b6feb1f1ced501a157b06a4782e05;
assign I17867f12563819dd7b89f9079fb0a385 = Ie8c0fac00a9de74870e59cbf9e87a39b;
assign I93b69bfb228db4b569a6772179d603be             = Ie99b8f3190ee307e743255156b7f7f90;
assign I2a2b4eaef143deb9e61110334dc5c2ea = Ie4827dc0983c1a63053c08de6e36d375;
assign I85c4d3d6c8408c6f38741257ed177ca6             = Iac858597facbc0025a4760eac49531fe;
assign Ieb02d465c1ac76962dd663067ebcd445 = Ib71611afdd0381cc1884f5ddbbae1acc;
assign I23a74ea5e7174d95e6d16a5e85ac236b             = I18c2833554a5b358578e7b6901c91c0c;
assign I6ad4bc4bc7c0f005307199814893faee = Idf8d15c7bd7705b9aafbda09c3a5b46c;
assign Ide530e6f4622c8a7b101b6dce9650e42             = I0cc6945a47b3ffadd1e52e3f71c9728d;
assign If9a814db74759469b79411ed7038c860 = I7f720a18542528f0c9bfb14f699ff4da;
assign Ic95191bccb18e26c10e56be395ca6b1a             = If2807866c5d481cd31c69b67ec537a4f;
assign I3d0f05a6136e0c14536830bc53a5333d = I70a4926e9e6a05fa9ee51a26988862fe;
assign Id0f75e19b94541ed5c5c352d13390d2d             = Ib24d495a86e15d9c8b2c8d360445e511;
assign I1f168715063587b7dfb01e0fefbca615 = I38fc49afce0298846ae8ed63ae715e81;
assign Ie697d28d757df82b3901564bda43251c             = Iad2cdac80bc26a0c50335c6467921c94;
assign Ida3cc6922fe4edded7f2e59b909d6d72 = Ic6fd9592d2ffcb8f4ca83c6f0bd19975;
assign Iaf0bbbe791bb71d0f557dc71caa5fb87             = I18c93f107d0520171864b789ae9707b9;
assign Ic2b81c5409d555402164dd12ae7decc4 = Ie4cda4648f6ceb76b8fb74f290ab6439;
assign Ie4ae993ddb776bdffec843db0def2f5c             = Ifd40aae90a89d2420e43fe4ee533a1a2;
assign I8edabaa27753c6f70325108c9c1b12b6 = I5707d30ca29842b6a96cfaeb44ac6668;
assign I4dca2dd40a7127ce44f83b430a34c738             = If46a176f32240b03ae959e9ad889fc2c;
assign Ie58289ff961fc431fbf10f78fda337ab = Iddc3e44d83e8253e5129b6cbf5082df7;
assign I8572aedc94f7243ce5eacb332c81eae2             = I5e7b386298be05835cd24554966cdedc;
assign I3ee219716889ea93423603105de22c6c = I94009bb7239be96243902ab0f0abea7e;
assign I4102100fa5f1dd299af0190862efcc42             = I5258d2bd4ae07dcfe7e022b046800856;
assign I957518cfe822b5afcc1f7153e07e26c4 = Ic308610ea8bb62ecb6094192e02dbdba;
assign I224bbdf94ac86c5c376d1db4f4d4e060             = I14da6601ba08fd3e9a2bcdd20bb43536;
assign Id8fb66bc4afa4f7f7f4ca0d7ce3f5543 = I85654bd3a07b4329aba17d8b27777f4e;
assign I6d83efa9f988328f487e9232bf2633a2             = I76bbfed1a115c2f503531682cd171185;
assign I3beb0bdc4242c12a068f7aec11bf022a = I975a87bdda30c5b6be8d2f0e4b107450;
assign I6734123aaf6320da75638b212812732f             = I64f37f25618c6bf5b35e863e3be05a3e;
assign I629a5a30684270d00605b4fc02eab693 = I8bd2a9d90074500698b302cb8db7f03a;
assign I52403a0454e5fa002e79eaab7ea497bd             = Iba3b847497a7572624a3a1f172b47d3e;
assign I32aa431be1c47b8c52c3b3f6d371f439 = Ib5ee5a6ffc45ed1fece0822dc4619b57;
assign I96fe3eb633eff6958ac575b997460bb9             = Ic9885fd472d244d4810bc9ff0971dc65;
assign I88d8124a68d50e1730a87914ed6b2a55 = I235c3a9fd3e8ea1cee762c10bc8e2c53;
assign I69f563e7b7ad483893ac9c4684349769             = I5753bb74c9d925b91c0173bcc320af36;
assign I474bd0d0a044aae82cfb1afbd3d40f74 = I582bd96afa764ded148202f738b7a1df;
assign I7f6dc6f0f403c58f9aaaa70c2383a666             = I66cf73ce0a93f90287df52adb628716d;
assign I2bcfe7aeef8f2b772605c9ad10a289ea = I5490039998187a1a2efc3549e3dee7d6;
assign I4f1221ce7880729fe584b42ef3afe6b2             = I84a477263ea86f2014d28e9ec928fa1b;
assign Id4a7c3a22060cfcaff64e2a3980dea91 = I0615acb0f7cf79b5f6ae8e91cb525dc9;
assign Ic08e85346f61da036a15345a13ac12f0             = Idda9e2f9a5e24406700b04e6035dafc7;
assign I6085d7398ccd685c1a60a21e4a15a606 = I7ec15b73b2811b44e1e50c74a9f921e9;
assign I9160d11439c5140c0109b5190eb82e6b             = I694ec5f3a1e7cfc02c1af8369064967c;
assign I203cd1948326fb3fa3dc14423bf3f992 = I6fb88d97bc9ed37a06b729020a1df140;
assign I66391978843c39b6acbdb4847a01050a             = Id0c6285ee3789c104e483a5626b5827d;
assign I67412169057453e2fb39c3b0760039c0 = Ic5cb81c821716a8aabf8cc2283ff73ba;
assign I6a6eb62960b616043415406ebfc21346             = If9bc7b1498733ed921b51cb613c2cf53;
assign I520d93aaf6b72a2ec7c23ae4e253aa07 = Iffa06a336949f56f4e5a88a06d8b7e60;
assign Id667c80003b5541de9f84d3b8709c828             = Ieeda4b6b301d662ab9be9f6b979bb1f1;
assign I34a77904a4a75d2907acd173bf27800c = Ic68f500938d80460ffdb33a0adc48298;
assign Ia030c08757123aae947f86ab8bfb6d94             = Icad98c93196218a7dbd25af042b4a32d;
assign I7a4ea8ffce8d52bb241553a681408dec = I1500943c4a550e78fc169437b0a663b7;
assign I4f756e4125c8af5c412944b273e01cb0             = I408e198b0eeade8b94c27ab7e04a8776;
assign I8e89fb1ed1d604bbf0177e0c61da6e94 = I22f5bb821a2571d1764978fd76c8f1d0;
assign Iaec1f186cb4a65da21d41e637fc628f7             = I24b90526a93dc177a5d23b61d20f8797;
assign I5d2148b5809cd169c41663caa441c464 = Id962beade26396738ba0e97f67d5e261;
assign I123a212546a8ac394051425db4924812             = I4da324410e88d8c9738949c287e7bff9;
assign I5bb0ab59e3468a9a95b65bfe58acd6a5 = I7c965c047d862c973d09a81abe03a845;
assign I730634ea15ac94d241f3ad2d6393a227             = Ie24b89ee61bddac2f2bbf1b8b5dd437f;
assign I3e9c216d05b6a9c1040616a42af371ff = I0b83f4ef8ba9badb27e81b32765ec5b6;
assign Id2c9f7ac95de07148c54803f69347f56             = I27b99df87eefd6fcd484ec321bb73dc7;
assign I4902647240aca7d98844546130944322 = I42ae0c42360c977b35429ce290516a6f;
assign I45c5e6710240685bf54b73b0d7a64271             = Iaac7f8ca30f4e74e1ae5016a222673d7;
assign Ia4c22694be7c5db34c1b875db1e91ff3 = Ia03836a4e93d2f36513227d1dfaea0fa;
assign Iebdc41368d57498a04fa73e30b10a966             = Id3076c8e12f28723096148d8cf91a13d;
assign I0760280d5f5f23d9e06752908f0bbd96 = I6d423a7d17e05a3c597ec6ef6c5a7cba;
assign I47b878f27c30f79a37e97e022307e9e9             = Ib2e36c2d0a51f5b953b9f368f11bb295;
assign Ic807e0ddc985cffca6a389b468aeae49 = I2c420acf428e44cdd9ca9998e276f258;
assign I5061e13a179d27e1ba5f89ce8ee0fd4a             = I9ef5138c78fee50aeb2568def8bc62a0;
assign I9e3643f805ebd6623b9ab7ab41c41ec2 = I14bf11ad80890227e47fda26ae1b9c24;
assign Ic7ff9cde71054c1ee9eef81eabdd7061             = Ic1cac944a0ed80e5b6e3821e8451045d;
assign I0dcf2ac5c06f517ea62c1ccd5acd9298 = Idd474d80b50992537d6f527faf279800;
assign Ia0a02781c674fe5d769206448d475245             = I915f18e8333d52f6ec4162fe35317d17;
assign I26879becf6ee094c9b8b4969c9377af7 = I2eed3d32a27d51036e17c4a21382b4c1;
assign Id66c47fd69c175a4393e975a269cf053             = Idbcf9e41a431a42028cc99d6be0c46da;
assign I3daa291236c162f58fdb9587a880dddb = Ic7b6dae3017b55dd3cd27423d5f1b0ec;
assign I0f7c32fc1548fb49b8041f55c157498a             = Ic46dd35355bcd4470886fbd416b3c75c;
assign I2e150157b54bedd2bc6d31435e29af0e = Iae7b72abf4d3c536330a229e3836b441;
assign I4939f69abb1eac56d5021e06406a93b5             = I0765c8beae32257c6c37dabd94cbab7c;
assign If392bba16edcc39c846dc23bdf59f976 = Idc5e98f6958786ccf95d39b922b42ea9;
assign Ife1190f76c2e251704c2960c23330a48             = Ibc002286423e5ddf50b8ea25ea1b3377;
assign Id0838a2f54127e6e86536294821b8fd2 = I2a4bbedf880a9a7b4e1bf946f9f96c0e;
assign Ib06b60cf9933dd8952206c5f3ccced8e             = I714b85ebaccb1e11d16d53cf6bcf65b9;
assign I3d11d3dc5ad053fd7a82b00d4ab4b180 = I4a91a7c9b2a0f3552b8f2ef4e2398be2;
assign I89ffab735ee30423c82e079ed98216c5             = I864ca16e4e93b435a94fb012d995c7e5;
assign I1f67b8b8a325071662e006b730b1cc8a = I3b8cdfb1440732ce98cd1676e05a2af1;
assign I634f0ce28934600a1a31ab0d8e59b4a9             = I227ef7de18494a9f62b2e8cf37687840;
assign Icd7c05e9200f346555aa6b82827ad164 = I3fbd40faa4c3b78b547b8348c466fd1f;
assign I1a24e98165afa62bd14986911a36fb6e             = I535a78cff546aed9fbd1d79827d56fe6;
assign Id136b4b678027d89c31614cd5baa6282 = Id6b508145cd21ba088ab8fda34577c35;
assign I9c4b34b5fb1d59c132bcaeb6258675df             = I90cf52bd1332ea1b955e8c193b670218;
assign I08dad437a9b452f65231279ae25ab7e1 = I99ff29c7ba68b5d0819f1e1bead51287;
assign I9494921d8487ee0b314f75cf0380fd2f             = If7dc2cec6ded3b32d42281d08e871513;
assign Ief01dd5ab84a9f9b05e48b07e0d1ed54 = I2aea17846a53e2eb2968581ee2c48226;
assign Ibaf00a6780325882067a79f0c4d693d2             = Iee43875ccb00a79e67acbd3e12cb516d;
assign Iba8886370777ea357fd7c1e13bf03cd2 = Ibf2a253afde05c905d0b2404c5a808a0;
assign Ic23e01562c8a753fd70c343297be288a             = I7aaad9fdd239670e028a896695c01216;
assign I9e1e97a64e15a82443cc946178c11d52 = I24f82a3f2c0e8df486fe495dd95cf8bc;
assign I61cc8a0f49e393721a62a776e4793deb             = I4a992ed2550a3c5b346158ffe18c255d;
assign Ib830e17254cac0158be2b443e3dd4d43 = If06b00be0356a2be5074d958ddcdb2f9;
assign If2b3e7d1541cbd8ffc2b4cfc3ad13a57             = Ib2eb28843cf201e8c6f8900b7029d42d;
assign I819741033c6737000bcf4a07a78e0938 = Iae5d6faac1f5685cb1d400ee2b1d85e0;
assign I71afab29cdb962e1f1ca21b61dfb50c6             = Ic9a5b2c8aee24c3fbc7e92b8fdaed5dc;
assign Ief41b57c092906a598c1cdcfea9b1062 = Ia98a6f01e4eb5bc74d50d350e79be426;
assign Ia284f974dd8a526f31eb81ed71a06e94             = I6996efa8115f38da03518dcb7dd42a4d;
assign Ibea5db121c78f1b6d5288231ef59d04b = Iabb01dc9980b4879a7356712b51df0d6;
assign I3e3ce8b4ead150a6eae2e5c701c7b598             = I1c4bf7954b4bd5f4e9c176a3ae1fc28a;
assign If9d3ee7956572ceb26e7d60077de7e00 = I604283449f13c7b225ea03f99f2e296a;
assign Idf3d79da44f2d686f5bd43c3c1427430             = I55d0fd8eda9c128cacdebab55a8dda5b;
assign I46fa901f3606f4d2ef11e13cdf029826 = I68b152a599887c0039dd9d45c528c219;
assign Iefd370d0df1a93639af482f78a1e8706             = I02fcd92b426929f24b9a8c063a56c0ed;
assign I9918607fc0fdd746a6830800696a9439 = I24135210c23b2422a42c90ee25594191;
assign I3ed2da9b53daac0852a06ad1acfad21b             = I3202a0ce45afe072eb955cd6e0789cd6;
assign Iac50ab3381392442d8e7f18bd9ecacd8 = If4308ed204e33952c9931f8fe257aca4;
assign I453fdf4fbb5af5bd28a20d7643da9eb2             = I06c82466a2ca646abb62bcaad3d63748;
assign Ie8bd9deffa3345851a9ff645b5bd1ddf = I2b600e5f5c146ee97c4044c08e1f5ad5;
assign If8125ad3c9e7f0a2b84106064d320996             = I23af695cf96a03638f0c1ef719d8d530;
assign Ia7d6b9edd50a4046aab863855f9491ee = I852d5295a32984af00c95f6d9389555e;
assign Ifb6c65a00d9a2c31d8b1119b949828d8             = Ie20b7fc4110631c1da7de4c7f38e2581;
assign If8c22f4e0850faaa35f617a99c827f84 = I33ee415d85e2bcd8f975d34b880f6ea7;
assign I43f2b69c6b427de3095c44d4166b77cd             = Ic6983ef65e0de21992fa0b90ddbdce9d;
assign Iee22d62b28aee7dfc6c9304c92214e55 = Ifb89e7ad8ef661959d82b7c22f187243;
assign Ie9cce5746a83479a567bbaeac6dbf497             = Ie7c2317cef621a89ad24c8b5bc79a39c;
assign Idd235ad7cda4d67de5992f50db3b8de3 = I9fe16403fc21bb1159a5e0305fd1ef69;
assign Ic9018b88fa91fb638bbab0613795ae13             = Ic58955d8604cb1a6a20a199372d44774;
assign I6bb6fc0f5773f1386ac5af0688f224db = I207a0f6184a0b3be71766a8b47ea5535;
assign I56873feb8418005b5661c7382f2dbeec             = I8198473d2a666821cdf398dcf1b0fdc1;
assign If44d50ac2bf54fad8236b3fcd9484792 = I86ba73ee348f80e2f9891d2ebc8a02ed;
assign Iefdcb71f2903b11f5cb0b8857f7a1727             = Ic60bdcbc8a55bc760e52c37aa3030001;
assign I9039a46d1a19d43e6c1cb3f0c162efb1 = Ib6ae81df8db1dae269437861ee11ec0d;
assign Ic57eb4a034247a4c952d8224ea9f2bac             = I987cca9a9fcbe4b617a7e524476431be;
assign Ib3c48b1a31a7198cc8d4fdd10d0c2db8 = Iabdb9374e5caee281c25b003624b2c4e;
assign Iad4ea0196eb32f9a152c9e6fe5059e46             = I765c7209f3c7173362057fdb60aab732;
assign If37efa97b30f1c80267e986fc90f759b = Ie5d9cc18b2dd300132470f206452ff17;
assign Iadbd245bf842aebb456417579a3e6296             = I2c117c8ea4060a5094453cc6140c9bb6;
assign I42e35cda79f11acac889996660ec32ab = I1b695aa715615662eff7065c742b0859;
assign I9c15a6a5c0db11ede80ff6d04c9a56d8             = I56a6be4115d52bd49fc003b164fbcdb0;
assign I0ac3076614fbc543f41c76c6be389a37 = Id0ab747d92288f23cef793567b2363d1;
assign Ie95f1a7e0effcec0aa423dc803056a13             = Ib834a7e4f3a491e351e2e49d809d2448;
assign Iefae454b50cfb5b83c8016d5826e7670 = Ibd12036702fe60b57354b3aac921559d;
assign Ia8ff29ed728e7f2ae4213f00328b495d             = Ifdcb28209b39b8d99c2eb00a72921a75;
assign I86cd5db563b397776c52a89f0b44e442 = I671de3d408b5b783541663c7f1e3a6fa;
assign I7103aa739616a39c03e675ea0efb0335             = Id721a94e50637fa39c5bf6124ecfae6f;
assign Ibbf7f6c104c9f3163fc8d6b8a33ff5fe = Ibe01835305315fab50269c72ef849b61;
assign I5827bc87b5db1801b7db16e1e61515db             = I72ee7b62c165dc693cc6b5185970f7f5;
assign Ife8ac54e4431329086b20d2111eb4f28 = I138fb0c48f2d27e3315e237d9e61d653;
assign I5b4305bef5b4350c1d7ae143667afddd             = I564ae36637e0cd6a8a06289e95823572;
assign I38c2a0e463853ac84b1f4e5c92f44243 = Ib1639811de6eb1c38257800c201fb704;
assign I70717726200ec02929f679ef05496455             = I085e99650c86078bf02f1b2aed141add;
assign Ib73515d47a61e4a795005e8ae6bb2968 = I169d8f2bb5fde5b202b4239b7a7f1ed5;
assign I16e3559c63ebfed83d6698fc9a9cd93a             = Ie4e63cba44dee9885eeae32cc844c3f5;
assign I48b52a0f686c64c91c6ef4b1ca47593f = I2b97a79c90f6578c8b2f321f8d598cc8;
assign Ie7f3f1d6cee7f02ae1b17740ed54c049             = Ic054b062712da78ddd4a148bafeb1a0d;
assign I9ed8d0fadbdab4e176b2d03549e41c91 = Ieed4c810a5bb69de112522dcf00b16ed;
assign If5dfdadb3868ed5a495007362f7db648             = I81b01fc018ad1c79ec03a123763e95d9;
assign Ibed24a9317d456b1a27bf71649c9a751 = If926d98f659e8fe4bbf36ad2c5c852c5;
assign Iaf1e4c7dae6ad89567836877c08f57d2             = I1d38ff144c3dcfe4c04778e50a044d5e;
assign If6b0b5b913b2f16e0354a62459f87487 = I8ca17b6cf35e1b1f8f601604575d3f27;
assign I88c10c47ae424fbdcb852fbf1e94127c             = I2e31a90886f87907d19d0c034caeee9c;
assign I6cf5556c5887ad4d2f85b26aefe2aabf = I9a6923c6368526a53ef70e16471386ef;
assign I06c7728ef64be8311f48d10d766d0c44             = I7c48130cd79566b1f1e30b7c709ee5cb;
assign I4fa8769d910cc70e158a0b649ce1e1d4 = Iaf82668eb49248709540f2f529f1b3e4;
assign I02cbb4255db2b21ea32140f9e9ddb36b             = I3868c6ed60d1f0ef9d3ad98e91931acf;
assign If25316f70adbd92abb74b4338c63d7d0 = I211f8d7f97ebb8eb3e50313513abfb1b;
assign Icd09aa81e9b43528af73e23b2f0f80cb             = I7fa57873a108e5894f837bdf45979b8d;
assign I38b3f467871a1646a7694cc6433b5c8b = I0fd2f706e374a4eb57ee26ab50201e15;
assign I6ff7b86cd7f63f9243646f1be10b2577             = I59d4025a86d065a84741dafb86b50cbd;
assign I0c7ee025ebd05956c96fd50885d627c6 = I83ecf12f3b38fc14c3b75e47b71ecc09;
assign Ie631e40caade823a196370fc3358f042             = Ib28a3fb3dcdea36c883c88b017fefa56;
assign I680660d6ba504eb445d2588ecfa046bf = I304ac9f96945546cdf1b6f1fa7136731;
assign I6ebb2b94f0f80425f8401ae823d92a1d             = I91e4dca55e1a5d1d8ddee5c3bd1048bc;
assign Ia861785bea48073ffcabfd97a16890de = If5ae6fbf843fdeee17945bc5ce81aec8;
assign I8c35c5b343b552c22000e194c517ca12             = I55dd62b8ff91323075533e896207c1e5;
assign I8619e41804844cd4d98818cb8387c3a7 = Ie039ab562e9cf90289047b5425186123;
assign I37dca40506d61bdeab1255ed4892ca20             = Ia30ca84355bb976cd045e969b2862856;
assign If916ac75b729dfffab3cf6b0029197ce = I7a9800418bd5c195fc47a72370680b56;
assign I4a2c3204a6a9936d4a215b46c0ffd045             = Ifa1359651fd7e160301261bdbb81b02c;
assign Id4f85daa963c656cff69ca2a821247fa = I9b8023f4dced915cd52c91bc9d4ed78f;
assign Iee367c535d9c39f872d2ec043e7e7b33             = I0b465f693268f6f56f52d41165bf66ef;
assign Ic39575e662d7843dcd7418a7e8cc4a75 = I49d35ec6369de10afb15be8e0cf135c3;
assign I67347c413b5efd8ff9e0d5bc7ab2a047             = I3deffa3a53b31688f28dfbfa66571d0c;
assign I7c445b4e53ebe960faa00a46e00d66b4 = I5f6a61c9f0c67510e148e596f553a4d6;
assign Ib02c0694762c4815448b2c8d3df767c2             = Id40c9857a5bb6c8cdc616fe68d8dc39d;
assign Iede71af4d6ced16d85e2576f035cc712 = I48e3309c61918c3991852b45d9c72ea5;
assign Ie76b0739aec66f8860870e66e87a6445             = I26754124b13858a3b925cddca5cd8c5b;
assign Ifffbd3dc45d11e43be5de5a276300bd4 = Ifa6e3541f5e12bf9677ffc51d0392749;
assign I613d4b1e3b9e812b785c9cf14fefdfe6             = I2ebc1a7d32a5457de4d35b6bb25507d1;
assign Ib7be21d644d545e6671098d3d8622fe0 = I8e313ceb21359bcc44114ab217b1c394;
assign I98cee6efbbe565d3a4de16703189782f             = I77bf5b03fa300d1dbf8df5ca4acbed14;
assign I1bcc55c2c22b349f421eac34341487c4 = I3c0a621dbef864fd1f566bc2e47f32c6;
assign I4a777f0dd62b19dd340ad31517c4e789             = I6c1c1e404f92fc80495e8e5d187934a6;
assign I5117b588204bc017b2a94a6e1097df82 = Ie61f299252b8fecfd3e8634b64df5a90;
assign I1e50c90010a3df1a8ce1cff811cc7a0c             = I126a2b15cdc34d88d17ebacb3681625f;
assign I7c6e35ef749c858168d55bcabea9078b = I33ddee677715877c11a1df45cbfb01ac;
assign Ia642db613c0ec1ca4e69afde7a14a839             = I9c5ec8e21febe3ebe00c53ac8b21d1f1;
assign I84a9bd349a6cd85859437ad4f9e70693 = I4c9518755c33d725221ad79ee6badba9;
assign Ibf981c01a9d44cbea3c6d8ead92bc2ab             = If27eaa7cc4d1b5d2b7a962b48f0919df;
assign I27b66137a39cb30b8059289cf98f8a19 = I5cac08dabbb6de3b01c821d4db93a8e3;
assign Ib6ea4a822da2ea32e0abf6cf8a33d295             = Ic15f443512d68537f9764a3ba88334f6;
assign I89b31cd7510ff82f89398b8682f040f7 = I1e96d5af3d0e3fdce39530dfd0131a7d;
assign I2eb90278aaa54b9c8212b3b4af7c3617             = I47b266262fb5a98f66706f460f1248e6;
assign I801f6e47b9e4f6b6acfaf6f8369ea217 = I373841aa2bcbad8232d54ac9035a3ef9;
assign I45bc13ae0e0554a79c62cd9c6aa8f2a5             = Id301f31702270a4f8e9964e3a75e3d62;
assign I6f7db7eb1e5bc6d08ea9059ef7c31949 = I3c3cffec9f47c9979cb9503f222f370c;
assign I864c33e8ea204d20a9baef4584f22d4e             = I097ba3ae5a0232ae6aa35478635640b3;
assign Idd01178431a1c4a53be45095dc897c33 = Ib62b02ddf0f57bee49838d19783ef6c3;
assign I9905e2686b350e8a6e7f790563a91294             = I3b65eb49005aee57f61279c5a172d158;
assign I64ae03b30dd467619e71498ce8126df4 = I182b43872d50de6f7afb700f178b160e;
assign Icc93450a007cee4c0a42717ed7600528             = I8573059885be4373531275502affd59d;
assign I36eba1bdcf4eac1c5c4b458515ed3f6e = Iddcfab4a7022e0f12fd20cb34e9b9d02;
assign Ic4a6c02880a9aead7353332708e3f388             = I627f9d9ac0c07ded7306fd14773fbee4;
assign Ibb1a5ae8240913132795df9605e82ce8 = I68d6769541fdc3df321e192f645c667f;
assign I6ad3228e0e2e1f19648d73e83ba5a229             = Ib559f45098803b21622fa96ade885abc;
assign I597865149cd8d3e173f8aed514cec357 = Id051f1d5454802e0eb37e22248efe8ca;
assign I995d2809ffaf0ecda6a004d01cb9c8c4             = I10e294379879538ecbf65fd423e7355d;
assign I667f0a049c87ac48820b60b2346de1c4 = Ib08897f9216599042f7b97b137e07fe1;
assign Idefa29d4d4e2a6e9147f84893520096f             = Ice861034cd3b2f3847f325dbc9f52d08;
assign Ieb1c4ec26a969a2c1cb60e0d1c67b5cf = Id1dce2b9eafc35fa71df33ada4aac539;
assign Ic044d7419cc43736d278c2df33b4a3cc             = If201eea7e0023bb17fe41dbb4b5ec076;
assign Id3293a3ac3bb53134fade82ddb8aace1 = Ided55428cbb77f454c2607ac783d7548;
assign Ie099210a99a4899c53baf39559592690             = Ib15f9bf401d734008d6a2b9a00c572d1;
assign If7ed4187de370efdc1b9798bb6b05232 = I275cd09649a750edb8ae8313e4e1e279;
assign Icd2e75e47cab1d539ba9ff1b6e1d7155             = I581f4e137ec21e639eec32a1675f4750;
assign Iefc40b941a682059aca6ac8abffe1cfb = If533578cacb685a95afbb8e1c05d3c07;
assign Ia1ee5579358b564de06c08ca418a9bf4             = Ib7ff7b93c88fc8d9bcd915f0c678acff;
assign I746ebc4b00c09f116eb087dfed4bf89a = I8879df010bbdf6e5fc9370e2fb3289b4;
assign Id3e0c98bff2636e216b4d3a0ffd51054             = I34dc9dff97e78a2d711f75675944b0d1;
assign I69683a0683ab00462065f6c3069fb6f3 = Ifd3d4f3e2a388b3c70e7704d6351e0ba;
assign Ieeec71d9df4613555fade2ced7b3baf1             = I8bc35065fe56bb75e6595937aaf9ef2a;
assign I183ad57174d779bab96973fc5ba5efd9 = I7c791c854d0bc28e8dd787545f8fbda0;
assign Ifc8ece44a4e68c3117eda9e65f3084d2             = I1822ab8ed690d872380ef820dc4282fe;
assign Ic4e5558ac995583236747a83b3f54f33 = I90b3708abdf742370f06cc513ee307e1;
assign I65354f2069de0c25bbe7cd50fbe892aa             = I1a1965726584c6c91a7e20de63f0fce3;
assign I12899b73e235f01bce4137c479f6b300 = I9a403c511fe2d44472ab319a9477199c;
assign Ife1164cad7cda4aa9a08d94dfe86add6             = I08c5dcac6674c1671b85d07a55a005b0;
assign I8dc3438a0d2b1c000f2b581f9a7ee588 = I17d32f292758416fe02527dfd938fa0d;
assign I4931884e3544af182bcda9061091a42d             = I40d67287bf525ab2696c30755d6babd5;
assign Ia589b25714c687f50bfa26ead5cfae55 = I446857735e680cae93a24dccb59b1924;
assign I0296d01fd3f9a269a617efd4beea9b8b             = I60dc8e5b6204e3a5fa32e79c5cceae94;
assign I7e4263d478638c2f3127394328deea11 = Ie536879e6fa9be65376d7f00e0fc40d0;
assign I106deaff50b8480eac31ddbae2ec7c61             = I0074b447046d75787aa872d8167171aa;
assign I1c432aa61cf7d02567ef990929a15696 = I3ade5535a79ce83857481ac771cd8618;
assign I5669856f88f5e2c98f64df696db76414             = I384965816ec3b915b9b623ad68fcc4c9;
assign I64531ff978fb8892605f2b0dd8422873 = I9ce3942aba354c1fd7d6b9a39c994d7b;
assign Ib3fb10da528d450251764a9b9ede0dba             = Ic0e2656bee7174384f7f952dbb9da619;
assign Ib8c44be17e150cbd0b49d41c060f95f1 = I40a223380fb4414a3f26a08cb90025ec;
assign I9747a02384abb1c2dd1f52b3a5a999cc             = I4cc3b0546ddc14d78da59e4981a77b58;
assign Ic45b89f2b51ee014d9a0fb19a7ed7619 = Id0b1c46fa4caa63a4c63a44ba3c5ef8a;
assign I2795d21d343b83a69146314a2407cfa2             = I7b680caf7d0d94114fae1d96ba374e68;
assign I338e32162153b4ed5d991c44c38aca27 = I88a89b2d938552458dab9bc34728959b;
assign I1b7a401bc11741e6f011fb9895b5c797             = I7f8986a922c03b6afb5786cd2e1d5288;
assign I06c60ff1b8b447112b28f71eb9e3944d = I2c6c6041c9c69c84f4d64af6458955f5;
assign Icdc9e676957b2223d60c413331fa982f             = Ie7814643e3833736c0f54b39f91fe792;
assign Ic2cc5a2da05052c4a68cadde2745b44e = I0c616f736879c28a5222de3d6f49a587;
assign Ib196f5bcf9152703dc32c5101076600a             = Id1f0c95b85ee041818da4fd9b5466c7d;
assign I8073ab2d9dc1d68d0bb4694ff206995f = I44f170d02bae7fe044456e125a98451d;
assign I165653ab165cfafe2b74cd441331f9e1             = Iefa8421c0c908de69fccffbe22f40911;
assign I6aec90f4d15da8590fe767c4facfe19b = Iefbdf686d9452a62cb99cf023a4d9fe7;
assign I340c98b886123c541a1b8d9fc8a6d48c             = I4319bf1bbb31debc7f58157b75025134;
assign I39a8cf4c424841d2b367cb3a1207fe03 = I830a4fffe1244e071eb82c28ddc4a308;
assign I381f6051282c062ccf53866830344cd4             = I4a349021efeeda16b646979a959bff6e;
assign I031f3e2575360f675bed8e87a71755d7 = I620b8ecdcaccc1ec80ebcf9fa6af0017;
assign I9fe11f6c8147391aa4a5afd1a4e4f731             = Iaae0c136077ecc36fc382a76abd550e7;
assign I40feba64660df64a02c3df651a2ca26c = I94460b6ce7b776bcc5eca149eab80c26;
assign Ibf80bb564263ea85bd886a8617f09bb2             = I4a442564148493664046e7b38cc6cfe4;
assign I985f121a0212a4d64ca4a47c1c210b40 = Ic3ba4531855366e9a060cec1c7694844;
assign I72b1bb104bf2843f161448baf7aab44b             = I12cc5eec3de8ceb3ca084194d430d9a5;
assign Id4ce64c9f467d1b1c4bc9099ab855db2 = Ifad8e46fc3844bbfaf434a14f6b5869d;
assign Icfc21935c007fbbceb2a67ebe1a68a0b             = I56db71b7df11c35080cbaee80c389c59;
assign I01c6d49bf9698d7621a545481b129692 = Iec91b3ca3b54010755d57f8b8ea4a544;
assign I8922487573e02d684a3d71448c3828f5             = Ifd1431230378775456efa4bdd5bfc397;
assign I73164ee0df8db9282850f1b325afc7ae = Idc6b6357741c9887a9db1037ccc2d922;
assign I68bb1f26f878862f288c1f57049cf58b             = I6f0cef6d870e38e5ba192463a3920818;
assign Ic985d004f7feb36aaa6415dc7365e617 = I21e72a7e5870151c3247d15121e5fb4f;
assign I848ed394bd4f0b199d11c0ff458394a7             = I3ee87c05f23571b687611fdce84a1b91;
assign Ia09ac88781a570aead25d43447ff9afc = I10a6c6a8fdb0003de1f360c148777d0f;
assign I120d597a80158374726e064fb0f099fb             = Ide521f7523b897bb6fb747202f730ac5;
assign I17cb6dfd1374c74d63862703fa6665ce = Id806a2df1c4519bbbe811791cb4072f9;
assign I1c85c8f73ef80a6808c6aec0c8eca8ab             = I314b64e5fbbc14807fd7fe3c7bca101f;
assign I6c05d39d4c7a50f019474562f741e591 = I472352e7027b9df2fa957d9fd68443ff;
assign I50383e3d7c172eedfa00aa50a9faac4c             = Id5ad2e12b160bc6a9f96f2524f849c8e;
assign I413638a340bf1e686e718453f1b243b6 = I74cbc0ec3bb682e0f927890eef8d7a58;
assign I4c971e714427664c59c6371e14781bae             = I2b2bf6d4e879b8f53b02f94f1e964344;
assign I904a05d4a23c6d15438654f937811877 = I4cde586fc28f8d03fc9934d56f7ff7b8;
assign I2520aa556aadf851f58f0b1820498730             = Ic60cb038b4b90d8035059b1e06f8d765;
assign Iab36b17e472fde9a92c4dc5ebb75ca6c = Ibd59d0e5a062f149bd0e91ba76985a13;
assign I524e78ae6a4204e17ba4532dba047d4b             = I707e2d6d9807076bfc91417fb9e198e6;
assign I4d265ef808b1e19fb1dcef26a6dd4204 = I51e14ece9ab6607f83e6ba27f3f046a9;
assign Id1fbbe0594dae272856566522633bb3d             = I49f5797b92e17562e6dfde42c20c7a37;
assign I535542d9580a449d24a712ef814d5e58 = I433dd5092cf1851cd196feade3cfa6d8;
assign I432aa7cb844286c442356954f8814260             = I0a9f0274dc61d574c40e0e2048fb0b9e;
assign I82298047310dc4da0ea3762c6a48e07f = Ib83a067fb08e118dcf794902beef9405;
assign I6203f49a08107f7185ebadeecf2c16b0             = I53ae3de5769255a9e69a2ae690d44ba9;
assign I761dfdefbc96fec3c2ac79f0a1de18b7 = Ic4c6f707f461cebbc4c93f2ba664ae7b;
assign I4e8ebc46bc068c3f9889d970db131112             = I1390f0ff082dbff11a64cdfcbe1b681d;
assign Ib68e4d694df8e44519916724104f7962 = Icc67656ad2dd3fffae4e5abe02f8fff9;
assign Ie1817cbf3a80dae435a5571dfbd2f5ad             = Id2f8816659d3881ee1b1d14668a53a08;
assign I3284ce21b5d114a7127917f8b261b21a = Ib6124faff821158c6a2c9a9c454ab68c;
assign I92678f5b52c9c55556ff7f17f0f607b7             = I286bacc5a8a77b89cb99dbb00962555b;
assign I30b857065185101e8e4cb0270e747cae = I358cf9609272a4562423a85f9b2f56bf;
assign Ia706fb593b63cebbee0321c154cb859b             = Icda8e8a6ba7607752ed282114a542b67;
assign If9be63889327fc1b68abc628c9a0a78d = Ic04828ba2db8239b093043c27476d345;
assign Ib75747cb32130d44b338ed8c8af8ca11             = I2da4a59f9a6bd71af95790a75b172df0;
assign If0c3ec1e3a80a23b2506621ec2d9f02a = I38352b363fa37f6f822fbc1a39100968;
assign I43493f70f0336453d77caf7f27503daa             = I1bcf01b7fde13919f5d7c4df4483e61c;
assign I2842882109b7ef022421ab185471ab33 = I759409e242eaeb144a53e630a8cfd514;
assign I7fb3b66cb48521f8715f66bf5642cdb2             = Id5f000c37734979d057f7887739a5615;
assign Iecb13253abbfb0a891a4e526f05841f3 = Ic1e9d9113150ad57954c0e369259dc62;
assign Ia4b5f2b07556629673fc6576bc49a5dc             = Ibccd7142ba951dadbeca13178458bb3a;
assign I899cefdf3938be01e93d011e046c1e49 = Ibe6b8c57d7ff47b6fdad5fadf1f6b841;
assign Id1659ccdeaea3e59eb2d3f65a65ebd05             = Ic1fe6b93bc8d517686ba430d3d1fe7ab;
assign Ib96a9bf253b178aa920a63c8493932fb = Ic9b72b2a91d951cf08cf54ed215ecaa8;
assign I9ec9f389d0489908d497487e44c6edcd             = Ib1c8d1d733e91f052f6d6824e734b1e3;
assign I5f534382562a3394100cdadb3ad1e0be = Ied19cb51636bfb029ba8a2c390f97105;
assign I6714551e8885ef5e4490673fe1b2dad1             = I08348d0a177e264af1a4769422878a06;
assign I137e343ba2386bbe31813bbe37e87dd9 = If7fe3f5ccbb5b279e41fd183c8ff3974;
assign Ic532c6b85b156f821e0742f47239a65c             = I2d2c2997dcc5167fc6ddc1e90f0ebc49;

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          I3c62d5bd891bd3750b7bd1d32612f589 <= 1'b0;
          I699819696b0299ab80e7233d054ec590 <= 1'b0;
          //Iac11baea9832d6493626d2fe40fd385f <= 1'b0;
          //I92354deea988f3beb25bfba90735c6ac <= 1'b0;
          I6d3acefe6d7dfb94a5d66dcaa1bbbb76 <= 1'b0;
          Ibd047e2643dc68affb5b4f25b82ded31 <= 1'b0;
          I65e382d77592c7d1af308d171b27ff3c <= 1'b0;
          I7d4dc5e91ba3d952184d90de12f67bd3 <= 1'b0;
       end else begin
          I3c62d5bd891bd3750b7bd1d32612f589 <= start_dec | iter_start_int;//I3931f8f1df3ef8a71a54685fd9eccd76;
          I699819696b0299ab80e7233d054ec590 <= I3c62d5bd891bd3750b7bd1d32612f589;
          //Iac11baea9832d6493626d2fe40fd385f <= I699819696b0299ab80e7233d054ec590;
          //I92354deea988f3beb25bfba90735c6ac <= Iac11baea9832d6493626d2fe40fd385f;
          I6d3acefe6d7dfb94a5d66dcaa1bbbb76 <= I92354deea988f3beb25bfba90735c6ac;
          Ibd047e2643dc68affb5b4f25b82ded31 <= I6d3acefe6d7dfb94a5d66dcaa1bbbb76;
          I65e382d77592c7d1af308d171b27ff3c <= Ibd047e2643dc68affb5b4f25b82ded31;
          I7d4dc5e91ba3d952184d90de12f67bd3 <= I65e382d77592c7d1af308d171b27ff3c ;
       end
   end


assign I43864225be03ea8e9379eb28dfa6c599 = ~I5f68368511b59d2e365cc91b806b334e+ 1;
assign I31cb0c699cffcd2fedfbed0e1b86490e = ~I71e4d98dca37256fcc84248a26d703e2+ 1;
assign Ibed5004d869a01005768ba694c2234d6 = ~Ib8380902ac4082f834744ddef6d0cc6a+ 1;
assign Ia4b2db3d48f946b0bfd0be0e32d7518d = ~I9570f8498d95bee230bb3c5e720bb857+ 1;
assign I4d908bbe633c193cd9fc93dd33c60bd2 = ~I55c425102db0a6838012a165c0597680+ 1;
assign Ib14733d3585dbf7f196cfc068e9508f0 = ~Ic970a88c435a85d21ed71c6060b8a8e4+ 1;
assign Idfcf7f3240d92bfc87d44833bc00ff9d = ~Iec8dc328edd6cbaa2d697e05ed222746+ 1;
assign I1cff7306aaf303bb3342ea3d72048908 = ~I16d2084ccfb102c3bafc701872f5ef2d+ 1;
assign I26bdcc44692db066911c8d5b0a1aae0c = ~Id680a9affed622577164b3a8380494f5+ 1;
assign Id144785da9b171f1e2d0e9182d693e31 = ~Ifcd68be4bea38622d2d57d3a4e6fc5bb+ 1;
assign I6b7a8ba12de5b44817ec99faebe54617 = ~I16deb9107193a3536979e4b5e5654b9c+ 1;
assign I4a403449a9ba75243369032e1cca1a0d = ~I28cac65a4db3f708cc90a1b023bfe894+ 1;
assign If85d9a95c1c02ce2da1dc3486b53eb81 = ~Ie763738b7faf253837e1c45de255cb5e+ 1;
assign I8e470b68bf35c647af42b6e46201e570 = ~Icfef12499b53cd84f0aae067f30c17d0+ 1;
assign I484ec87270fcc959a486ebce40a9a03c = ~I0982b8d7f99aceb8871c9c10448f54c5+ 1;
assign I079932780612fbce79cbe9b58bb6c2b5 = ~I6c661048307c23c699d4b3636564de0f+ 1;
assign Ibb157b97546cb19fa7c1c0a7c79b1d38 = ~I786dfcaa131b99c254aaff15bd2c2b6d+ 1;
assign I45cb51c25c426c296f97a5d23a08c063 = ~I2b49d74cb130542f2ca99534e2c513b1+ 1;
assign Iff1d4b06901796098f91e87a3c30f7a5 = ~I0f6cb7a5a31d6f2f6178632c0c898bc6+ 1;
assign I16db9cab1981451a02dab21e2ca221b4 = ~I03bea609a189246a2375b355df47cf81+ 1;
assign I72756ea6a4997bc4afd4bfde1dfb2d26 = ~If56555b7cf539750706cf678030ccdb2+ 1;
assign I2882ae2eb6d79a5b96d1ed937dcfd8bf = ~I94e89b3a841f9760e3967c97e86d7160+ 1;
assign I1a632a3e06ad738d5865acc77e204f48 = ~I8cab6f6faf0758f26d1a8851fae43896+ 1;
assign I4d4ec5540257040d10182ed478a71918 = ~I6ecf7249e6151477fe74a79d0b126b21+ 1;
assign I8da7e01f56dc9a70eb6b3f110dc005c2 = ~I3753b2c4ba8f1bee70def390a96586b0+ 1;
assign Icc5d7bcbd7fcdb5092e6d8e18f6de6ec = ~I9b919f3d4ee3f33506b87bcdaf2d43a3+ 1;
assign I83cec264bd378f1dc23f87e439e7310e = ~Ib3be128b6704cc04c61e0fc9814dcf20+ 1;
assign Ied7e494fb288f78d110ed06662f1926a = ~If365a3c3ef86dca7c7315b91298c2db8+ 1;
assign Idd5b362dab4f93bba0c39af78c4c5981 = ~I83560e8d0f8cd37815cca6336fb2208d+ 1;
assign Id033e7adfcfb0420cc592a1fb6c297b6 = ~I099441ae3d3dffe49b18bc578af54dc7+ 1;
assign Iaee91a5e94c3f174682f72a1ebfd0021 = ~I58f89947eead94b5054a0fea3520ae33+ 1;
assign I0cd8a6e719305ee3fbe8228081993957 = ~Ibf565bf1803ed43120fa54b80f6f1f29+ 1;
assign I9b8cfdb69b76453a3ac687a1e098417f = ~I619957528c630e7f64924a25127c93fb+ 1;
assign Ic2159627df2efa5e677fa6f4498bdd31 = ~If3cc31fd16469339470702045fc6d0da+ 1;
assign I59fba74472ded0a985cb237104ac127f = ~I338ccc17dc6158aec0129c8b0c02c429+ 1;
assign Ia526539cc0f844b802d412b7a17cb6a6 = ~I83d71a89f35eb73265ee3e54184e1277+ 1;
assign I5d80b7c7d102d2c2bfa73a68c73376be = ~I7362f08ed4e4ae309dfbfda112c56ad6+ 1;
assign Ia92defa0ca87c7c30fbe901da40a575e = ~I8be4be8471625db0749e6385f87d2dcc+ 1;
assign I8fb1602dcdcd2912ea8aec42e2b7848f = ~I3d6a685a1913bd8be01fddbce1edec2e+ 1;
assign I0cedca0e2c589104d6f3318505910594 = ~Ifd77e040c5f82790b1d5636a42fca602+ 1;
assign I54c260db5c1b2c76527c8fc1cee229fe = ~Ifbe479e5cab3cba43444bec1e12e72a0+ 1;
assign I3d700e050cb7f22b0e381f3c72a20124 = ~Ia784f35a5a46837b69eb048dabf84052+ 1;
assign I63c0c8bef1dea4e499a16ce01e781951 = ~I8d0f440df332ea96e2d56eec490fbd51+ 1;
assign Ia8abcb8cf8d9ecc17c27ff015aa0b71f = ~I8d431a0524241fa54cf6dd1e79de4c74+ 1;
assign I3f59174b3764a0b0741462024be9fb92 = ~If49f97cc0c42b23ce393b534015559a0+ 1;
assign If0c2d002c315b21e11ae776bb48c9338 = ~Ie932a22a7f1fa37087cbc9e8d73efef4+ 1;
assign I18e548b082364c75686f2b7ad2ef46ab = ~I2956687a5fc2fba7149889624ef85647+ 1;
assign I5e0d6b44474a226ab2ce916a6d46072a = ~Iebf28886bd39c2540c90e808a9c20d3d+ 1;
assign I0c53d8d6a5b92960e29fc31cf456c23b = ~I8d4f3e64c8e3b0710a4a6b30d27c8be8+ 1;
assign Ib16c6096ce80e2f15a5ccea145e28510 = ~I16e3f3a6802fd206654bb622fa1393fe+ 1;
assign I0e7ca2d6470b9bfc6a1ca6143b468507 = ~I4b5713aee09999592256c407d4b8a95a+ 1;
assign I4ba05e74c2f63e2f4c59268775d549aa = ~Ieb1dbb98d5e5bda5b9ce803857f2ca26+ 1;
assign Iaed26e1c4a2578d16b111d15d31339d2 = ~Ife1c8d014675240a94f1133a78703ed5+ 1;
assign Ic566fe27ccaf2220101cbc49fc187a6b = ~I94d9412a7b43fa0bd4b9a6d32d313fc7+ 1;
assign Ibf9f6d7baed9e761b69fb41442761ac6 = ~If13e359e530823319046ce20027445dd+ 1;
assign Id5b4ee69444e5b499476c05a7f1d6e60 = ~I221777352b48c4e228c6637410113854+ 1;
assign Id6105518ade80c89d4f20222a2382efb = ~I1ee46fec2b82cf8e5142f8e2ac5d9d8a+ 1;
assign I26cf25e680483bf4e556d74efec35ee7 = ~Ie45aaf966aa0a94803050b5f43d69e6c+ 1;
assign I8636f5c91b567780d3324e4b8a320fc2 = ~I88aedd7f52399f5fd435c3415f2218ca+ 1;
assign I914bef0326cf82d350344317eb1359be = ~I7651176b0a74846108fbaabc5cc4900a+ 1;
assign I7de222bc26e38b8b6543819701740302 = ~I57ac487adc18165136e9b3c7c50f95ad+ 1;
assign Ie3361a270ebc41698ef4651bb3548a49 = ~Ic95668328a2121027436f682bac50b9c+ 1;
assign I1240c9410b897a4d0504affca5ba139e = ~I118726375ca9381e45f001965fcefc5b+ 1;
assign If17b4f86674bc5fb212a1f7751fb043a = ~Ic8d47ff5d6c31601a57df868da78c2d4+ 1;
assign I275f6334127640b2de3f0f87f54fd74c = ~I7cdc5ada6fc68ee31fd4062e2ff004d3+ 1;
assign Iec844d10736440b96f9d6c651e604efd = ~I59547aacdcfde31dc016ec2acbb2f4b4+ 1;
assign Ie04ce30f26a4ef1ee5b34474368dbac7 = ~Ia7f53f0cd86055da72c13ac474f052a1+ 1;
assign Ibfee0b4ad5cdf16e88fcf469c5e031e9 = ~I915054f2fbb8b93516d8748a3e3e29e2+ 1;
assign I3a4a965f22487553dec2a3e8e7836264 = ~If257757fa31c2f4cc9ec322e4ecccf83+ 1;
assign I2a2d014f94d7a3b9fb3024a3e9107a73 = ~If91268e2b84df18785cd6a53e53eb4e9+ 1;
assign I5bab5ae46114c487f67b8e779d7461df = ~Ia072f1d679429d3c3180f8eb67fc7dd7+ 1;
assign I45373bff54eccf8137da2931d841934e = ~I91a8168d3b087ab3891cd6d479427b95+ 1;
assign Ib9322ec1d3866ba3cb42e96b5ff5cfb2 = ~Id1dce8c1542f1279badb381aca3c9b51+ 1;
assign I0a9cb91319cc0d0c1c4d0020cce321d7 = ~I8983f003c30a218543f39f5bbcd9a25c+ 1;
assign I299b37fd45c6ee2031fb2c74caac73be = ~Id1b5c33bc63f75561b7cce6fc0981c69+ 1;
assign Ic2f450f7ab60ba57dfc1406c92c0f077 = ~I003f95fb8f2027efa41a1936e8b53986+ 1;
assign Ieca5b21b91e150c9d509964bdcea500d = ~Ie16dc913f571ae73ce03d755077345a9+ 1;
assign I48b39ee498563e23c3a4be079b6100d8 = ~I86e53eed5b857c439039238bb486067c+ 1;
assign Iac8cb32c2d86b975f51a2ed605002e51 = ~I89433799cfa534afd66e8d6b9f1b62b9+ 1;
assign Ic989dc794ce4356856b3916ab1889589 = ~I80f2e8f6743e28e86e4d85b295e2f768+ 1;
assign Ie380b37a78242e6d45b659d568887457 = ~I1391018fb93372ccc2fcc08700e38b65+ 1;
assign Ie43a7f8082f91c2955076a6373028b55 = ~I8fd26d47ecd4cdd08294cf6133468d17+ 1;
assign Iea765ae5e9c65b3186445b15c56f69e5 = ~I7097c9518bb3351818b96f31ed49c6d3+ 1;
assign I74b55d2f94073ba8f948e4b02386867c = ~Id683d693cd50645c3d6d657aa1c8bdb2+ 1;
assign I015630502f5cb4eb27b2a673e810f1dc = ~I88bd8012c93dd9e2ed52ea5e9b8b0004+ 1;
assign I5085f161323433d8d38be2e4511b0c46 = ~Ia8d3667adc34b2b50acf7edb970538d8+ 1;
assign Ie9fd8f7dc0c3849c0437a2a3d8607b4c = ~I3f0bba472e912f11dea8e788fbc1cb63+ 1;
assign I9306d9ef7934ffe5902306b9783c351e = ~I6dc671e73b4e9c70cabfdeaac2e5c40b+ 1;
assign I70e68beb262fbdeba621b3794adf9f84 = ~Ia6255a136d5f36ea6cba654bd5823850+ 1;
assign Ie7bf11bab3d601fd0a6e3eb415e263c8 = ~I2b9584392ef9a7828ff57bd4c522a302+ 1;
assign Ica3d4ebff001fb6ee69a66eb898eb5bd = ~I6c1235e88ae444a96ea64fd1bfd04d8f+ 1;
assign I27951ef3d612004abdc639662807426b = ~Id09b8242c22851fb960d55222fe733d4+ 1;
assign Ice4f4ba8bb3381c8846941d5d5fe4534 = ~Ie355fa27abbc41291eaf08f2cf9a6ff7+ 1;
assign I223151b6414d9979d71023053dd3f5e2 = ~I566224393f6bb27bfd8b0b0d6b8e53d6+ 1;
assign I73d2731c1b1ae5ef73ce0eb9c8995912 = ~I8fcad6e7d5ffc9f79eaaf634f6fe8cda+ 1;
assign I5ca15c7da1f49580ddedd9ff8ba822c0 = ~I6f0f74dcc830fdcb0af9df75a2b722f7+ 1;
assign I8289bfc08a5d8979ec26825bcb6e3d18 = ~Idd95fd099dd2b53c46d02f09575b8032+ 1;
assign Ie3c88bc240576aa220f0f110b13bfdd3 = ~I0f277bc88d46a4e6e9f1f2c410b503fd+ 1;
assign I583c6d23506c7d7b84403bfe977ec1ec = ~I66b92f1de2cf408c3af53b161a6ffa60+ 1;
assign I768afe193d9d79b136736abc6846d945 = ~Id28d9545e8d20ac080fbac5e345692da+ 1;
assign I277d7065150714e33d8ba64875d18190 = ~I4a5cfd6ebd47cda4fa2e06ba9ad6e5b2+ 1;
assign Ia5c77c9be26d62b026f24ee5a5e25fb8 = ~I62bda8dc70e0b5eb38abe094bbe92fc6+ 1;
assign I88a325547ccfe4eabf90792abd60e356 = ~I223b05d94c09b095d1988df121aa5e37+ 1;
assign I21842d06e25948ef461d1fd03485f86c = ~I5f73e5faf1aca83ee0a415c9ac4a1b9a+ 1;
assign Id65f22fa8fc9c47bfd00c796b63c9fa4 = ~I75f9d3a41019dca3044a1c2cf7069662+ 1;
assign I288ff69a7395e74f7de8da5a6a7f9062 = ~I820fa56328e3919970dd64adb1d4d8e7+ 1;
assign I2ba94ef71f97b9ba731b306d4a5fd02c = ~I05eadf11cdc6c2f2b021e33f2438fa49+ 1;
assign I26ae9e570a101c6f8237d7941285b924 = ~I2c487770d606451440eecf358202db32+ 1;
assign Icb92c7c10f0bfc5d287228f98d8a235c = ~I082aa8c413d7ef8f054b1c2857cbe39f+ 1;
assign Iba4972a3b71a3101ab23190ed905dc17 = ~I420e2c5a8745133f6263a71b458f1e2f+ 1;
assign I33703f538ec70268e6c00ad6eef6c4e0 = ~I4b8d520ee88fd39d83a16432e962f731+ 1;
assign I71b93abe4b20e6a17ff17e0f33ac2ca5 = ~Ia3f7f07ddb09ea33218afe14281ac3c6+ 1;
assign I91c2f3cdd7cc98a60090ec6e46d52ae7 = ~I25aefb53f59a00abe88b9dcf6be6907a+ 1;
assign I4254f2987cd014ed703ae18e9963e585 = ~I22c3140a8db02352d2e2a2a11eeba117+ 1;
assign I9068cca0de6ecff56ca542d0998fcab2 = ~I954dd66f60316803a8f13a39c460a39a+ 1;
assign Ib3ec015a3d43d46e0b7142b21a81cfee = ~I37b3988d699a1ed42923e3fd1584ecc0+ 1;
assign I8cb171677016e4309034dc5d83981a48 = ~If79bc5a35cb55036a367efb88c7d5510+ 1;
assign I2a4b3573ae7c3b38ec34591f20c1d076 = ~Ideab06dc2448a6950cd1a06a0c90c2c6+ 1;
assign I276c2ce5d3a1b7551c2790971071b094 = ~I1d7d7a68fc53b8be89c4637ac8f29380+ 1;
assign I9dff504e40aaddefedbb7b0f822c844a = ~Ib34ad1d14978608d1440f59998a31672+ 1;
assign I4ed5da534afbfe9ecbc10ef4cc649a55 = ~Id081512cd113e4d09df0fb13e443d76b+ 1;
assign I618363a8ac413dd0ee52eb658940eaed = ~I57a0f8c3710cf8e216d6dc2420f7621c+ 1;
assign I54166b387c02e12374d6febc425bfb7a = ~Iaa164a078c8cdaad694a053c9c1e0313+ 1;
assign I0b6cdfa1dbfa774fc9a12d856e61cddb = ~I7eb76b3d17296fdae702d8f820f1428d+ 1;
assign Ic4af6c9097257c9b22a57ce4b79b40fe = ~I00ecb5e329390023b318a2ceba0df231+ 1;
assign Iae21bdea20a6266d3f69aa680b6b2817 = ~Iea32ebc385c6cfc9212ff37973a0a05d+ 1;
assign I37e360420c7dd061de93a6647513676d = ~If845af0d620024f04525244753ba5d18+ 1;
assign Ia81c31ea4f4786136b539c9766987596 = ~I08e907b0619bec3ef2cf4cb3779e0794+ 1;
assign I5a4f0749acdc34fd0786e4b3d062f88b = ~I68e5b12792a86dda0576742831d3b728+ 1;
assign I5529d6db17b6184c45cc4487e5a2c24a = ~I72db05084d30d7c59ba1cb06d3b09400+ 1;
assign Iabe5aea929c668c9b9728d073ffb00c8 = ~Ib1f1aef6c0a9291553b62fd555feb2e7+ 1;
assign I4fb3fe065daa2708e55c812e57c19fb6 = ~Ib504b808f724ca6032e7c746517cd4fd+ 1;
assign I4bd98e902e805426fdd4606fcb5a5214 = ~Ia47f7fb27f2d965cfd2989569c257356+ 1;
assign Ia5e26c2417aba1005971749f4ab2f367 = ~If2b17f9e9186542117f43d0dd342326e+ 1;
assign I0e112f1d4e9c934a118f79f3856744a9 = ~I6c4ba0863ab4c8d1a56324a4d89ccbeb+ 1;
assign I005e8b590924f9486cb23191d35c9797 = ~I4dbd1bb8f1641f15e3a4f1e309962811+ 1;
assign I8c5f98353b5b082dc3cf056469945a08 = ~I26781ef851ed43c6f88ff1215cddca6b+ 1;
assign I9aa11f30712f1779339b985212a7979c = ~Ia349e1f7c10a63ddccb3f300c73b4572+ 1;
assign I65928407b1d5447dbc815cd2d2e7b37d = ~I50c4e1d3a3f63b93bc36b5141226fb3c+ 1;
assign If5b3850da967f6f3d7a71d680341ad1c = ~I12334038c2be8634c47869f397503019+ 1;
assign I0aa5522190c741b7df4c4d7d34e46987 = ~I64692d5168554dfd7ce1c7a046aecf72+ 1;
assign Iff777b2c4a3939e330c4cbb36cbe1ac5 = ~Ia4b438844530fff602ea04e72b07db8d+ 1;
assign I2d839c10960739097d449efab58b9fd4 = ~I9574759e112f27778f3645d5d49126b7+ 1;
assign Ice8765807beffd3acf59fa137ee0baac = ~I2ffb7c2ad09bac694ef13ec41e5de327+ 1;
assign I529eaa7e5eeb6d0a1aba78df5d5a2fa0 = ~Ib190f589f4d663dbc0a3c166a8dcf5fa+ 1;
assign Icb2805685607d5fedd0300c9d800f863 = ~I459c59ac61179d74170db53bf45ba89e+ 1;
assign Idadf072247b351cf51d718f797c3b375 = ~Ie5e432a991aff25577639f1b4ffd594f+ 1;
assign I6fcb3b133a6a654b69f41468a713d922 = ~I72064a6a84ff956d76a5aa590bbc05a9+ 1;
assign I77e1f5f504a794edbb89c66cf1ffcf66 = ~Iea74ecbac92e1b8f2ec7ad68d10b8e7d+ 1;
assign I185085cbf8da6df921ba32442b28bcca = ~I4f72d0db9fcc358c6fbec9964fbe0bbb+ 1;
assign Ibcb80df5bed66f8498561e3f3ffa4ec4 = ~Ifd958901d2ea2284f506e04a058012fa+ 1;
assign I2cf5304a672431888916e08b3c15f0c7 = ~Ie317bbd70b9092b840c0f2713204fb9d+ 1;
assign Icf266f710358631b7119ef526acb301c = ~I2f9e56d570e72714a06c59aa9e4334c0+ 1;
assign Ia209e5b03deaf4fcb8ae12b731a49e0a = ~I5b53fd45210b92703cb10d583f471ab9+ 1;
assign Iffb7fe9c74dfc01a43e99a099c4e7e04 = ~I8edbe77bacf1975e014faeee6b861980+ 1;
assign I43f52bcba1bd2e8ee5fac03320e4f19f = ~I174fcbc2ee01fc55edbc8238e5da7f0c+ 1;
assign I9fdfe73e77c384d33196c0f2d2a2fde2 = ~Id4dc304aef5f35f6ceb91796c278e716+ 1;
assign I546657528d591e8bb44c32fed7707af5 = ~I0cbdfae6f75a639eb591d9c0022f5838+ 1;
assign I6e4ae763dc4e8aa8afc4599de96c75d3 = ~I088898ee932a96c14f2f0f568f5455b6+ 1;
assign Id8c36004ae8e550569a491f6b514945a = ~Ide0abde3644a4fafb436aa59768d016e+ 1;
assign I111ac0aadbdd3e4479ca0786491a7b08 = ~I08581dc8d42be712cfb36d744f2786e0+ 1;
assign Ib83242b57ab050b0e5f9bdf91fa118fb = ~I29fb3830a5fc5922f1ec687a38941e97+ 1;
assign I7be8b2f8a9fe8e13001c2a1fce4a8a3f = ~I715d59fb27e519a9b76bdd8b5139a619+ 1;
assign If4d030e5858f325debc6f37abf4a7d6c = ~Ibe6a876a041198a581c95457a7d1fcf8+ 1;
assign I627e4bdc8061c69e3fcac17535b9f1e0 = ~Iec078a95a69b081cfb5e987ba9c5a613+ 1;
assign Ia443284a35e0873de59b3ae55b7f809d = ~I0e8f3f56bce3be1ee4d5f780a2f2a9fe+ 1;
assign Ibafedcf9f2990ed9c1efa973a0b1d81d = ~Ia73cacadbf80c0701a5b5b430c0d5c98+ 1;
assign I439c7c302b535bfd7db655c3c607d71f = ~Ic634d26fc09589a29a160e4efb5613a8+ 1;
assign I2133d362ba45ceb3dceaa84e95ace1e6 = ~Ie1374cac341cf353b1863dae9f544e8b+ 1;
assign I67534b68fee8f76ac0c5e64cd02aba42 = ~Ia07447985347e9a7f3739bd98867cdfb+ 1;
assign I8613cac4ccd4f956e8a0ae7b627f5be2 = ~I2121318f589878b4a9260625f97de518+ 1;
assign I8493e2dac01f009db1d2d5504b49d135 = ~Ibd8424c228f87f85df3da6204edff2b5+ 1;
assign I5c278aad08b7c4b0237d68f88fcb3f3a = ~I8a7fb51566bf215af214cd2fb5209974+ 1;
assign Iba75ff0f3b67c7e28cf627706733d528 = ~I7c0f872988488ac69815d288885dfd2f+ 1;
assign I9164fa2a9a33da6612ea692cf3fa7d2f = ~I3521b10b97b0e74888ce385cfc772945+ 1;
assign I0f3c4fb63ef1e88168b4d28175a0b68c = ~I58f0b81a46549cab8e74ecbc285df23a+ 1;
assign I99d236d41be79090ca7ba1fb6faaec4c = ~I7095040b38bf9d6b5229c11d2a0d7c57+ 1;
assign I487b9b236d118786e475ccc5e4e56a6d = ~I675ab6c4fb93b006f3fcafc985fbc405+ 1;
assign I6cb09ac924c3b3b44443263e08c3315c = ~I239a992ebb62899120a74b1c9e6cc4b4+ 1;
assign Id924dafd31fd0af0b28c7e6b7e95ec37 = ~I927c870d09285dcb47e6d399f319471e+ 1;
assign I9184110e3e9b8614460fc0abe5fff2d9 = ~Ie23ed3ee61f468f59f2baf661cb7f85d+ 1;
assign If8865fee7dbf593b34ea54692d947f10 = ~I68e58664be09261e5a80d6f8ecdd1b60+ 1;
assign I4854ff71aa885da3d07acaaa24740d7c = ~Id2808e0f40992c79ead4da7c734e5b79+ 1;
assign Ie8befb003fe83e774e8d1d01d4e2f4ad = ~Icb2b390266bff241a688961136db0f51+ 1;
assign Ie7e196fbb66ba6bee51ef0064ca519c2 = ~I54cfd68212d97a2cc8241ef429429453+ 1;
assign I685699f60c76b00df87c9c53e9a8e448 = ~I8d4e3962525c424786ae822a6981a5e6+ 1;
assign Ib6c0e635e659f54724737f0cffd1b0fc = ~I1a5f22b4e326d1684c0a8c7a7e754ab4+ 1;
assign I3a8bcfdab631a268d21c87b98e9d1c49 = ~I8c2e0c83a8204d6b21e0e3e458d56f05+ 1;
assign I3faeba79f7af7a006ab5cd256352e2db = ~Ie0622ff815747e4a9f368c74787026ec+ 1;
assign I02e672436ade3ee620c72c0d9ceee664 = ~I5ffed139764d90825b9f2eddacd0eddc+ 1;
assign I65708fb59e90bb79b8107da619fe63eb = ~I5a3297f48e1045273db6522744582b05+ 1;
assign I840a1a7c0bf49f4f42499b33f32fa02d = ~I9858bb2a3cc458aca5bf7eb077ee55dd+ 1;
assign If7543e2f5a158b1f3f3a4078ec54cab5 = ~I6e7e27bb176196e4493bf9c45ca19719+ 1;
assign I98a2aa729628adde0b6047869bd12743 = ~I4cff1804df738cbf4f940c775236df9c+ 1;
assign Ibfb57f2b507c27759a3556759f23977b = ~I0c1e22375d5e023c24519901b92eceb5+ 1;
assign Ib20dec1346f227042c749ec1abfa4d39 = ~Ida5b16851dc06534844a0b037d74feb3+ 1;
assign Ifba318d4faf308168c5eac8fe92395b4 = ~Iac3cb5b4481687fcf430c8bf52cfb74d+ 1;
assign I95b923444062b4a98918c685c65996d0 = ~Ia1499972c4995268acd828c1289f353d+ 1;
assign I45a6ef43e6e42594444adcbda26700ab = ~Ie559401a3a913400dc5e3e5641297fa6+ 1;
assign I508cea40d87bec2672f980d145c89b55 = ~Ie0667fbe76244eaec0b155d69dcc9447+ 1;
assign I0ace1d51fdee91f8f3826a945c4e66a4 = ~I1d0f031e8ae9c0335d501d1565118220+ 1;
assign I99ff3922e018c409dc8ce5f3503e3c56 = ~Ie2c801b2de066c3218d7312615b7bfda+ 1;
assign I6a3824a6598bbaa138e1e763ad85f5f7 = ~I64c4bb0d40d80ec52aab61ce46954f43+ 1;
assign I283107989a436e2c720123b8d9e335c2 = ~I512f57a40c7c8cb2f040bdde73e44ca3+ 1;
assign I7b12345fe53174cadef6811fb8869b42 = ~Id60cbf534604e5dba988050ef5abe625+ 1;
assign Iac6fcccf3a0cfe04edc0d998b60c2681 = ~I37998a91d20db2248ebdd8e661d42f70+ 1;
assign Ic9678deca4bf44a7b99f853334f6a05c = ~Ib65ff82aff398f6ff7ba711a36f41ee4+ 1;
assign Ie40c90fdb38b3e4046ba89295ed77d7c = ~I3d1dd8b9c7c6d3913f7ac369ad7e625c+ 1;
assign Iea4a7766d3b9d5d030ade1739859ef0d = ~I097722547450582dc5776bdaff914741+ 1;
assign I844b9a89ffb7a5e48979fdea546e244a = ~Id4a213e494f9c9be0fd1a307e87c756a+ 1;
assign I656852be6f5b3542862e0f68d48be518 = ~I21594c8b0169efd7c2aa6cbc31f4a901+ 1;
assign Id6551b6b053952162b90792ab73a1a49 = ~I15022e1b349eee259d3567837283dbf6+ 1;
assign Ib7fde6a2ec1ff0a3af10bccf3012e63f = ~I1070940dc2ef6e8ee3d1227ec9ff3162+ 1;
assign I989091b3586964ab598f166a89279d16 = ~I8922cc37cde6ba132f632743113e42af+ 1;
assign I9785922874bba479ce4a9bf1759e2933 = ~Ia66c399023e500ed67197dcf236f5d42+ 1;
assign Ifbaae8b3da03911a4c96d4efdb9283c5 = ~I1171dc208d5db1024dc3f09a90c78ca0+ 1;
assign I77a54091bc2c3d9006ecb3471b94d8c8 = ~Ic28b148967a5b3d05409976fa9001ac8+ 1;
assign I9859b94cda465ceaaa5674eb19e94824 = ~I79fe46308b93fbb24245fe1c75edf4a5+ 1;
assign I5a7746e9fbb8c009f83ae57423296cdf = ~I3bfcd63e92f1949234ab1d2701dbb499+ 1;
assign Ibddcc2e26fba20dfe2a2d399be2bc45b = ~I5e2331edf6e881e9f3a8c47eebda0ac4+ 1;
assign I8dbe6497a8deabcc60783bfe7548d0fb = ~I4b66c202450986ef0df05e979cc8bc7f+ 1;
assign Ifef870b405335975988b58b2273d4e1a = ~I737daf208eccf95feb3192897586cdce+ 1;
assign Ic1f6842b4f246d624d91daa6ada10ca9 = ~I29c8133231cfda17668bbe7b692bdfe2+ 1;
assign Ibc8679379ddc43ee4bc508a1f577eb2c = ~Id9d56f09595e80d66c2ac300f7d1d972+ 1;
assign Ibdd9957b7f1a319b797c021933ff75d7 = ~I97e89a2ee18d2688d7c1a640318a1e0d+ 1;
assign I041f9455435bfa375395eb330a34993d = ~Ife123bf57fe693dabe6aeaa236c4e058+ 1;
assign Ifbe29365e7035c78af9f42902b0d303e = ~I0c0d844fe3b7d35c1ed6bd7cc4e0dc24+ 1;
assign Ic8759e2f58848b33082bd1b02acc9c0b = ~I2d9632ae6a0f3ba44c3da8f56ba3fedf+ 1;
assign Ie2e3d64640c339dc51512979dbd6a173 = ~I38cc7b117c0bcd5e3060cd370d710d7e+ 1;
assign Ib2c327648cce481482eaf0467e9227d4 = ~I793ddbf6a5d026a57ab72984ca19deac+ 1;
assign I535cad8c919a4330257eb5b4bed61b3a = ~I79458089b042e181e37cc44c06d08681+ 1;
assign Ib2afdf9534deaae465d99b7e377788bb = ~I42460fae0acff25fa2b829e39ddcc4fd+ 1;
assign I6eaffd980e4d77fdbda5e63bad9489d7 = ~Id3670a6f05d40ab69624544de92b9c64+ 1;
assign I6e4786234b286b12c83e06e93c628534 = ~I81800fb49855a4fd2737faa07ff15d29+ 1;
assign Idcc745602c4b7b34df9c3d68f9a9d76d = ~Ibfe325e48511372569e0d98d9c4e70e3+ 1;
assign I0fc42ce9cc31d781ea3013318c25a571 = ~I326660e98f61bb2ced4c23c7bcc9324a+ 1;
assign I4363ca6b3d9ca9863f70958aa7c23777 = ~Ic6fa98631d742b27f252fe7c95caef55+ 1;
assign Ic902e09b33db1b919c102f7971cdef7b = ~Iab6d0f72579687407e029c630b107f7d+ 1;
assign Icf4405d4a4063448a2be8ad0354ab1a8 = ~I19eae741ef89baa1a64c403fb29f14f4+ 1;
assign I72108531a608f6d5e51a481c68d7b271 = ~I749b9c345f23aae03c595a2c76126ecb+ 1;
assign I6922b510e432e06d209095bcc6297e7e = ~Idc77c7d5123717fc2596a51d904c6d82+ 1;
assign Ief90f8a8efca2b06eff0d4cba1cbb342 = ~I779da979707d9712c1626d6025f97599+ 1;
assign Ib5334df42ee8f1574e41cb30b903fae9 = ~I97aede8502e443f98938487a5a5c072c+ 1;
assign I535b29f7177b4fc009ee998f1f4f7d7f = ~Ie7820d1a242bc28c19ec32d2c91e47b7+ 1;
assign Id0842da8068ee88d99af7acea50e7b77 = ~I82a14e1ee4723e7d9a13c1f2b8b13691+ 1;
assign Ib6cdbbb765694d822639b7c8fbfc50c4 = ~I77a94cd9186ca546ca9664942ea3537f+ 1;
assign Ibdaa6d215d34aa0cc27d5234da6fd991 = ~I3c0ddec25c53c166d30eb78d4518840e+ 1;
assign Id769d4a92f5f6da262ce0521e5509368 = ~I98bbe3b75958f10195dee6460cf2aca6+ 1;
assign Iaf3a0b5ea5d9eda47fcced9260922bc6 = ~If6d436031f68ef587750c5c1dfcfffc2+ 1;
assign I03a8a458ee0942c35001cbfe8e589222 = ~I461398638cb8280f1779915298540b00+ 1;
assign I25eb943ea517a4827efb1e797bfdc4f5 = ~I20c65000bbc10299168af7390776a03c+ 1;
assign Iac4b8906947fc90bfe76cee2f1d4c4ab = ~Ia840e19ca36795a50ab1a6e6a1729edb+ 1;
assign I58a490344f87b4d5bb319e3e85ba9278 = ~I7d98d1e5f07fccff5f20eaca6363c700+ 1;
assign I9222c4c0eb2b110fd80547d46ba17036 = ~I97a75b8625ae2a143cf364790ae77753+ 1;
assign Ic1af7410a9d11c5324f3ee5b2e0e9dac = ~Idbea892c8109117f90b453efe8ae25af+ 1;
assign I9e0a36d0be66b4c02b03e5b75b686226 = ~Icfc1c6d96a3598af73e99a350c387d72+ 1;
assign I1eef40a71c8d1e2da9802929a5347e90 = ~I523e9b6f828ec7f166750112f8a3f676+ 1;
assign Ied41909cd443432dafadba42672151c1 = ~I79259217f63b2f6263552c434d0e5c93+ 1;
assign Ib2c1636a66f6479d6123a038cbc668d5 = ~Ice6db5ba70d3c7499df6723a2df56bfe+ 1;
assign Ica02d19b129c8b1d491ea4747a55113e = ~I28aa517220bf597cf898660f698ef19d+ 1;
assign I31bf4597a3b776962f5c820378254065 = ~I07048dc5cbe24ff72d24902d572face0+ 1;
assign I58361fb97f1b5aff0a2751d35c8da672 = ~Iab3876e5107e3a56b1fafe41e16d9482+ 1;
assign I8ab7efc436a0f2cc3efbc299a0ddf914 = ~I511a55c2f4d6d3727dff5825597f55a9+ 1;
assign I3934ed7170967ff3852944cc39ba1de9 = ~I2493237a24acdcab8b5bda10e804a5cf+ 1;
assign Ic690477b1672dea4905a5e1c92b47366 = ~I03829256e357ac17c7ca7cae2f980f41+ 1;
assign I5eaa11e26f19b94dcb7eaee7f09d24b4 = ~Iae32c44b88fe7ddb5d4f19cf8fff3ba6+ 1;
assign Iaf1d3be13e6441a7a9ab3f286a7dc21b = ~I3bdc5ba374f85dc61346e4868c41a6bf+ 1;
assign I61f5ebea2bbe443b644c95ee559c2234 = ~I557ef77ce931535467a07a8d70145f55+ 1;
assign I1fbcaf2f6be01b129ebc24dee8a65396 = ~Ib4695d4389db72c5ac7e31809072c290+ 1;
assign I1c0df8c2c64b688ae417a238263f33db = ~Ie81315a3a14a5ef879d8e3f405936365+ 1;
assign I4f169c2c8c0768f2725ed655a03acfc2 = ~Ia7520053a7c4a94437c6a780b03a28a5+ 1;
assign I96f65790e2cacf7b529ce5b88598da00 = ~Ic308a5413f38b96d244cac3b0bc9462c+ 1;
assign I6b5720d71a0b4cd10ea34affa6631a25 = ~I034fb3850485fae2d1358041a1c41888+ 1;
assign Ifc7eec6765af08463751db128f8818b3 = ~I0e7079db66c15210046b997f319ece89+ 1;
assign I8dddcade21ad3bb330c1c25970c32b73 = ~I9a5388f8aa6e9924a309aa8db4c1983b+ 1;
assign I74a7b85ddacad06ab1c6b0db9b084bd3 = ~Ief76663994991118b1899ea4ddf4527d+ 1;
assign I2b0b168ce4fe8aa4a2e7cb69fe532aa3 = ~I6fb63ea54e492bdbc6d1145affc683e9+ 1;
assign I3e8d26ea83937cae01aadf1092c59bdf = ~If83ce1cbe3a73472419520c225b288a6+ 1;
assign I90a4190941651d885d04deb86a163365 = ~Id1df78ab32daf524b77c0431c782f2bf+ 1;
assign I7d85b73e85379bf3a480e954c05516f3 = ~Iff142b88493149045fc0de355b767c16+ 1;
assign Id5c9a9b9c34c8f9d56df0aa8d780c9d3 = ~I28c3818247c7c6de11790f6692882b5a+ 1;
assign I21255a0ad20a9668c958faf68d53b2bc = ~Ib451127b69a0a800332a712af77c6d29+ 1;
assign Ifba1584d599da13b98a3b76b4db10974 = ~I3d601db540da359ae4d22f960d3d5af8+ 1;
assign Iad0f4602ec545dc6ef12aa34add00ed3 = ~I2c1f2476efe593829ade470fe8ec2526+ 1;
assign I8bb46c3eb9f54c5d1b28dc6aa0154358 = ~I7e685b06df8a8c2ac351fa9f9b76a81d+ 1;
assign Ic09b4671e867144fe9f54a09e74c5519 = ~I1338d211b5d2d409bfe0df76d2ca2701+ 1;
assign I391a2f354262558ff17d7d80b8c39e8c = ~Ia40dad546d9c852e2fa8942c62a1c1f8+ 1;
assign If6b40a030cb120fe017bf9d39e1a35d1 = ~I0b0dd019d8bd24684403a29aed668b6d+ 1;
assign I490996026af34eba5bcd8d553af818eb = ~I66a304016a9adfd85a2abb6f8fd39afc+ 1;
assign Icbc12ab47f586b12402ae5d4361c967d = ~I177be24718c59688752097fe2a4085c4+ 1;
assign Iee0e45914c52a357e1e32922299d6937 = ~I7e66a42eb7cdb820cd1297c39f0625e8+ 1;
assign Iefe423653d454e21324a6857b52f98ac = ~If2021f0735c6c5649ebac0d230fda87c+ 1;
assign I6d6a242cdfadfc97fe656510bef73adc = ~Ie1bf5d97b8f679095d2442bbf9f95608+ 1;
assign Ib5c8d91204a2d313c9c23110a53cd0cf = ~I632469889d6bb1c268b45fb805467ebd+ 1;
assign Ic9740baafb1c92e3a25f0a1e7bc46486 = ~Ie230ba3c73808e102eee9e5868595e7c+ 1;
assign I6f69796a6fe6da57066319ec8210c1a3 = ~Ie1e9326e4eee006ec07abb6bb7d269a5+ 1;
assign Idb862697f62a6c678072de760e176096 = ~Ica4ec1647bdb5a3aad6db6b447bd7995+ 1;
assign I06e05a1ed002175a75d02b8b76f52c50 = ~Ia17295aec0a40c2b46a595dacfede2d5+ 1;
assign I1e110e27162231650875dd1152d96e64 = ~I4c6d3d6fc2d10066a744fdd9405a7902+ 1;
assign Ic46357bb77f6183329946f7e28294365 = ~Ia9c043c5e8873fd13e39cf6bd8136c51+ 1;
assign I8741c5cc763512d16cb1186fa3323f45 = ~I2e802c75c6ce34b05943b678ecbfacb1+ 1;
assign I30b5c7aadb5312ce96e833704bb3a320 = ~Ieb3f28762410fb40a0c8a8556b4b3ca0+ 1;
assign If404a00ab81d6ebbc0dbdf4aecdce389 = ~Ie3e0c0e40c7a67ce7f957e74bd2a895d+ 1;
assign I19875f52f79482b477f1febaa7e97090 = ~I491f2373b2df19a4c22e1787ef034179+ 1;
assign Ic7855ca956651bd368cbdde7ec93ba6d = ~Ief96603d41b4f670d2bbfa3d3875c903+ 1;
assign Ic57a2627a194099105a2908a41feddfb = ~I7a029c27d92754041eb6d605837238dd+ 1;
assign I4d1ba6ee8fb9505ba3b58b2b7553245b = ~I00dad36628d2fa923120fdaa79bf0045+ 1;
assign Ieb7b388ff89e352dd239e0ccbe7b9ecc = ~I3707f68de059df0af5c652fc0478e543+ 1;
assign Ib1461f456ebc14f449eee77e386a4c69 = ~I94af4b6b9dc11935db54ba872889392d+ 1;
assign I8786eb767f02164cdc32f14f41b5d0e1 = ~I38e2dbba093928b874d447362d89b291+ 1;
assign Id6fa8ec5d1062fc3e09bdac65ff79f45 = ~Ia48f0029e9e76386f3dd70aacd9adbfa+ 1;
assign I83b77ad1a40dc102f28153f692516eb4 = ~Ic2b20168744fafbe15037ed7fa83da72+ 1;
assign I55e54359961ef6e5a63f1c2eb0ad4aa1 = ~I62fdc8936121a2707d94cf3bd6e660ac+ 1;
assign I90001da8c360ccff128f637cd672ad42 = ~Ia0932b3fd6a5ae6da2bacd2b86ba3a43+ 1;
assign Ib38a46dc131d635b81fb7c196110fc4b = ~I9fce6091885f1bb97d29fb1f543b1a38+ 1;
assign I926c049036f53f0a0a6ad369de116c57 = ~Ib402cdbfaa9900820b85bd625415c547+ 1;
assign Iac48d2ccf6c6e0c555e874ae77123f2e = ~I518a2736384c14c02f27bfa3d8ea7aff+ 1;
assign Ic6f40833f5f6284c9015304fd3fc00f0 = ~I847cf7ff866f8a666872c12d6b67b1b1+ 1;
assign I3f2507530dd648814af0964f7da11d35 = ~I9e45e3d7117ce48cdbfc5db8c0ccfcf4+ 1;
assign Id9edc6ac95a260bf5af3de25f00e9e9c = ~I380ff8528cdba4026fac3c4eda8b2c52+ 1;
assign I28fa295ebd90c2b7255d48ca9ffcfcf3 = ~Iee8f9b0654f6f6797f11cae0947e454e+ 1;
assign Ia308e09137af1cb50167562efb5da628 = ~Ie3e54a4700d8d0f6478187e06cb6f85d+ 1;
assign I5aa85d9503b0e4ff46bbd63e873053ca = ~I8c0069e8756bcff203ce21ae3170aa42+ 1;
assign I7ea8fe50c45e213f3257060e2813240b = ~I856eada207c5006beb8f83f01d5d74c9+ 1;
assign Ic3e6e38a2986c7f14fd0db2246367a1c = ~I79a46279070c53678a5af54f661c5821+ 1;
assign I581eb136fdd08302e02c1fafb5d5c90b = ~Ica807adc510a2e32580ca77c18ea0b45+ 1;
assign I080832c25509f7003ed50d71210bc7f7 = ~Ia8094903aed8dd0ce8e9ff459a5287b0+ 1;
assign Ib43383830037df764b48c637a28ab6b5 = ~Ie018f3003c5f124bddd13c359257bf35+ 1;
assign Iddf65ccb4396288264a400ba37cbb655 = ~Ice18bceb10fec484ffc96155e14c4974+ 1;
assign Ia7673d73f0535906a99d6cb467892104 = ~Ib484aa64b795f7e36198b800f302164f+ 1;
assign I8bc3210e86a523accdbeefe7e72ee4fc = ~Icdb143a4ce96029c2441758bf2edd7b0+ 1;
assign Ib63574478126e6ee30a388d9648cb548 = ~I3a76f70ca3bfbcacc6f3342aa71f1912+ 1;
assign Ic4501a8a1fb34c30a97e18a0ab189e3a = ~I9470c7ab9634c01bb832c9e4ff5496bf+ 1;
assign I2b807c16cfc6d65cb2a7f28ffa837974 = ~I218ee96418a4f5d734d3d71685bc09c7+ 1;
assign I0aa93075086164fdbab3814d60633141 = ~I924514226fdb5bac110a2650bcb2e85f+ 1;
assign I886750aaf8d2040c3f12ff113294f658 = ~Idc57f37015a48393608e2b026bc7065c+ 1;
assign I103ec7cf279f527fc6e3648a19a12a8a = ~I41af7e4c97fc04154fe6de66b82499f5+ 1;
assign I9a57f2f03cf8a154c3a7d48ec089306d = ~I972bee4216f8e532e8fa4bd25fbb9c57+ 1;
assign I9d8f8c1792427975a9e7024041f59be9 = ~Ib303ea0240e7ab5f000dd10e975b2274+ 1;
assign Ie8644d7edbadf19937c399cf275946e5 = ~I5971253546899e9a82f387d5eabcc7b3+ 1;
assign I2b32537c9178028493af165398a60875 = ~I1fc36e6f738fab96df356979e1e3a612+ 1;
assign If06a1563b9d7348de03a98d31bd85b06 = ~Ie2d8c84d8c9a4c8f637068a2ae39fdde+ 1;
assign I58a7c7b05b84d292cd06d68e96ecb9f8 = ~I114c595caa67a3f777f087a634130a6d+ 1;
assign I3fdec80112b3fc543b217d1c253406da = ~Idad14b6383b9af54eb35e72ff3d10035+ 1;
assign Ia1aedd38250e76763aaee3de2f832b3c = ~I46e9c76b19ed1ff21f102efe6ee5c732+ 1;
assign I2087576fbc15119bf5d9e8afa2603b69 = ~Ic75b8bbb1b80001ec188a0cd25623420+ 1;
assign I7a6ab9e700bd94208ab6528af413f3a9 = ~Idc7df6877bdb7e7d392307d78183d31c+ 1;
assign I4481555c402ba99bee05658ba6017984 = ~Ib8b95ece5da3877b261a06e6d0571921+ 1;
assign Ib849494e5087777f646ee0947b4f634a = ~Ic99654bf4833c9132912eeb4c0dc92fa+ 1;
assign I18d0dd7a10d6533f721a2392d4ad2d02 = ~I2461055ef9b1aa2ffca0f5cac3300e71+ 1;
assign Ib8603cb82ceb97c2f35bf8209306a457 = ~I2bc3ffbe5b42b0833206437d3863278e+ 1;
assign I2418ae211f327ed45cc70c42078180dc = ~Id5e02d4c48fa6c3b0d45a9e66f09448f+ 1;
assign I6521c9167261db6eb37f50b66159ddb7 = ~I40e99289d5762e77a3766eb8251eef00+ 1;
assign I920f95bb52cdc9b07f93afc3a6b5c009 = ~I20beb3fdbe91936f74a200cd8ec9817b+ 1;
assign Iad0ecc5208263d239e4a62c5563f52ab = ~Id435b68afb53bef4afc7b70a9512e955+ 1;
assign I0c0be3347a7df9cc39997208b013f17b = ~I0cf5cb4cd472502b84dbf6fe1af0be78+ 1;
assign I70dc03a46e1ac0da826388abd3bdc503 = ~Iacf6340a29a5592b61ea875304a2de48+ 1;
assign I452ba61d5fb5c7ead1824dade4bd7801 = ~I5dfc71255cba279420b7545df4d35c40+ 1;
assign I8b5d10c412daccdcb07645bf239d61bd = ~Ibadcb205c7e9a0f3345cac7eb41b5985+ 1;
assign I9b1390839ee2b9ba591e3873e967c8e2 = ~I762b2abb876381eff6de97cef0798405+ 1;
assign I17e818b67440efaba9a5d19e7467bf85 = ~Ib3e7633767b6e09e4ee54f6feaddd31e+ 1;
assign Ifa67d343acc6f3ec50c2b01fc26b4374 = ~I3f193e9c265c1dfaeada63d59db5b79f+ 1;
assign If0676ef300628c4097565b13ef2d8854 = ~Ie72268e979cf069b88f6eadde789e5ab+ 1;
assign I8d26e73fafa909f1e26e329828cf4888 = ~I5732fdb805258fc13c8ba4aaf56574ca+ 1;
assign If29fcea810adbdb1c4d8a4ace1d8081b = ~I3afe987d8f2c93cc19534a3221d1939c+ 1;
assign I0e3286fca6cd040758950259ab663df7 = ~Ic66af6c3c0268cfb0e9f0776c4f4e961+ 1;
assign I696db0b98e27dcc4657dc7feb23a881b = ~Ia605d14205926b3edc6d1c2f69f70ac0+ 1;
assign I06c0921675f464807a63c7965796f0d0 = ~I0071f2168787bd42ab7f2370aed9d0f5+ 1;
assign If36016df78d833c80e1355151c038225 = ~I4936f823841b0ffe32f801f5134c0211+ 1;
assign I0dbf900b4f430b4c1106aa86b640bb37 = ~I5975ef8f6cf53cf2132cdd9d707e7912+ 1;
assign Ib8664a2abe9d6326d6e45bb2a7ad59d0 = ~I954ff0f9ee871a31774a3d786128fa13+ 1;
assign I91893028c4409cfeceeb7976815b2d31 = ~I31f6bbfbbbd4c20d0c5c71663da1d4c1+ 1;
assign I2e14fb1e667e967ab4c116e0c7438aec = ~I1898bc3cc6a8b6f71d65c758d1f08366+ 1;
assign I0fb60c4f56f6d7b4007cf0dae39f4573 = ~If86532f849bd392dbf599eeb2fae0545+ 1;
assign I24b4c998d19ae97f7178e37f75c77d06 = ~Ia344734d285ac29b53cf401c08a0f987+ 1;
assign Idb73eba1bd4ce25a6109e296f51e7dc4 = ~I502a8e382aa0881dc86f3c13e0566ca3+ 1;
assign Ibc1a16427d8dfa5ee20dac15327a53ea = ~Ic462cebbfc39190b22d20013259e39eb+ 1;
assign I0e52c25aa840402d944cbd81f73c1ffe = ~I385d03def4cfb49f54867687ebd710ed+ 1;
assign Id7619819e1297844d92c8bf3a1d61926 = ~If8aa3ec1b5a4a3c122da82467be917da+ 1;
assign Idfa432a87877e1ce103e56891745b62a = ~I8daf79a0a2ee1bac7f055af441539fa4+ 1;
assign I13b9e098622d90a1074f636d8f351aca = ~I6261e0d339762cb2364421e6b87086cb+ 1;
assign I78e1205de9119fac3ae8f43c72ac71f4 = ~I0e2f746715b901feb69f6b3c94f3a828+ 1;
assign I5bbbc4eedb7c61516769f429a8498ea7 = ~I7b8da162c08f8aa2ae90522ee1526cf6+ 1;
assign Ia1d9dee7a9821283498d17de0cfacb32 = ~I5e8ecdbb018402b2fbc0049ee44bae8c+ 1;
assign Idd8643af2515f65fd9a1dfe66494ccf2 = ~I06d859184884c07a14c83d2f06587ad5+ 1;
assign I1684820afb9d9cec38cfdfcd6ca8b36a = ~I79e3e49f57d47231c0fe6aaafdbc57f1+ 1;
assign Ice8a82bdd966719098a8d5f2a826f73d = ~I12c07042202f66db926861c9ce7c2b25+ 1;
assign I338400586daa58006c0a3dcd82ea8f4a = ~I9d0fdb45b9e86bd409740e538a690320+ 1;
assign Ie467c5fde1d123da4e9587b5a56748a0 = ~Id5fd6f25dc3df22a322434ae3c90dea6+ 1;
assign Ifc52604a4f9f9de392a35f2f9fe885b8 = ~Id812a8ea2a3b4a912d151be582833fcf+ 1;
assign I20c4e393929b875521e5316f4d8e2d42 = ~Ifd3638d44e1ba2285891fac152dee327+ 1;
assign I064499f0315fbeec7b6cb50583388a07 = ~Idd1b6014de2f053554ed09c29bf3e640+ 1;
assign I894ef04bfa1b7b39ef51b7c82f7686eb = ~I0d96336eb4d5071d7e1d350e86513b25+ 1;
assign I8d6927b0bcbbb318cf52987c121a07b5 = ~I31e5b2cdc3dc571eafa37510076bcc64+ 1;
assign Ie0ce2826fd13b0e0b23c91e97787691f = ~Ia8849f78971a45ed0daa2489e7d27dd7+ 1;
assign I7dbd1aeba00bb8b257990b7bb294211f = ~Ie4749f8e9ad2b370f9f9814b5a463c43+ 1;
assign Id5ddf5331aba567aaf5b7eb88b31a52e = ~I3096d11098113da669ee0a94686e600d+ 1;
assign I0f46a17f14ab18e6338aa3d06678b0a5 = ~I09a1d04c307fcb8a0e30925d86df3fe9+ 1;
assign If1ec4241fd12255369f72b3f3310b6e7 = ~Idb0a98cea3ee6cd4308bfc2414a003e1+ 1;
assign Iedf37dac8b3a5331277ae4f0176968aa = ~Id4788855f9a503e8b506d012aaeea445+ 1;
assign Ia422fbdf8f318ff3ddc049d1374e7939 = ~I5b937934e7aae1f916c2848889f12685+ 1;
assign I9cbe73d708c561d43d05945552d32dde = ~I9275bb36e58e0f17964e13ee7f027ab7+ 1;
assign I7e36dcae438a712fca2320117b7e3356 = ~I02330ade2eed926076cc071e45eed82c+ 1;
assign I0f9bc36c9d40290f83489aac3d674924 = ~I296bc392d4223cbdd6f77be6523df819+ 1;
assign I3a09554ca009781e28ef1b3ea70d39ad = ~I31b0f2fe98cfddbc05dbd14be8be394b+ 1;
assign I28ea268c5b51ac1d9249e96599bb6b0d = ~Ia71663e8f563041c27cd21a0c9c27a28+ 1;
assign I1d648ed8f07f0743a6d616584270c513 = ~Ib46b13498ec14ceaa56719f26f18febb+ 1;
assign I82a225237aeb1ceb31e8cd18b1e45c6f = ~I9bc2d5692474b8368c570d92835191b3+ 1;
assign I36ed1a0d0d618f90443fbea17b7c97ec = ~If8b0b96a659183e3651c691a2848b86b+ 1;
assign I612a41511db375f10f3c2b10d13edb24 = ~I87d958c00fc6209d901147831b0c951c+ 1;
assign I19032091a26dfdfffff60818041ec79e = ~Ie4e4eaf3e5d2f581210af8054df71c6c+ 1;
assign I6aba8ca0e4b20a6355b43a70f19d9d8c = ~I0b557cf102da41afd26936cbdb64b6e8+ 1;
assign I839895c8614ff28df83314c44824900b = ~I49eb064043f91112c854e31e4eb9b885+ 1;
assign I8cbafa797ef136d7e50c909dc160deb1 = ~I1039bc43e88eee527d2ed6adb8c7d1ba+ 1;
assign Ibac0851ce1a3c23f18b072d263afff36 = ~I9aab16e89f1b64117caece8ca8af5940+ 1;
assign Id58474582f209a3859f65a447fe99191 = ~I343df614f97cf732e57cf2ad3f95dc9e+ 1;
assign Ic9e06a355beabfacc053ec48f17f49de = ~Ie02de90d8eb06b16314946d21299500c+ 1;
assign I77fd8001d879fc9e9117464fba27902d = ~I3353a7916b569f2c0ca122180608dccc+ 1;
assign I2a0dc4ed573a544cb13544e049514903 = ~Ibfe760474fcac99f1e5ffa2e008fef99+ 1;
assign I71bc7271cc432bb3c5d0b7a416cdfc60 = ~I3caf1211dcbcdc746a3e4c7fbbdae4a8+ 1;
assign Ib76e892d1a1271844338042381b5690b = ~I2dcc0d17b9fcac35693bf32b5c5540fd+ 1;
assign Icb158c031d434cb419c15e0510511231 = ~Ie6764a631310e312ba5c2c1e601d828f+ 1;
assign I563802213afb6abe2f6e8c6f4d1e5b08 = ~I220f8e45e5fe6e69f02cded87f12e1e5+ 1;
assign Ia5b779ef95333736b08f63770900e275 = ~I896cd566a3d078b0f697a788efd223f2+ 1;
assign Ic1120eb027841908cd64fe5c7274da14 = ~I7caa41076a293edf18c7c4309fdcfc91+ 1;
assign I5160de2c5ce4782d8f8be10dc740694b = ~I928a0e4951208aab170656596f456209+ 1;
assign I5f7b6e6a30348ae86057f7e56f625846 = ~Ia3d129fd297905bee180293c0c39d9ef+ 1;
assign I9de41d0b279b84366640880dbd18c502 = ~Id555c88cf7f0904db74d45cc75c8f5d6+ 1;
assign Ifec9abca21cf476b70e0befa3926b46a = ~I1ddfd31bbf062aa5c3c71d61e492e3a2+ 1;
assign Ifc527b6af9486df7f52d7eb9637c671f = ~Iae9e023628eb6686708b2656f15616cc+ 1;
assign I31d94aae2e3721045fe850d84dd2225a = ~If4b100d26126e460c41b8c1bc8fbbb96+ 1;
assign If3bdbb4c20efca0c5af78614b4271ed1 = ~I85a7fede715578be0634d71e9c7951cd+ 1;
assign I4037f1b207aa101f354e59eddd7c9eb4 = ~I2d7715a3af03d9664729fa6df85034a2+ 1;
assign If4d63635a5f99c4dc9e5b57712830c20 = ~I571ddcb0a10938e4c0816c965214b4a8+ 1;
assign I1f1f2fefd3381ee48ab0ec9c9301754b = ~I8bf8b0cf27a2654a0e7fdf3255945b67+ 1;
assign Iba52b84e6e215842e0ca8e72c42ebce7 = ~I63f82f075d53205b5b556c0054f1a0b8+ 1;
assign I597c3f5c14e235f90dc8c796bc3e931d = ~I3c6fb0df5846a19228a4e6cf9f9106ac+ 1;
assign I397a69dab323c7148b620dd6fe0b0c51 = ~I7168b0efdd2fae57292379c9d15c62eb+ 1;
assign I401ab1ad994f5018061a3f57d3a51ad1 = ~Ibe502ebbb366f54a8f8fda4e361308e3+ 1;
assign I3a47540f34ce47bcfa1da66cc4e6e088 = ~Ifce70fefde8f5ea4d2c1857236f66d65+ 1;
assign I18916d0023ca275d84c52af07dcc5ca2 = ~Ice2c390d296e09b117d60905343e9098+ 1;
assign Ic79072d9e42dbc9974231f1d642b3f12 = ~I4b94402a53d981e953c21ef316c709b7+ 1;
assign I1140fa91b5e22ba0c094c03295781e5a = ~I450c0d6ad5d3b1f18bb28e3a432b5442+ 1;
assign Id2989aaee3930698cd374e6c9feedf82 = ~I2587a5800a5a9ffeabc4dca503e3d964+ 1;
assign Icda9a86a25dbe516a93b46fe487029e3 = ~I1182655739d7ab5bbe4a6546a5ca36fd+ 1;
assign I53971b75cbd7ebc74b579776a6ea4778 = ~I8110a5a62607093b21b7cd088b1d9ee0+ 1;
assign I37e5c3118e8536e37bd797aeaa92476c = ~I8b611f7c12ddd81de403ba74e212857f+ 1;
assign I9c68bfa3b888b6a6d41e38e674578284 = ~I84a62a133dbceb5a32a7c907f371663d+ 1;
assign I2c72d6c5fa6968dffa6517cf81219875 = ~Ia2fc8a1bbc3cb0dd7d89a7f05b04909c+ 1;
assign I9bb4d58b1fe80549451b00c4ed2b3885 = ~I2a3eb42a4402e873d081f94a14a99c20+ 1;
assign Ic488e78b5c73251b673301e84c4b5b0b = ~I58447d6ae49a6be2d043477a06f83df0+ 1;
assign I8d07beccef519ab4ce4024d911ac2346 = ~I83292bcda4645233d8e8a1dfe8e5f60b+ 1;
assign I7c191c2c2be09886d0f31e4368797afd = ~Ic5e0a84cf1a2ef907b2456559ea26c75+ 1;
assign Ia3bfd86e26efbef2cf6bb72be7ac1453 = ~I2cefbf897bb7f6f67ca500727e85c683+ 1;
assign I4ae59dd2f57bda295e11b077e8668f1a = ~If47be2ca4617a426258c51f8d977ba3f+ 1;
assign I3f6fad8bb0fba790fcdb1612b6fa7712 = ~I7c68e0ae30efc4ca4d68b6047119c6c3+ 1;
assign I58416287b268462d28f55c6c2705e613 = ~Iccca1936f4c1c9496205e77b588e9985+ 1;
assign I106d0e71b7378d110b0a624e5cbf0d6e = ~I59d4567d3355fdae5660a1364d1b8d00+ 1;
assign I59adad4fd84c1fc233dc58f70a12779d = ~I4600963866dcb9bbea2515c805f885cb+ 1;
assign I8e01532a1ab9534b8de0474549d41a2e = ~If26d90629e70c5a871e6f5b14471b8cf+ 1;
assign I80af3dcb716f3474a7257700aef89b81 = ~Iedb9bb14951bf67bc8865b0983490c14+ 1;
assign I07d68462362d8453e83570cc793c55db = ~I6a3854ed571e8c262aa3ec377c247778+ 1;
assign I9a2bba3f62de5f750dc8161a488dc331 = ~I05028975b49ec0c089bd981696f85a8b+ 1;
assign I71da7e172b2b967040b6e6d02ef9949e = ~Ife732309efcc740cfff5c747aab2e3d6+ 1;
assign Ib97b2670a6cd88b2327f07f62d887900 = ~Idcef10a0465614cf38e0d6f503b5174a+ 1;
assign Ib2963b82260024e1853d297798d88d3c = ~Ibd4aaf02982068ffbfd1b8b3795d9217+ 1;
assign I0722ec4e9d400f8eaeacd060e42de79c = ~I788c64785b992c675fe348a1fa181525+ 1;
assign I1972375d51767f0cffa5395a354b3493 = ~Ib235af5b28d56f24372d3f0af816f2c2+ 1;
assign Ifb19d75cfa0051107b5fba57bfc002b5 = ~I4c03a6569d1b954d088053e38827e811+ 1;
assign I9d05dc0e39e85c23b62f343a8de12e64 = ~Idda26504e422367082caeafbb29871f9+ 1;
assign I64ae3cd6f36b8bde29cd3e1fcba7bade = ~I195c3a82123142d509886ee37dc6fc98+ 1;
assign Ia6a78664c080829664158f53ba330312 = ~I1abb512ca0383c9e7104418e07281841+ 1;
assign I2ba16a10a82c20d54c776a9804ee50e4 = ~I00ff1331b1900bb031ee81d2a58c1bd5+ 1;
assign Ie9a316de516ec4fb828a614c67e38b2a = ~If65eb5e743a7b1878fb232ef2fe13cb0+ 1;
assign Ie945349d77442536992d9ad52ce84218 = ~I24ae7de3549a84f4f88f561b6017b7a8+ 1;
assign Ic6a7a82d16e6106071934ba79d3698cd = ~I449c77140475475b138d839a74078337+ 1;
assign Ide40b1bf9c0b642c49a5685a62af1c93 = ~Ia9e102d8679943c079f16c0228f0f0d1+ 1;
assign I79280400a4c9bed015106e5d006de757 = ~Ibf1c9d86665f696d91c554db748ff42b+ 1;
assign Ic6e3847f035738243f4c5f71f296da57 = ~Ieb0336a1974a2aec0966f4f59f460802+ 1;
assign I45b64b2b963963d2d0a8318133941f1d = ~Ic0819ccefe784a6379716b3633ae0196+ 1;
assign I1939152ddbede923cde577984e0aa743 = ~I0c4bbd1827b1859caabb067e864ce4b3+ 1;
assign Ifbcebda2bb0ce58a0e1764c392a816df = ~I004c98da87996b77b5761d366210f782+ 1;
assign I6d0d098e6d47dea04d6d7be67b648a0d = ~Ia457938da4efe847cb06f645f2a54a52+ 1;
assign Icaeb9a2ec8ec5822658fa85b88cca04b = ~I7e0474089ebc1c34747be1bc17a81d72+ 1;
assign I3cc30aaba3dcd3eda262a19e85e53117 = ~Ib0b46b99e61d724ae664d9d1fec1e29f+ 1;
assign Ic0b2f9717b8aacb34325fd5aaf03a366 = ~I56d1025271f1f7704a40dd7f0df02b0b+ 1;
assign I002869e450d79649d27441ce00bfb575 = ~I72c2256ba47cf03f95143df8f741fd83+ 1;
assign Ie4d20df6b1e7a42f0df9a3cc26b12ac1 = ~I733c3fa4d84e5680792b16a70bb1a51d+ 1;
assign Idd01d014f0469f893305057ae3f4cb2e = ~If367d63311c96726517240de13bd2a4b+ 1;
assign I79444eef1875b6ad1a0675b66392ff9d = ~Icc6d895d943e14f2801c22e79ce190e8+ 1;
assign I7caf8c7496dd96c1ed08e98b415f5775 = ~Ieb664ac9be65fba2e25960141f7fb4b6+ 1;
assign I7fc6e2aecff5bd691872d1e10a39103b = ~I66071f20991b414140869a2e3b750471+ 1;
assign I49321308413cb4dbe5e6c01ba5b9023c = ~Iffeefa89a2ba7d032db5db64cbf05e20+ 1;
assign Id27560fb44b4f2fda98d47e9f20d6898 = ~I9ab3cea6ee8d8473221da21bae06066b+ 1;
assign I745187336b8a5ae4eac66e90539752cf = ~I3403ce6e697b523a9f441d8fd5e2d420+ 1;
assign I772e844c41387e7079259875e0ba3fa0 = ~Ia98a70144e466b356d2998948dc4b602+ 1;
assign I32c35da92922c5b477f8aba837fa6d92 = ~Ie4ca0836695d951ee09622892ee35928+ 1;
assign I3bc01b072987a0c980615abbc2251e5f = ~I485a48b4ff4da08f977425fd10e6d392+ 1;
assign If08adda7d796da7c7849e472a73282a3 = ~Ie8c79e6a5378808c0ead5a4b24319ce9+ 1;
assign Ife3bb8945e14d8746c82b66886293997 = ~I9ca81c841a75a9ac242835956509e0fe+ 1;
assign I45ef0ac486fe043f57e8a46aa91461a3 = ~Id50f18f642f3b00ffa34986f78a0eae6+ 1;
assign Ic0ae1191869e636f9e4391efe93309ae = ~I75838ca09e301b8e1301cbf603a1f8c2+ 1;
assign Id92d779518ae724b5fef5221372f8f26 = ~Id968b34075e351ab01d65abcb4ed8cca+ 1;
assign Id0762ac7710c93249bc11c6ce4ae51a0 = ~I84da4ce7441e132e775167c1cd81dbe5+ 1;
assign Ife6be241bc50560a14f97650e5cc2959 = ~If19dc22d45cc4664c85a043ec4c00617+ 1;
assign I1062442edb2bff727ca6283c8270bf28 = ~Ibf482db0f5058be72061267c42ebc292+ 1;
assign I6c9ae8b8191507f908c27bbde53bf2d5 = ~I6d2dbb953a58b91dafa7f0d34d41bdc3+ 1;
assign Iec936eeebd1f8c95307bd8705e6def81 = ~Ib393146d81d3cf031466543311cee2ad+ 1;
assign I6332af145d560e3f22a4a88106749f98 = ~I42564ec6a794ea803795f0b5b3523a93+ 1;
assign I0c121fa3e9e6e0e2e8291a594d6b4ceb = ~I4a0033a180d7edce81fcfef603532e28+ 1;
assign Ic3c59a5167cb83fd76ec6236572b1f3d = ~Ic7a21921e2716fba55aad2e351f4498a+ 1;
assign I3e8e280553edaa5c8555ace81ecc10e0 = ~I9a3f0b4867087790c78f674b719dbf7b+ 1;
assign I3e466d40a4447a23953d96d2e6d61d47 = ~I138f008a6206a1067bb0e22ce3d90990+ 1;
assign I76e4c55148effeba62a4837cd19c5e51 = ~I48ad9b737892d7c49340ed679f46e034+ 1;
assign Ie335e68643fd2b0a53351f4bd45c3475 = ~I04a9c9765fd468a7e841577f09fc287b+ 1;
assign I89f75107ea95f207b9e664a1f4f0746a = ~I7b929c228c865112f00bc6b4dcc95b52+ 1;
assign Ic8f0049e1298b14b4e039075dc0d5f74 = ~I2b54a135e59945901e9c11580a29ee3d+ 1;
assign I382153cec6f7d6258574e7c532186473 = ~I566221060f06e724676ec9bec861d7de+ 1;
assign I351dc309e916f282cc1e19303eee4112 = ~Icd9a876a0feb16ea62bcad5be2004dac+ 1;
assign I9de5e90485b3f22e9003dc8a7b22a79b = ~I8f8273c4cb2a9ace8a09847efd4bdec7+ 1;
assign Idc4171a40dd2470e852af37a461013c7 = ~I96ef4b631a7f63e19f67f3920685f0e6+ 1;
assign Ifae488cb68d95ea517376319eb11f1bf = ~I9e2de71442b8f504358e582087a6d19f+ 1;
assign I9cab38b69794ab661e12750cf69c822c = ~I1fb13d7500f5ac3821c424bd3688cf4e+ 1;
assign I24180fba17c21bacefa8a4514e4b685c = ~I2aabda12ff89e708d04b4399472b5203+ 1;
assign I83bbe6fa947f9f909e1a6785ab31901f = ~I8c733a5d394e6b8d045eede5cc7451f6+ 1;
assign I202c385beeccee309104b66f8f096b2c = ~I4f45dd50d2825ab338b8a2a8264096c0+ 1;
assign Idc549661d6694035874a3366704801c7 = ~Ib45caf6b563d22144be3e9225a99a1cd+ 1;
assign I778fbaea65beeb6de599490daf3b7e3c = ~I9d6730140c690037b5ca58aa30103f5b+ 1;
assign I4fd45670f88265e5d7aa6582f3ad3ff8 = ~I9df5b63f66c162d517daa69f5d0e6095+ 1;
assign I2d636a246d815a4d12c478794860dd40 = ~I1b40adfd6fa6c943dfa8d230d9e65514+ 1;
assign I3319313fe1d2b4ec2626711b187b4a5a = ~I0eb3df4d4094e09e6c4b3c788baed61f+ 1;
assign I586aaa5c55efd37996b01febd3bc60a4 = ~Id6f7923a16cc5adc96a730083153ca6d+ 1;
assign I95ccc219b5f5038641b38dff6db0b222 = ~Idf8ebc0d747ae143aa61866e33d458c0+ 1;
assign I5001118df37d08bd19d322aca8ff3996 = ~Id682e531735437bc24abbf3d3d51e18b+ 1;
assign I22c15857572603cc24d8a87cb47c33b0 = ~I05ecce409cca00ea5b0df25de5a50cf2+ 1;
assign Ifdcd91f925b63e0817798aa6e9200e50 = ~I831d214dcb4f8d534b5ddaaeaeeb81ce+ 1;
assign I8435e69bc1ff06e7edfabbee7b9aa49e = ~Ia540866403683bc30504bace19bdda7b+ 1;
assign Ibeff607ba15fd8ef504224a9c1d102fc = ~I05fb1982415bd3fa78dd9a00af7a3d4a+ 1;
assign Id15c3bdce785df234c68432ccec8f959 = ~I977864efb0d94149cce7dc4d165f11de+ 1;
assign I25888aa2135fc403ca9eac4df634549a = ~I9362b615a612599239e3b752a9334e8c+ 1;
assign I632ffd09a9091335b3aa91ab2a8f1cce = ~I5d4fb4b5a5ad3dc48beebfa0e0cebbed+ 1;
assign I283331db80e6d0891b13dc55e6a7d76c = ~Ifb9b29c43f435452cc761218c509f5df+ 1;
assign I134a734d93e62f6ac6635015fe3a2096 = ~If2143db72bf9a02b64eb45b3a4faa39d+ 1;
assign Id66798f8ea67e74a67f264fe6b4503a3 = ~Ice780b1695a8e80607a03dee3c426ffe+ 1;
assign If2ce7b8d2573494564393f7d426fa47f = ~I90b0296f5ef87dfaa6110fc2e9d6ed9d+ 1;
assign Id59cf860d9f4aff11b205b8970d93df3 = ~Icd37da8ea84a606529e32b2db4eb7f5f+ 1;
assign I75aaeab4f372e28a8e51453540f9c6b2 = ~Ie626a24e3680f7d3995dd0c2ce60cbcc+ 1;
assign I2266afbacf1ba750ce18f296aba1181d = ~Iebee55168fb47664095b11c9f6641124+ 1;
assign I69c2b063e61e14f5d49b907095ece00f = ~Ic0954671eb1dc893c3932e456800fadf+ 1;
assign If077c67a062095cfe69f2260cee82833 = ~Ia4131464996aabab8aae1db85f6a50e4+ 1;
assign Ibc03a9b6115d0941ce9233df7ef2fa57 = ~I2de1ca2c390bdd3011fff4a359bb5332+ 1;
assign Ia18bdb8d2f02b50281f0acd4a45ac973 = ~I6fb55222b69475b7168874423226ec9c+ 1;
assign Ib88c884e54d6e6ecf5ac015bc304e4f3 = ~I9b09b800a9dcd8ac36f25cb0324e748d+ 1;
assign If6f5efee5e1f9709d86bf28cfb741955 = ~I74ac0327175f50f508a5013df298df02+ 1;
assign Ia0caf6693d441ac622f416a86b665166 = ~Ica26f542586d50c56ce0f3c00f36b388+ 1;
assign I85dd6a9634284c22027b4241551ea628 = ~I7c6862830daffc98cb2c1fc121d82c38+ 1;
assign Id5cedaa397ebfc2567efcc2f8a648db5 = ~Icf19dd665616a8c96146b3ab9f46c741+ 1;
assign Ica0a119af1728ae253c16cc3eb93f802 = ~I97f2813ec39bbf1513faf66b3e38838a+ 1;
assign Ie7274a7ffa053ced4f12a67986d3c81b = ~I716ee53e79883f69aa045380a357e913+ 1;
assign Ife7985db888089ea618413810611bfca = ~I25c324feaca84e80f58075597e8c448f+ 1;
assign If49068db99aa9d09302eda27ab51fcb7 = ~I7fc190647082a3d71614f46f670167bc+ 1;
assign I2959f2dc554e599d675eb6912757e413 = ~Iebdf938a28594624f4d4a337356485cb+ 1;
assign I898d1b59aab3d5d4adce8ec3c0e14a0d = ~I3fd068d55154441ffd005999ea823fd0+ 1;
assign Ibb6e54edb9d277242c06d386a9a75a26 = ~Ic5ca74b66763c6e5591c7c2bfeeb0663+ 1;
assign I51b1cd475d0e389326b182cbe680a402 = ~I5ab556386d2973354a5551ba9823e4ba+ 1;
assign If12366160fdc899bd71cb0de5bcfd84d = ~I64f65df774d29696425ba460dda09b68+ 1;
assign I44e5ce0cdf812c5b73e6e638da36e414 = ~I9e09c25be9f877c1e1aaf79bf12c7943+ 1;
assign I4f38c3d620b72f21cf6d54c7df4ba816 = ~I42c1d469ff97913cbf15e3ebee6fdfa8+ 1;
assign Ib66b897398ea0702b74bdd03774f3ae4 = ~If9f2a53dbf6e9b9a335a7657b7a2b468+ 1;
assign I0b3a936c3f7e0391111e696b2445803b = ~I495f8be463b15db906474c518e0741e2+ 1;
assign I10f045edf47784a91a5599494c2d3de2 = ~I3e265a7dcf29687248b9275df49771fb+ 1;
assign I6a81b4485598387e4656c35e83866209 = ~Iffd94cf3a8a4681ff3327c90bf89bd8b+ 1;
assign Icf7630b6002db2f9b59d5323d6cc8105 = ~Iea71417e738c6ca54c50aa014cc38627+ 1;
assign I3db0adb3457cb22c755f5d29a8fe7ed8 = ~Ic8df04756f67e6dd29f3374c5f86d451+ 1;
assign I887911fd9466f4d4fa7f50642d610d88 = ~I546122346a22ad64a6ab2b4978cde095+ 1;
assign I9ae284c0089ae462a1bb9d168bde2fd0 = ~Icaae0fb0f460f68d690ab00697355a49+ 1;
assign I342a563de39175fe4a6eb7e3e1ccac9a = ~I42455e7e4d0c63f97702d204d18a446e+ 1;
assign Idc758f8e6fabb6b31b0a7d9c0c590310 = ~Iaec2f15665e83416bc140890f3cdde9a+ 1;
assign I72b4ef48363856af7faacc85eafbaf2f = ~I487391402b6aa27bf212724a37ea9c33+ 1;
assign I4ae2f2330a8ee7d5626499f2a030c7a5 = ~Ia9f375709014a9d553d46cff2799b59f+ 1;
assign I4aa98503fc71292d42dba1cab6db952f = ~I34d428a56bd0142a9be9f627f1c3c87f+ 1;
assign Ic35d5ac4dac46d47b2796bbac6452161 = ~I57db98eb439d59a895dabe029c6a3a8b+ 1;
assign I32679702c19eab37b46d13bb372967ea = ~I9937af6fcf9d834f308bc3683d524981+ 1;
assign I6a86b03402bd2e35208d3fc74601f9cf = ~I463f4f370e1ecad71de44780eff10df4+ 1;
assign If8a259e0c4f1839e852abec6e1b904ee = ~I53309409a6059c3bd39f037c23ec3458+ 1;
assign I938dd59e4cdf3434086f60d000113430 = ~I2603e0b8b93f6680e44c9c8883f6512c+ 1;
assign Idc198bd5732ca5760d1a700a25273ce3 = ~Iab354cc9ac1173335c0efeef694f3567+ 1;
assign I9dfdffbfdb83572cc3205f674e5db753 = ~I6c19936ca2edeb0e261e880a1055e964+ 1;
assign I60520c850a95b893528569c4069bd677 = ~Ifebfa58419ecd22a334ed4b67f5c3581+ 1;
assign If525ac3dc97e3187e036d70e9984939d = ~I71a28e8525f07dabeabe4b4f45f353d0+ 1;
assign I0c1e4d400520935c5c78b792a9d554ba = ~I514830acdad20c4ff3d078477e939b4b+ 1;
assign Ic7d5fe6c4b1dcb97d10ba3de2f95d1df = ~I036342f6be0f2e2f1f4927099a5c4a78+ 1;
assign I8efad9622c05177563ab8a2747879044 = ~Iedb655aa25e5f0e35137ec6c3acdc527+ 1;
assign Ied4ddedaf801fbd7238d8a55c17c8090 = ~I0c59e8c82a31aacbf5977ff778a7ff49+ 1;
assign Ieb9720b6beb2363d651346ef0233cd49 = ~I1b6d20c64b9f23fb6c30f723546aa285+ 1;
assign I202aa0814e7e28a6bd21db116b652b4d = ~I0d66aa55747362354aa81d96057bc4c2+ 1;
assign Id201f81bbd80a70006a10866b8efeeff = ~I1ea33707e40a2e41513fdb3118371437+ 1;
assign Ic227f42a20219c6638ee3343ca445acf = ~I68c85727adecde0aa8aa66ed08c4b502+ 1;
assign I507e9bd0265d9ca6cd21a46fa21ba084 = ~Iebd050e29044153d5881ef80b2db8c28+ 1;
assign Ie04e44d8e0756cdf34cf9ad53da76e47 = ~I3c057d64cf4fca0238a874f0ced99c76+ 1;
assign Ic92ab3dac1a151d6ff0b4e0c21003eb0 = ~I066cd52173ec5dbce9a3f470d73325af+ 1;
assign I3da241c7f221413abfbf1b4384bfca5a = ~Ic7ad59f6a232a997706d17b4098e0324+ 1;
assign I0807a826e91f92ef279ccf0b6512a428 = ~Icf8cfc800f0a2aa5140a7f83f035b0cc+ 1;
assign I05aabdf73200996b7bea8db700fa8930 = ~I6bfbf7ff79ff0a6facc9ba5031239644+ 1;
assign I03038b940be8bd21bd26b150b28754a6 = ~I78ade92efd265027807c861be44a10af+ 1;
assign Ibf547f8a5e1059ffaabeb3f447904dcf = ~I2bc5a10c587d89d10021aa5eaafb490a+ 1;
assign I2ea27544ba4cc14d0f7ccf7158a27a2f = ~I30080cc6c03bbe933165d266558a822c+ 1;
assign Ib2f34922b0d5346500de093275bebc94 = ~I7e28234bdf66ab5489d36d15678db797+ 1;
assign Id2e223005a932987b6f60663773187f8 = ~I74b3c9dd3a8168aacd4369b9ff68fdfd+ 1;
assign I3188d354c2ba494ffe210dcd89c00620 = ~Ia7046faae1ab05978e4b32bd44049fb9+ 1;
assign I09faa07bf38acd96c4e29afd8a5167e8 = ~I0c5250aaca86185fed5978438c8861b6+ 1;
assign I6d4867d03d9187e95e27e99f7aecddec = ~Ic78949e07e643f571f23df7e8f15d9fb+ 1;
assign Ifb09b84f9681c7bc28ffd562b633ffd9 = ~Ifb8b3586a5b69b20cf03eabf51344ab6+ 1;
assign Ib55b0e4c45ebbdb605f0ba9d62bff21c = ~I9ea09f27ce4484f2e7fc3a6b6d6ecb7c+ 1;
assign I4319fa23d59f4e690e31fb7e3a823d17 = ~If0b9225e759438be175c4128c78605ea+ 1;
assign I4ee3f608cc8f8df27345949f1a3713a7 = ~I33d941ad9d4858fcfb77f0f6cf99d2ec+ 1;
assign Iede5d56e52612e083407888da49470e5 = ~Ia0868eee7e7e0640ce1a4d3ca9c001cb+ 1;
assign I3b2739319710681986b9d3f8cd04f619 = ~Icb3ab2c67a87b2ee158e0021b72fc186+ 1;
assign I850c257a0412bd9bd6001817bd9d0ee1 = ~I5b64997d083769666741c794dd92fb7f+ 1;
assign Ib7875bf9d30d071e62a474c50d88ba06 = ~I0a3323aac825506435068f6746aee974+ 1;
assign Ia92b76ee5b7d82a992a1b58147c0c0be = ~Ibec442c099da091afcf75a7c970bf8ea+ 1;
assign I2253b32e46200a23dba243819fce02f0 = ~If3a79ede332c39a8d2a276de833242f6+ 1;
assign I1b01cadaac7d3d15007f0afe5c0ab0f2 = ~I49ccb3e14fe61618806e791ecb4f4eae+ 1;
assign Ie96877deef8b1676138f814c4a720800 = ~I461ebbf3a02ae63e2eb27531b1370f24+ 1;
assign I8ce945d9f70bb317064a8d2d4eafd2d3 = ~Ice66c108aa66981051df71e226cb0e4d+ 1;
assign Iaed105b99eae5b078521e3a94d8a79b7 = ~I645ff0d8c0a87ba7f792fc83f342b958+ 1;
assign I05a812cd935867d1e417c64c26ea0952 = ~Ica94017f26e96fb22a47add326ee126e+ 1;
assign Ic0a580f94f3d03f72e3a487f84bf6612 = ~Id32e7ad5b1aa825732d9b26d0fa02ca1+ 1;
assign I39d9044227c161f0163e58dd82aadc90 = ~I51b5e641856239367cf43f9b5679b268+ 1;
assign I5f607bdc9b276fdf07a17a11a20a6720 = ~I2d1a5645b126761fc7fb70d24e37189a+ 1;
assign I12e8b8cf609c2fbdc72efce9bb5dabee = ~I49f5f87662fbb540d72c94bfd1acd060+ 1;
assign I6fdccefd034e8b4b86cfa997502512ae = ~I30253dc91301ca27b5732312c01145e0+ 1;
assign Idcd5283cf7b42d403ee0e4404b5b311b = ~I143f5e324716a94d24ada126886bf895+ 1;
assign Ia020344403aad35e050765a4b0cc42b7 = ~If64aa8c220b9ab6652e081da7e404e80+ 1;
assign Id11fd3a31b70da0e64138e71840cfb83 = ~I1092325b801600fa7ec85fa640167da9+ 1;
assign Ie9c5e7c98281cd1deb6acc51590c9d9a = ~Ib028686da9c849e827cf249a744b7db3+ 1;
assign Ia0e77e9544481aa0f56dfdb6eb253137 = ~I5f3ff7fa8686f7a380302d71b88cfb4b+ 1;
assign Iec0d7ea31e0f1a75b15121090dcf1e11 = ~Ic01904f7c518990eff2dc1de127676c4+ 1;
assign Ia98bb3648ce3719b1c31ce0f41121c63 = ~I43f2ddd9780f86af489f8deae51168ec+ 1;
assign Id9c8055ef530f2cb8096cb7bb2af55a4 = ~I0a013fff6c792363bd7feb03d9691db8+ 1;
assign Ib9081d438413a627f5b16f68c2eabb80 = ~I7cf8401bf6893eab0b9f33a0f91ddd05+ 1;
assign I9c5bf5451736358f8c84e150004fa5a9 = ~Ic7ccbeaf4ab94d0660eb7a0533723e24+ 1;
assign I377933518c3807edb71f648c65ad5c85 = ~I08043393cb7f2558c145a698ea6652c9+ 1;
assign Icec98d794a64752081fadfa74308fad3 = ~I84865c4f872c0845124b78fabf695c2c+ 1;
assign I7bbe4d0a7d61d3f7da346de71b9a3a5f = ~I57b9dd7a7deea6695dcd03439c9723cf+ 1;
assign I197c05f74bf7fb8d44124d40bd7c6563 = ~I1cd6b35bcdfd461db69a4c1bdb1d387f+ 1;
assign I92acc55d81ec6e02880337b0a451ae21 = ~I40a1ecabded8add5bffe316f2d8beda9+ 1;
assign I35c0ca76b28cd2f9355276b5d2f29ad4 = ~I7c52ae4af926267b5e27a530202fcce0+ 1;
assign I29da0e5661f29bd8493c19885c998582 = ~I1a5c6c50817db8bde279d5f0b5095d76+ 1;
assign I9426c8c1b4d988d5cd7d89a7aed4f8fc = ~Idf0c1b85712fcbbbcc12915158ebff62+ 1;
assign Ibd010f15e36194cbd2ce9f01c98a2b6f = ~I6b32298e8c61e75d0a38bca3084c0528+ 1;
assign I7e86ab53e6d9647b230a94e076831ba2 = ~I5b0d72cedc120406402076148e2d30b0+ 1;
assign Ia0ecfaedbc1d546d484978fd50096d10 = ~Iaf624549f73b0d13c1a73c850b99f810+ 1;
assign I27098cbe2d4fdd634385d771cc290c2b = ~Iaaf7efeae9f6dc9e8222dc2b10122000+ 1;
assign I5d7a0739e447775e00115799c52b11dd = ~Iea1cd2321d2ac9b891b344e2ba2363d3+ 1;
assign Ie95793e09085b6de1383a37cc7fc41ac = ~Ia544fa24b953fe91800978895e3e610e+ 1;
assign Ib24b68cb35da39a743e1d90bba3f0836 = ~I7fa710c37f5f96c3cdc35612a702a71c+ 1;
assign Id4cdd72193e90dddd211af73d7f3634a = ~I98fd105696fca11c1075f9bd30013747+ 1;
assign Iccab4c19a9190689f90a42160e2379de = ~I61345963ceabdaa0f25f8a463fc9fe5d+ 1;
assign I275ea08a3dc0600d8ccb6300eb7f2a6b = ~I9e8375af6af10f4bac3e87e416d430ee+ 1;
assign I1b53098a7240d2b5dc1f5c5c3b4bcc11 = ~Ida1cd844022bbf1b8431225e66b2b78f+ 1;
assign I278659ca1a0b093fc883d01987989dc0 = ~I30e9ab592e97dbc5fb6ab58d2ffbf8d4+ 1;
assign If92e66cba66732798dd19f968a5ef8ce = ~I2ec2a6de2be39b1bc259b0be72e35a0f+ 1;
assign I784c4e9fb75c314f271477e0621aaf7c = ~Ic32e349efae2ca419e095ee5e15a501d+ 1;
assign I3d3aafdd4d9d3e9fdab1f487c48a0ea9 = ~I1befb935ee9cb871c9a7476c1fc0da3f+ 1;
assign Idb4c722992139f39914af7085378c6cc = ~I01c57f697f2af7d2c6ae904319f10725+ 1;
assign I63c9deb7e6a4b400e0aff6887a09e647 = ~Id580f8a2748efff9b6b747c497c16e9c+ 1;
assign Ie6f67c6e4c5e2b8357c0a902979e8722 = ~I77b54488bd26318f14b4364035cd1836+ 1;
assign I1d7a4f99e3975fd01bfe5a9a1da84765 = ~I786338397f55073dce91e1c8c5f8e298+ 1;
assign I059d847e09f5aa3f6a8147062f4b13bf = ~I0e5931219d94c8e8e1f4af081404dcab+ 1;
assign I48e5256ade4d061a3b5ba08a53252bc3 = ~I8d96b419b010f8076311420d7b9c8a18+ 1;
assign I635fb29c55e0fb5cff0b6f443c2e3de5 = ~Ife13f962c7a8df3845cde104a959f678+ 1;
assign I088c5b971a2def57248769a33b7d2a2d = ~I7f701ff37ad3fc34d2f4efafe5ff5351+ 1;
assign Ide22394fce1658f9e7002bdb30d03c2f = ~I43c815a8ce0b2df9744a525328969691+ 1;
assign I9ff276a14d3205b98174a8a736f79774 = ~I6c4a1ded9bf39091cf302ebe0103e2f0+ 1;
assign I123255637493b9c7924e3a72d1b86ee9 = ~Icd4ff8d14af2699db2b5168027894ebb+ 1;
assign I87e6ef84894cfc86b94e19c9d3065bc6 = ~Ia79d52fe2130426c07890fcaa50137db+ 1;
assign I4c32900878260a261bc5403e8abd6258 = ~I308aaa8ac500b5589aa4af533a9062bf+ 1;
assign Ifc100357ae3f754fb0e3863334bcc764 = ~Iac91f4037e542d9fda30fadafe7e79ac+ 1;
assign Iefe9e5376010997c0ee52eeb28e57a25 = ~I8cd5970682bc84881489c12ff073212c+ 1;
assign Ie6060acdcb16b6fa6aeeb649ed621053 = ~I1ee27be7e1a38aff0039b21c45f406d1+ 1;
assign I46c2b923860b0d1c01b9475f4467f280 = ~Idf90f01353ad1057e11fd060442f4e53+ 1;
assign I38b4eceb159ecb0dda3920290a21a02a = ~Id45f4e0f142b6c3925f24a37dcf7c0ae+ 1;
assign Ic45561ffe1837c3d5bb42c695a377f82 = ~I52a9bcfbd2d3a763671f19cfeaf7bb8b+ 1;
assign I3e76abc721bf7ed186f4d0f8f4bbf4e3 = ~Ia3cc6acf2cae41e560e09993007ffd2b+ 1;
assign I1afb4061458e9d2f5799afa1f2373bd2 = ~Iba0d2f08788f2208a648ae7b5414195d+ 1;
assign I18bb9a781a4c314fe6bd990e4c275f67 = ~I9f7df6ad60284c812aeb522974578e0b+ 1;
assign I49d7342f105c4502377abd23db973752 = ~Iab1fb7006598181bd8749ed90c519b13+ 1;
assign Ieeb12d463444ca36af1ecf2e09504c06 = ~Ieef3b299ec35075c71ef9fb10525bfc4+ 1;
assign I17525df1798fa2c1c4bbc4a1ddcdd0a5 = ~I58a7c08adf48d0737c5803e2a818c045+ 1;
assign I90c44c31fa7903a81826c1c568597362 = ~I30a1c8fcd9a510a6ed559f07dd809b90+ 1;
assign I3997cf122743b612f49cd5dd125a9201 = ~Ic4f5e9d49419e1c57cfa387761ab643d+ 1;
assign I1112c4267582ddb8148ee40d9529beee = ~Id3dd71ea0bf0f2996fbe42b8c3318762+ 1;
assign I21c207af859b94634d3750482b42a2ca = ~Ib834b91bf81067e8efa9d470023e8b9d+ 1;
assign I2ff2421bd86bf9ec110724460f1171e9 = ~Ic6ead78ed741442f17a15a157cd6ef9c+ 1;
assign I6ba5c453b17e4b33c61caf5d70041c4a = ~I4e257dbd6f196a02dc0f5a2e5f6047d7+ 1;
assign I08318099725fbe033ab8d5427eb8b278 = ~I3dbfbd34d1fdfd4f422d900154123b6b+ 1;
assign If36cb462cdf20b0b1758cd6417e524fa = ~I529b763dace1924613d184c6c70c2708+ 1;
assign I40e8463645b1122b7cb224770fa00447 = ~I7a600aeb6cf8c3311c10afa4d82767a1+ 1;
assign Ide386e751e06dd5df0c042cd76f0f800 = ~I8c7aab31f8cb705ea13a41a5bd349303+ 1;
assign If63bb4681bf1116c0d1db3aa21bf52ac = ~I171149dcaab2c0f0e2a10547ad95084d+ 1;
assign I566c72342c69969892480fae41232c37 = ~I23b60ca4da2df0ec40c1df62d058deef+ 1;
assign Ia0f7deea6b1ce1050dcf97fa99de9178 = ~I7978d2d800b4438d0644ae3df6bcac9c+ 1;
assign I992b9876530d53c1b62d98511bf41942 = ~Ibc4eddc0f1768e9ec7e38e951a28ec42+ 1;
assign Ib8861f627f6273c0a031bf43e7812a5d = ~I1c97fd1d21a31af8b5498a79b1a3e7b6+ 1;
assign Ieb5bac4ef0f5e4e0b826cdc43ae71471 = ~Ie4f063eeaf7ee3f033e2a01ffaca623e+ 1;
assign I3cd0883d9f0ba7475f474f1e318ef023 = ~Ibb3d57d510cad00064a331f61f6400a2+ 1;
assign I5f8a41ab83a9257e534973e981e28e9b = ~I9485ae915474a31562ce358666d66245+ 1;
assign I0e420136675d5f0d1aa027d589ee8741 = ~Ia54b6f7044a831020e49f1bf48bc063a+ 1;
assign I4aab6ff52e3fba90bb7417cb50766125 = ~Ie71c7babb5d17378d40444b6bbd4e7a6+ 1;
assign I1ba7f209cb735471073e8051026a148c = ~Ia0977b79857bdbf058535c30e338c38a+ 1;
assign I711c5cf9fd8c5161bac36060b3443503 = ~I600ea1371a2be66430ac9534583b512b+ 1;
assign Ie3591b22e0e127f04658da68d4846be9 = ~Ife5b9afdbb30c122b84d5378f9cb366d+ 1;
assign I409129c0bf5d361e9916b6dc98e69a7d = ~I27556d599dd1a27ee8f49e819ccbf29a+ 1;
assign Ie4f4faa470f572da2081b63b6df6e392 = ~Icce595233ce089eafcca3eae5e71e5f8+ 1;
assign I5011dfbbb0eccfebcff255e4a2c5e64c = ~Icc3cadf40c09be1a8c2847caf0e3e63c+ 1;
assign Ie32ca6b91d1c55883be8f63acca78764 = ~Ib43886d923b8c683004713ff25b2f90d+ 1;
assign I6c7965d39dc839a9df56e628c77a5457 = ~I132d9671c582876568c0f7f5335f5227+ 1;
assign Ieac9cea5f36bd82f87105b530e8fb614 = ~I0859c80b42a8c60dade8f05d58ee3701+ 1;
assign I79657595561eac53237215fb4110f09d = ~Ib3690ec149adde94343d3e617931a287+ 1;
assign I9b46463a6c54c3668e76190d942b7b38 = ~I41f2bf9ff00f983ad1298c8c83b041cb+ 1;
assign I3ff883ad434cd5153b67186b6b21418d = ~Ib5414585cd6976cfce42e42190cc08d7+ 1;
assign I92abaae6fb89206885616877cca1e25a = ~I1ca59325ff30db83df5bf0a2cd9706b6+ 1;
assign I33668b0ef7defef974b7a4c0f87689c0 = ~Ie2f5b03f3b136e651b8aba92a30d298a+ 1;
assign I338daeacf82ad288b14c6b5bd4099870 = ~I312ce79a8dd2ce3d37c930d42640509b+ 1;
assign Ibe085a39ecb07a8dca62002afa38df93 = ~I467d5e2554ef25873e0b44e947ee0011+ 1;
assign I1f88dddf05f255942e2749891a7733da = ~Ice73b514709469fd21cd254bf4ceadd9+ 1;
assign If1d0be4e9b995ec98c346e8392b9518a = ~I45ba06a6d6f00c174b1439a6f226a085+ 1;
assign I56a4443759b3d786bc9a34a0dc32abf0 = ~Ic8a272f82736fd599fb3250e970edf9b+ 1;
assign Ic826d371f2cfc503f5d9e43dc17481e1 = ~I5b9710b16effc8bf0695517c6e651836+ 1;
assign I5502f383dff392ef1be4cbbf9dbc3c2f = ~I038b42a83025f5eaebf45799d1ebe7b0+ 1;
assign I96e6f1dc0cd451da6ac9170d5f83976d = ~I73ddd7cf9272ceab5a663e2244e72d7e+ 1;
assign I10cd840a369d3e25556a41beede2be27 = ~I16507fab8f9076bfeb419896fa7cdc1d+ 1;
assign Id85c2285fcc45211f0fa6963b74a663a = ~I3dd1f28cf199299aba54e47a429c9b11+ 1;
assign Ie0bdfac78159144aa65090028931a3bf = ~I49d9203dc6f8c17f17383e8f7e01f005+ 1;
assign I28fa30cd1f3b476fa6a354863108cbcf = ~Ibeec86c75d950ee00dd63a2930f08a24+ 1;
assign I7a927f4f266cc5253ec30f5c127bb17a = ~I47b2438c3680b2d816168df37d7c491c+ 1;
assign I7571c7c306861230de71a75fca79c5dc = ~I5983bf2c6c90b872ee6cf58b5e520311+ 1;
assign Ic79811a48840357d0b6303e7b19413dc = ~I6745cacecb7ee86cf3c7ad7eeee6048f+ 1;
assign I0f29300446f020dd23cf847d3e3d3530 = ~Ib9672d20643d856ff31905ab14c0ac87+ 1;
assign I802bd5b13c183c37e842f7e9278f35a9 = ~Ib9dfea1f34a120eda30d5bd919365a6a+ 1;
assign I0297905b35f06697625420b7fc2434f7 = ~Ia7bf82c9e5ca4467b5e50beeaeb975e9+ 1;
assign I8487a819dcb61016798cde56f9662fcf = ~I327c9acb8934729b4ea5486787afa2e8+ 1;
assign Ia2904a5d5db43a209bd4b358ace68c6a = ~Ieddef08050c38d07e5d38f5bb7b099c0+ 1;
assign Ia8b29ca047a643f47bd3a0ffb50bf8cb = ~I39f9e8430db114991bfb27cc46ef3e39+ 1;
assign Ic45d0537b94bc30713c0a0ee07b1ec40 = ~I56aa548618a4a15e9a35e04f5eeb823f+ 1;
assign I337231f0dc7eb85f7d950262e0adb724 = ~I1908897b529ca04df7e7da395be4a8ce+ 1;
assign I530cf1f747d1df44b913f49eee90c079 = ~Ib2bbd59cd6098608ed53ac556036534f+ 1;
assign Ief52461e4a5ddb128be5e439edf34862 = ~If004552b2047ab1cf23bb50375460b01+ 1;
assign I46d86bfa6de26f3cfef9d802549ef2ad = ~If97092e1e2147de199c94a23831cf6b9+ 1;
assign If6a3bd6f002d91e0773c4ab9caaaa01e = ~Ibf74a4dfaab7f7f538d2b5fac7394b63+ 1;
assign Ib33e1c6d57e5e6fc465dc9c9a7cf29fa = ~I991a7a7d562eb0a8b4b8d8f008ef2225+ 1;
assign Id92a319da408be46970faf524513fdd8 = ~I64c3d7be41abaa17d6992f9af8e72789+ 1;
assign Iae182ffae6cea89363f0ccc8b5679561 = ~Icb91e63ebabc7a75a54eb7c731df4fa0+ 1;
assign Idfe6aecb694385ce8c3c1544a4992a20 = ~I673d1d0d0daab99bd940c46cc14ef55a+ 1;
assign Idfbc5726963cfa31bb4324143ffd08c7 = ~I62cadbd70b07a6a7a2974c7c392696b3+ 1;
assign I205d5fdeae55fae7be2f06f11c949244 = ~Icd8257d7f53d93db989eb56eaeb7e593+ 1;
assign Ie667e1755ae1561a2eefae9b63845dec = ~I05931ceae6eff26e5a66a44a54d628ae+ 1;
assign If7348fdbe0400aab92e8fd6a7cf6c267 = ~I306fec0aa68a0396053a6e0fa1cda38f+ 1;
assign I143b91852fddcdcc30bf1041332c4ed7 = ~Idee8c8144207d676d1f2f9064bbdff45+ 1;
assign Iee5e74945ba15220f0f707c9c1927ba1 = ~I5855124d566af739caa6511f8598f2c5+ 1;
assign I4d1c47569b0bc8c651c897ac8e88bd1f = ~I50729db4a8e04f18979707df14cb2419+ 1;
assign Ib9d6c5be487a434fbafcda25ca9351dc = ~Ia3cb3ea64576a3e7332e1fb55953aa3e+ 1;
assign Ib0d033ba28e8c606ed92207049c76884 = ~I3cb1f233951d49f985b0deac6e052bfd+ 1;
assign I300d9f403e33d860ff5dde9f91bae11b = ~I7015def91103398e54f446ce3e43af01+ 1;
assign Iebfe0fa45e4b34e142e82ddaa15243cf = ~I04874bd1bf257f205b5189c8c20e5a12+ 1;
assign Ieb778442bc855e93e11c9b13f1a7ae06 = ~I937e3a8ede2305ea7c1750283224a870+ 1;
assign I57a393cc9cc9e1abc7962aa2cc840a7c = ~Ia7206430a739a11af4d860096eedd6c3+ 1;
assign I0ffb8b65525af38861280645ac310e3d = ~Ibf4c2c00f8e012e9498361bfd3c5b06e+ 1;
assign I30fb41a57460a0b1f21065b4b97ddd42 = ~I899e5f03cd1d52d11f898959559aaeea+ 1;
assign Ie8298c5c8ff538a3e37af46798f6d753 = ~I59c80c7ec26f43308b1a646c47160568+ 1;
assign Ie7dc322fee8ca0b6b9659e5183e0d6d6 = ~I8a954a331d36266465a0813d2e8b319b+ 1;
assign I91bbec0523f77fc52a88ebcc49267e9c = ~Ib49e53ca8efd9564ee9572eb3089bb51+ 1;
assign I38ae79956762380fadc94f8126dc1c90 = ~Icbde2c6230e9cc67ef12031e38bb344f+ 1;
assign Id55a1ab9d158ea509e5f57286a3d1b67 = ~I2e22e867f6f84a7807b82f64a147022e+ 1;
assign Ice615e7e18356ae4c3f615dd997be943 = ~Id9704e1d8096cd28577c5c357d30b7a4+ 1;
assign I57b40c72004f2c3072cbdefbeef72b7c = ~I4b8554cab486a4fc1e14884a6495016e+ 1;
assign Ie38351e19bdc4f2ce9caf75fc3937dd4 = ~Iaa235d085a5916a3b0814c3ed2a9026f+ 1;
assign Ibba6269b560db9d4913e1e515ed8270d = ~I5d86ce0b58c0b281d747116a9069ef33+ 1;
assign Ie392719059587a201c0148138ba2a2d4 = ~Id20394136fb036435bb4680aac64581f+ 1;
assign I4852d6bacfd82fef6fab4502d61e9a37 = ~I8a16afac6e470ca69634d7fe9656387a+ 1;
assign I9200526d94c38e638370e9a2d7fed75c = ~Ic4e7f690bc050f1d1f84eae7ca193e1c+ 1;
assign I15b8aa7d973edcf3b2365040f5570d82 = ~Ia60421aa427236540b4d0d08d52ff507+ 1;
assign Ic3f8e77259ee3eb5be80e11b607818bd = ~Icace650ee3865bd7bbddd2d9435c5561+ 1;
assign Iabf228f57ac154c417389f6711af1950 = ~I7d27d070b96b7810f667e1d1845342d3+ 1;
assign If37de611ce4fa330c4fc9dcb87d4d95c = ~Ida7ec09c913caa0e78a2c4cbaae517c8+ 1;
assign If3c44eb85217da3b6bddb5aed97a9bb7 = ~Ic5eba898858be1f768841ead792d6d86+ 1;
assign I8c36318c45dabe6bf540381373f09fe5 = ~I72197797a307c611fa8952533e63d7bf+ 1;


Ic3da32f100a43f826b89a492544e7812 I8bed3fb56eecc27b4fcbb5cfc2f52746 (
.flogtanh_sel( Ic93835a022c46b7aa00a465c407d7da2[flogtanh_SEL-1:0]),
.flogtanh( Ia67805b59c3011bc4fc5cb1d2996f90d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(Iac11baea9832d6493626d2fe40fd385f),
.rstn(rstn),
.clk(clk)
);

assign I5f68368511b59d2e365cc91b806b334e = (Ic93835a022c46b7aa00a465c407d7da2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia67805b59c3011bc4fc5cb1d2996f90d;


Ic3da32f100a43f826b89a492544e7812 Ie7b83a9c62be138cc7fd9250dffea62a (
.flogtanh_sel( I2e30088bf29cedd7debc15b1e6ec4ada[flogtanh_SEL-1:0]),
.flogtanh( I61fb47b07547e09c746b1fb5d7c8710d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I71e4d98dca37256fcc84248a26d703e2 = (I2e30088bf29cedd7debc15b1e6ec4ada[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I61fb47b07547e09c746b1fb5d7c8710d;


Ic3da32f100a43f826b89a492544e7812 If7365105b4359266502e1931893366fa (
.flogtanh_sel( I38f512bfb84094d1e92a10a345d5505f[flogtanh_SEL-1:0]),
.flogtanh( Ib2220549c84e87683ccf85798b2bb22f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib8380902ac4082f834744ddef6d0cc6a = (I38f512bfb84094d1e92a10a345d5505f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib2220549c84e87683ccf85798b2bb22f;


Ic3da32f100a43f826b89a492544e7812 Ic00f96f8dc955b5e4979a2dc3a2a44b1 (
.flogtanh_sel( I1e878f00f056f637625cb013a93325a8[flogtanh_SEL-1:0]),
.flogtanh( I12f063ad18938c2ca008e1165f9119e9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9570f8498d95bee230bb3c5e720bb857 = (I1e878f00f056f637625cb013a93325a8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I12f063ad18938c2ca008e1165f9119e9;


Ic3da32f100a43f826b89a492544e7812 I69480aafea8257c5437ac4373ad1c1e6 (
.flogtanh_sel( I25db27464b31fee41ccd7a3cfe4d403e[flogtanh_SEL-1:0]),
.flogtanh( Iae6b4023f9f2641ca00636181f4fb028),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I55c425102db0a6838012a165c0597680 = (I25db27464b31fee41ccd7a3cfe4d403e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iae6b4023f9f2641ca00636181f4fb028;


Ic3da32f100a43f826b89a492544e7812 I271d4e9c0c6ca43854eeb7b986431d7c (
.flogtanh_sel( I19417a224c5cdf1211e9790aa29c4c5c[flogtanh_SEL-1:0]),
.flogtanh( Id11b7d1aeb413fd4920ef0e0097fc6c4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic970a88c435a85d21ed71c6060b8a8e4 = (I19417a224c5cdf1211e9790aa29c4c5c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id11b7d1aeb413fd4920ef0e0097fc6c4;


Ic3da32f100a43f826b89a492544e7812 Ibfd3c16dea8a2c68944ec5e93a234c1c (
.flogtanh_sel( I16dcafa854ea9c67d8a080feb2ba9166[flogtanh_SEL-1:0]),
.flogtanh( I3af03d3e0bb7e0e73e034dceda70ff3a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iec8dc328edd6cbaa2d697e05ed222746 = (I16dcafa854ea9c67d8a080feb2ba9166[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3af03d3e0bb7e0e73e034dceda70ff3a;


Ic3da32f100a43f826b89a492544e7812 Ie5a7b0dafa40187048c7e75670ac9cba (
.flogtanh_sel( I7f63338eee2663fbe61fffd248433310[flogtanh_SEL-1:0]),
.flogtanh( Iba30a494dc1b66bd2862f82c16017a99),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I16d2084ccfb102c3bafc701872f5ef2d = (I7f63338eee2663fbe61fffd248433310[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iba30a494dc1b66bd2862f82c16017a99;


Ic3da32f100a43f826b89a492544e7812 I535e8c8f08c8546ab637017ebbfb55fc (
.flogtanh_sel( Icb1e3c56c8729c32d43c69710e345db2[flogtanh_SEL-1:0]),
.flogtanh( Iefa075dc743d616eca65f76d2c03371c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id680a9affed622577164b3a8380494f5 = (Icb1e3c56c8729c32d43c69710e345db2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iefa075dc743d616eca65f76d2c03371c;


Ic3da32f100a43f826b89a492544e7812 I899ada2d26f95030e673433fb46d8a92 (
.flogtanh_sel( I6ece8e3c1e89613879336936f77d732f[flogtanh_SEL-1:0]),
.flogtanh( Icc7a632da404a9cda7b8247706391f85),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifcd68be4bea38622d2d57d3a4e6fc5bb = (I6ece8e3c1e89613879336936f77d732f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icc7a632da404a9cda7b8247706391f85;


Ic3da32f100a43f826b89a492544e7812 I00cf63ffb5c51cef81a8824d96eef6a6 (
.flogtanh_sel( I72a646ae7e32a16af0f5930a6e95b36a[flogtanh_SEL-1:0]),
.flogtanh( I708c5d8d6d8f7f16c2f348c3b97b906d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I16deb9107193a3536979e4b5e5654b9c = (I72a646ae7e32a16af0f5930a6e95b36a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I708c5d8d6d8f7f16c2f348c3b97b906d;


Ic3da32f100a43f826b89a492544e7812 I03b5eacbef8fd3e4d61df6c09d373ee6 (
.flogtanh_sel( I7e72d119dd93a6ab05a23fde0a865866[flogtanh_SEL-1:0]),
.flogtanh( I51ba1e25e01c39a77559089626bafa09),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I28cac65a4db3f708cc90a1b023bfe894 = (I7e72d119dd93a6ab05a23fde0a865866[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I51ba1e25e01c39a77559089626bafa09;


Ic3da32f100a43f826b89a492544e7812 I25a3636d0a391ac3a95169e451e49935 (
.flogtanh_sel( Ied4fdf5805039cd2fcd042fd13755fdc[flogtanh_SEL-1:0]),
.flogtanh( I2217e483aaf5124d9beb9baf5037326b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie763738b7faf253837e1c45de255cb5e = (Ied4fdf5805039cd2fcd042fd13755fdc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2217e483aaf5124d9beb9baf5037326b;


Ic3da32f100a43f826b89a492544e7812 Ib8648fb43b0b9d0a49a204accd49e601 (
.flogtanh_sel( Id44c2293b765cff450dd1d747c47c1f3[flogtanh_SEL-1:0]),
.flogtanh( Ib47f8220e7a319e690649f9d6cc9f0cc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icfef12499b53cd84f0aae067f30c17d0 = (Id44c2293b765cff450dd1d747c47c1f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib47f8220e7a319e690649f9d6cc9f0cc;


Ic3da32f100a43f826b89a492544e7812 I82d8ce125217b65528b7ad8a1005a894 (
.flogtanh_sel( I8f4ed02f7aeb823b745040f7f3f43ac7[flogtanh_SEL-1:0]),
.flogtanh( Iffc502b536d88d080c59eb3aedd55bd1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0982b8d7f99aceb8871c9c10448f54c5 = (I8f4ed02f7aeb823b745040f7f3f43ac7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iffc502b536d88d080c59eb3aedd55bd1;


Ic3da32f100a43f826b89a492544e7812 Iacfee3ae0e57744f4d474f386dc383c3 (
.flogtanh_sel( I6488b9b8f405d7d81a4874fab2678102[flogtanh_SEL-1:0]),
.flogtanh( Iaa823b6b13acb376f979dd52683a2231),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6c661048307c23c699d4b3636564de0f = (I6488b9b8f405d7d81a4874fab2678102[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaa823b6b13acb376f979dd52683a2231;


Ic3da32f100a43f826b89a492544e7812 I696328955cba7f8540e195046ce2341c (
.flogtanh_sel( Ifff612d16828ec907a348479e19ddf31[flogtanh_SEL-1:0]),
.flogtanh( Ic5f3f371b1ebfe733404b4165fe746dc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I786dfcaa131b99c254aaff15bd2c2b6d = (Ifff612d16828ec907a348479e19ddf31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic5f3f371b1ebfe733404b4165fe746dc;


Ic3da32f100a43f826b89a492544e7812 I977277221a170e898622260e22727cf3 (
.flogtanh_sel( I268262076f22bc6b1507bc8f91b98a0a[flogtanh_SEL-1:0]),
.flogtanh( I021d991730d154218106f00e74bf9d4c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2b49d74cb130542f2ca99534e2c513b1 = (I268262076f22bc6b1507bc8f91b98a0a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I021d991730d154218106f00e74bf9d4c;


Ic3da32f100a43f826b89a492544e7812 Ib9ff92e7058da35313862d7081d58dd8 (
.flogtanh_sel( If1f732841adb7c0cad1ba37c0f5fd517[flogtanh_SEL-1:0]),
.flogtanh( I688e5b6520508178afdf85bb2194186d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0f6cb7a5a31d6f2f6178632c0c898bc6 = (If1f732841adb7c0cad1ba37c0f5fd517[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I688e5b6520508178afdf85bb2194186d;


Ic3da32f100a43f826b89a492544e7812 I9e1dccf22f01d1ae330a488c70fc0a4d (
.flogtanh_sel( I0df8a24f31c027756d248c3bd1b9bf7b[flogtanh_SEL-1:0]),
.flogtanh( I658630f3cf0e86ea86c5fb78b025b0a5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I03bea609a189246a2375b355df47cf81 = (I0df8a24f31c027756d248c3bd1b9bf7b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I658630f3cf0e86ea86c5fb78b025b0a5;


Ic3da32f100a43f826b89a492544e7812 Id26df530f2fe0c907848c8f6bb3e8e71 (
.flogtanh_sel( I8ef901e733b12e76412eb36684e2b575[flogtanh_SEL-1:0]),
.flogtanh( I8b17f8bae259d829b52aba173bf10b4f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If56555b7cf539750706cf678030ccdb2 = (I8ef901e733b12e76412eb36684e2b575[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8b17f8bae259d829b52aba173bf10b4f;


Ic3da32f100a43f826b89a492544e7812 I3a008e7478eb890f467c2447ced05e42 (
.flogtanh_sel( Ia48916a02f68b1b8f5fc7fece04677bb[flogtanh_SEL-1:0]),
.flogtanh( I944da8181119550916eaf431c7b04c50),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I94e89b3a841f9760e3967c97e86d7160 = (Ia48916a02f68b1b8f5fc7fece04677bb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I944da8181119550916eaf431c7b04c50;


Ic3da32f100a43f826b89a492544e7812 I741118d8af6cfed44fbf85a975ed9088 (
.flogtanh_sel( Ia37409944d9fdd3b16e7007e13d82a79[flogtanh_SEL-1:0]),
.flogtanh( I3aa615fa11ad382432ca658ec233f094),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8cab6f6faf0758f26d1a8851fae43896 = (Ia37409944d9fdd3b16e7007e13d82a79[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3aa615fa11ad382432ca658ec233f094;


Ic3da32f100a43f826b89a492544e7812 I423a5b0b0ebc1a90d8f436ca8ed2440e (
.flogtanh_sel( Idd65f149afe9d5f63ddaf34b82b11e95[flogtanh_SEL-1:0]),
.flogtanh( Ib7c4f77c160ec436e93ca9de75b9fe42),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6ecf7249e6151477fe74a79d0b126b21 = (Idd65f149afe9d5f63ddaf34b82b11e95[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib7c4f77c160ec436e93ca9de75b9fe42;


Ic3da32f100a43f826b89a492544e7812 I018f2c494128a900c65ee1099848b918 (
.flogtanh_sel( If2886d560854faed32ebd8e33d868973[flogtanh_SEL-1:0]),
.flogtanh( Ic1e06942b276ee0933dc8b85dec58756),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3753b2c4ba8f1bee70def390a96586b0 = (If2886d560854faed32ebd8e33d868973[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic1e06942b276ee0933dc8b85dec58756;


Ic3da32f100a43f826b89a492544e7812 I564054cbca01fcf8c4afb77505e627e1 (
.flogtanh_sel( I77778118bb3ea900c080754ff4c49c26[flogtanh_SEL-1:0]),
.flogtanh( Idd96d8b4e7be386203ec3ed3a81391d9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9b919f3d4ee3f33506b87bcdaf2d43a3 = (I77778118bb3ea900c080754ff4c49c26[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idd96d8b4e7be386203ec3ed3a81391d9;


Ic3da32f100a43f826b89a492544e7812 I1e03de209c3c3bdc860d89cb5ab87ecf (
.flogtanh_sel( I7292ed752d8741594d757730950feea4[flogtanh_SEL-1:0]),
.flogtanh( I7df43eec4d78baa1e0680be2715c4495),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib3be128b6704cc04c61e0fc9814dcf20 = (I7292ed752d8741594d757730950feea4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7df43eec4d78baa1e0680be2715c4495;


Ic3da32f100a43f826b89a492544e7812 I7d56e9ad387ba285bc760f691fea84ab (
.flogtanh_sel( I68cfd7868e061793ee8a41e69e80219b[flogtanh_SEL-1:0]),
.flogtanh( Ief08536c38479e6bc7fe786cfaf9a10f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If365a3c3ef86dca7c7315b91298c2db8 = (I68cfd7868e061793ee8a41e69e80219b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ief08536c38479e6bc7fe786cfaf9a10f;


Ic3da32f100a43f826b89a492544e7812 I31e0860f6ffc1be7190f10f841d1c858 (
.flogtanh_sel( I667ead814b303fca64ef047bb8246b19[flogtanh_SEL-1:0]),
.flogtanh( I6ef440b2077563ebbe50dde593c3875a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I83560e8d0f8cd37815cca6336fb2208d = (I667ead814b303fca64ef047bb8246b19[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6ef440b2077563ebbe50dde593c3875a;


Ic3da32f100a43f826b89a492544e7812 I6c7a7abb57b8c9fd9cb6a7ea48563160 (
.flogtanh_sel( I4f25c7edb12e868cb5532e42b4ba5133[flogtanh_SEL-1:0]),
.flogtanh( I20cfad172f0a614687d72d2337ef1003),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I099441ae3d3dffe49b18bc578af54dc7 = (I4f25c7edb12e868cb5532e42b4ba5133[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I20cfad172f0a614687d72d2337ef1003;


Ic3da32f100a43f826b89a492544e7812 Ic356506f770623f8e3505df62d6ca688 (
.flogtanh_sel( I5aed2d82717f359bb5ac5a0ab91b7beb[flogtanh_SEL-1:0]),
.flogtanh( Icc6a92285959b25d53b452aed0718c8e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I58f89947eead94b5054a0fea3520ae33 = (I5aed2d82717f359bb5ac5a0ab91b7beb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icc6a92285959b25d53b452aed0718c8e;


Ic3da32f100a43f826b89a492544e7812 I772300d29a37ded7289001e5b6fd75b2 (
.flogtanh_sel( I92835fd54631deaefa7b214e2c4b9bff[flogtanh_SEL-1:0]),
.flogtanh( I132c12f1eafbe34bca7b070354bd5f43),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibf565bf1803ed43120fa54b80f6f1f29 = (I92835fd54631deaefa7b214e2c4b9bff[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I132c12f1eafbe34bca7b070354bd5f43;


Ic3da32f100a43f826b89a492544e7812 I7241058865140c737c113ee9a2a3c426 (
.flogtanh_sel( I67e067da565635fcff166e3a7d0c446b[flogtanh_SEL-1:0]),
.flogtanh( I0f327225758bc82a67a65b8714949a91),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I619957528c630e7f64924a25127c93fb = (I67e067da565635fcff166e3a7d0c446b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0f327225758bc82a67a65b8714949a91;


Ic3da32f100a43f826b89a492544e7812 Ic56e9245dfa44e3f60a947364bfa3217 (
.flogtanh_sel( Ifdb0f307b1b9458c0487a1574ccc094b[flogtanh_SEL-1:0]),
.flogtanh( Ia90d4bc44d3687e912b59e4b6ca02718),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If3cc31fd16469339470702045fc6d0da = (Ifdb0f307b1b9458c0487a1574ccc094b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia90d4bc44d3687e912b59e4b6ca02718;


Ic3da32f100a43f826b89a492544e7812 I4b06d92359835a1ee9d1d0f7fc92a387 (
.flogtanh_sel( I5c6b7d143e42fd3b8bcdb7d7ed4da2c2[flogtanh_SEL-1:0]),
.flogtanh( I21c1757545cc2732445c7f978f7247c4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I338ccc17dc6158aec0129c8b0c02c429 = (I5c6b7d143e42fd3b8bcdb7d7ed4da2c2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I21c1757545cc2732445c7f978f7247c4;


Ic3da32f100a43f826b89a492544e7812 I4c55988c9baabcfa9d505ed4193d4895 (
.flogtanh_sel( Ie679a21d0136a08cc5e6526e9f8d1843[flogtanh_SEL-1:0]),
.flogtanh( I096fb1aff9431ed667e5d85a6f3726a4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I83d71a89f35eb73265ee3e54184e1277 = (Ie679a21d0136a08cc5e6526e9f8d1843[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I096fb1aff9431ed667e5d85a6f3726a4;


Ic3da32f100a43f826b89a492544e7812 Iaa2713a943196d86c7b34fa93e5977fb (
.flogtanh_sel( I611942a72a5e12f6afaea6bde6699ef6[flogtanh_SEL-1:0]),
.flogtanh( Ia69d80cc1f2957ccd79cbd466dea987e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7362f08ed4e4ae309dfbfda112c56ad6 = (I611942a72a5e12f6afaea6bde6699ef6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia69d80cc1f2957ccd79cbd466dea987e;


Ic3da32f100a43f826b89a492544e7812 I6078e0efbdf6d793f388ebb21ffc369b (
.flogtanh_sel( Ica9883c97f823a4491cbee5b45c43590[flogtanh_SEL-1:0]),
.flogtanh( I2243822bb5cdbca7f2ea942c7b720da8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8be4be8471625db0749e6385f87d2dcc = (Ica9883c97f823a4491cbee5b45c43590[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2243822bb5cdbca7f2ea942c7b720da8;


Ic3da32f100a43f826b89a492544e7812 I67c595d9f8f2b459cb145d8128790843 (
.flogtanh_sel( I8e6addfc61f5bfb7af74fc2993639565[flogtanh_SEL-1:0]),
.flogtanh( Ia77953e90a0cb40984d138c2c209db01),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3d6a685a1913bd8be01fddbce1edec2e = (I8e6addfc61f5bfb7af74fc2993639565[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia77953e90a0cb40984d138c2c209db01;


Ic3da32f100a43f826b89a492544e7812 I80ab0c2ebe798763b2ac22dcb148b76c (
.flogtanh_sel( I9d53619f10e2a426f7297bbf7c81158a[flogtanh_SEL-1:0]),
.flogtanh( Id0b03e6dafabbe570f2626f51c9b7121),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifd77e040c5f82790b1d5636a42fca602 = (I9d53619f10e2a426f7297bbf7c81158a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id0b03e6dafabbe570f2626f51c9b7121;


Ic3da32f100a43f826b89a492544e7812 I96b6904ec785c131b076aafe2d86597c (
.flogtanh_sel( I8a055c27778913287ad951183fa0d4d6[flogtanh_SEL-1:0]),
.flogtanh( I5bfac7858439b218179c95c8d8669f17),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifbe479e5cab3cba43444bec1e12e72a0 = (I8a055c27778913287ad951183fa0d4d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5bfac7858439b218179c95c8d8669f17;


Ic3da32f100a43f826b89a492544e7812 I04e1872d4b35b4c3c071d7d981f794a9 (
.flogtanh_sel( I8f6ae5c80bb2f50084b5f5ee5ab0ffc3[flogtanh_SEL-1:0]),
.flogtanh( I52497c500164c2417f928196ddcdbf84),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia784f35a5a46837b69eb048dabf84052 = (I8f6ae5c80bb2f50084b5f5ee5ab0ffc3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I52497c500164c2417f928196ddcdbf84;


Ic3da32f100a43f826b89a492544e7812 Iaad65d61da236eeebf30744c7bda6126 (
.flogtanh_sel( I3db8b3a342e8e2f13a448246aa001c2f[flogtanh_SEL-1:0]),
.flogtanh( Ib499dd504da7e433bc1caa258d7e7101),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8d0f440df332ea96e2d56eec490fbd51 = (I3db8b3a342e8e2f13a448246aa001c2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib499dd504da7e433bc1caa258d7e7101;


Ic3da32f100a43f826b89a492544e7812 I23591a2c75507627957aeba252565b19 (
.flogtanh_sel( Ibbee0996ea0f5e16b1f711345be7f2ae[flogtanh_SEL-1:0]),
.flogtanh( I7af88e2be096e488d7269479f935d185),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8d431a0524241fa54cf6dd1e79de4c74 = (Ibbee0996ea0f5e16b1f711345be7f2ae[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7af88e2be096e488d7269479f935d185;


Ic3da32f100a43f826b89a492544e7812 I22d8cee416a0f827720e02957b13c074 (
.flogtanh_sel( Idb777f1eb4c3cbba103b9b43f948ccf9[flogtanh_SEL-1:0]),
.flogtanh( Ief51cc849e0034a9a6b3ff061064ad64),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If49f97cc0c42b23ce393b534015559a0 = (Idb777f1eb4c3cbba103b9b43f948ccf9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ief51cc849e0034a9a6b3ff061064ad64;


Ic3da32f100a43f826b89a492544e7812 I15aaa4edb37eb15195676a84ca44dbde (
.flogtanh_sel( Id5e46b1f8844c7587f99d22170581a24[flogtanh_SEL-1:0]),
.flogtanh( Ic5f096a42ae6fec933dcaf85faeeda49),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie932a22a7f1fa37087cbc9e8d73efef4 = (Id5e46b1f8844c7587f99d22170581a24[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic5f096a42ae6fec933dcaf85faeeda49;


Ic3da32f100a43f826b89a492544e7812 I93d5604164d223b8b1a5f196431f4da4 (
.flogtanh_sel( I67aadabd3cf49456cace7392a1e7a35a[flogtanh_SEL-1:0]),
.flogtanh( Ic9c0a2ce51d641ba7896c2c6911d0f96),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2956687a5fc2fba7149889624ef85647 = (I67aadabd3cf49456cace7392a1e7a35a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic9c0a2ce51d641ba7896c2c6911d0f96;


Ic3da32f100a43f826b89a492544e7812 I8832a7ffac105d2d57732b166dc51f2a (
.flogtanh_sel( Id5635595d6b7b6dd7e6d510a27ad6702[flogtanh_SEL-1:0]),
.flogtanh( Ia96b3ea2e8395671b3ac674f5a956771),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iebf28886bd39c2540c90e808a9c20d3d = (Id5635595d6b7b6dd7e6d510a27ad6702[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia96b3ea2e8395671b3ac674f5a956771;


Ic3da32f100a43f826b89a492544e7812 Id1e5aff4b204e2b5364dbb9e49840461 (
.flogtanh_sel( Ice783314a4868f0bba8bc3c5e3b65ae4[flogtanh_SEL-1:0]),
.flogtanh( Ib81d241e073c97c8c8d1d0abd9a9a64f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8d4f3e64c8e3b0710a4a6b30d27c8be8 = (Ice783314a4868f0bba8bc3c5e3b65ae4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib81d241e073c97c8c8d1d0abd9a9a64f;


Ic3da32f100a43f826b89a492544e7812 Icca1b593c5c92beb6812d268808f9d22 (
.flogtanh_sel( Ib2d9b7f58cf571b904be02e6073f9b94[flogtanh_SEL-1:0]),
.flogtanh( I0fc5e49719d7132c7724ee0d406ff93e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I16e3f3a6802fd206654bb622fa1393fe = (Ib2d9b7f58cf571b904be02e6073f9b94[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0fc5e49719d7132c7724ee0d406ff93e;


Ic3da32f100a43f826b89a492544e7812 Id3d956051c977537249d54b05abb3127 (
.flogtanh_sel( I61b6effae91ae4bdcce4550eb5cf0796[flogtanh_SEL-1:0]),
.flogtanh( I4479a0c26d4fa67dee328ecae12d14a4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4b5713aee09999592256c407d4b8a95a = (I61b6effae91ae4bdcce4550eb5cf0796[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4479a0c26d4fa67dee328ecae12d14a4;


Ic3da32f100a43f826b89a492544e7812 Iefb4b4f6c5d35224af9dda1b2bcb5e93 (
.flogtanh_sel( If5cf6e81b0e3b77f6a45f2555201acc2[flogtanh_SEL-1:0]),
.flogtanh( If5693e079544d04478ec3da9a0ba28d7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieb1dbb98d5e5bda5b9ce803857f2ca26 = (If5cf6e81b0e3b77f6a45f2555201acc2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If5693e079544d04478ec3da9a0ba28d7;


Ic3da32f100a43f826b89a492544e7812 Ief314496bb908b7eea2c32a68480b093 (
.flogtanh_sel( I62fae5bf51588f28c3521715b834909d[flogtanh_SEL-1:0]),
.flogtanh( I701a0ec899c88feef97aeb45fe19e639),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ife1c8d014675240a94f1133a78703ed5 = (I62fae5bf51588f28c3521715b834909d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I701a0ec899c88feef97aeb45fe19e639;


Ic3da32f100a43f826b89a492544e7812 I4d547789af8b24398e22c22015401a3a (
.flogtanh_sel( If5cbdab78a4cf86b6285a400d0e0ac90[flogtanh_SEL-1:0]),
.flogtanh( I6e9d61b111a45e4ea92ff12d33801755),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I94d9412a7b43fa0bd4b9a6d32d313fc7 = (If5cbdab78a4cf86b6285a400d0e0ac90[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6e9d61b111a45e4ea92ff12d33801755;


Ic3da32f100a43f826b89a492544e7812 Iead32f99096ab34ce26cd8a507537a26 (
.flogtanh_sel( I6e481cc49441c08bcd9fdcabbe90a000[flogtanh_SEL-1:0]),
.flogtanh( Ief65b0dab6ce1c2fc23cd297a21ac8de),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If13e359e530823319046ce20027445dd = (I6e481cc49441c08bcd9fdcabbe90a000[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ief65b0dab6ce1c2fc23cd297a21ac8de;


Ic3da32f100a43f826b89a492544e7812 Ib6ec46aa056c63d9255beb163a4ddda2 (
.flogtanh_sel( I3aa663be3dd604564ef68b9a2b9d7319[flogtanh_SEL-1:0]),
.flogtanh( Ibb843c4198a06c8e46bc954663c52a28),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I221777352b48c4e228c6637410113854 = (I3aa663be3dd604564ef68b9a2b9d7319[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibb843c4198a06c8e46bc954663c52a28;


Ic3da32f100a43f826b89a492544e7812 I51c25a9310e7baccb7abf1ae59f6cd5c (
.flogtanh_sel( I8031632ee8700c63c207e2d6a6bdb630[flogtanh_SEL-1:0]),
.flogtanh( I0c043ef5daa388e93fb3cf6465c217b5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1ee46fec2b82cf8e5142f8e2ac5d9d8a = (I8031632ee8700c63c207e2d6a6bdb630[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0c043ef5daa388e93fb3cf6465c217b5;


Ic3da32f100a43f826b89a492544e7812 I92420c9da0b36e4ce41b2b81c61e7b39 (
.flogtanh_sel( If9be2701858da0bdffbf2dff7bcfd7e1[flogtanh_SEL-1:0]),
.flogtanh( Ife3f07ad3ad5228f10da7020a01e7069),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie45aaf966aa0a94803050b5f43d69e6c = (If9be2701858da0bdffbf2dff7bcfd7e1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ife3f07ad3ad5228f10da7020a01e7069;


Ic3da32f100a43f826b89a492544e7812 Icbc2d07d815f28f31874a73ff31ef1d8 (
.flogtanh_sel( Ief209532f4cbf1c6a41bea414577f825[flogtanh_SEL-1:0]),
.flogtanh( I2dacd37cecd93c6e9134cb55ed917d78),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I88aedd7f52399f5fd435c3415f2218ca = (Ief209532f4cbf1c6a41bea414577f825[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2dacd37cecd93c6e9134cb55ed917d78;


Ic3da32f100a43f826b89a492544e7812 I576b5a8b10944760f3e55d1b03e9d19f (
.flogtanh_sel( I1c8953ad3f64f3c3cc506808aad29dab[flogtanh_SEL-1:0]),
.flogtanh( I2419bc316181acd41e29ad005241d812),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7651176b0a74846108fbaabc5cc4900a = (I1c8953ad3f64f3c3cc506808aad29dab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2419bc316181acd41e29ad005241d812;


Ic3da32f100a43f826b89a492544e7812 I4bccc68d2cd1c59e701eb9b8c5f3cf70 (
.flogtanh_sel( I1b519d88bbf86cfb080a50ea0480a128[flogtanh_SEL-1:0]),
.flogtanh( I35faf0af91f4972ae843883993fc84f4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I57ac487adc18165136e9b3c7c50f95ad = (I1b519d88bbf86cfb080a50ea0480a128[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I35faf0af91f4972ae843883993fc84f4;


Ic3da32f100a43f826b89a492544e7812 I8d5cd2bb516fa5bc6f5fd684fa6d2ce1 (
.flogtanh_sel( I5b8258f35d889071109216b464abb2a4[flogtanh_SEL-1:0]),
.flogtanh( I4dd2e7b6a685958d7aac77a38354e05f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic95668328a2121027436f682bac50b9c = (I5b8258f35d889071109216b464abb2a4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4dd2e7b6a685958d7aac77a38354e05f;


Ic3da32f100a43f826b89a492544e7812 I4142f6d5b9f94a60dc4c93f0c1a5e4ab (
.flogtanh_sel( Id9681d4e0e4d375f9279de115a4337a3[flogtanh_SEL-1:0]),
.flogtanh( Ib27460a2e2b13abc54f5ba37f32c8653),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I118726375ca9381e45f001965fcefc5b = (Id9681d4e0e4d375f9279de115a4337a3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib27460a2e2b13abc54f5ba37f32c8653;


Ic3da32f100a43f826b89a492544e7812 I22b6308113e975a22426ff3a2aa88296 (
.flogtanh_sel( Ib42144ece00b82debd70011724a29c91[flogtanh_SEL-1:0]),
.flogtanh( Ia3fa91387788798672eb6199a2eaa389),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic8d47ff5d6c31601a57df868da78c2d4 = (Ib42144ece00b82debd70011724a29c91[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia3fa91387788798672eb6199a2eaa389;


Ic3da32f100a43f826b89a492544e7812 I539bb7fc15c6311b643230dcbce52d5c (
.flogtanh_sel( Ic5717058a1815f63f164de1b1defe8cb[flogtanh_SEL-1:0]),
.flogtanh( Ieecd194ccc5698a2ba16efd969cfd621),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7cdc5ada6fc68ee31fd4062e2ff004d3 = (Ic5717058a1815f63f164de1b1defe8cb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieecd194ccc5698a2ba16efd969cfd621;


Ic3da32f100a43f826b89a492544e7812 I2fa2d9bec1881c9e6cd52d1d171e0ebf (
.flogtanh_sel( Iea41672f012f225d64d9c75b198c812f[flogtanh_SEL-1:0]),
.flogtanh( Ifb09fa1840c5a1ddbfc81cda21c11f1e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I59547aacdcfde31dc016ec2acbb2f4b4 = (Iea41672f012f225d64d9c75b198c812f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifb09fa1840c5a1ddbfc81cda21c11f1e;


Ic3da32f100a43f826b89a492544e7812 I43e111ddfbf6e973763f3a841b83d1aa (
.flogtanh_sel( I7a070bd014e1d2c5e55e5fcba88a5664[flogtanh_SEL-1:0]),
.flogtanh( I4ce505ae2025bab3abcf5a44e0ed5034),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia7f53f0cd86055da72c13ac474f052a1 = (I7a070bd014e1d2c5e55e5fcba88a5664[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4ce505ae2025bab3abcf5a44e0ed5034;


Ic3da32f100a43f826b89a492544e7812 Ia72461665ae08e77c1b7bc2239fdc2a2 (
.flogtanh_sel( I4a0a8b28429b708363458c74230b0fc2[flogtanh_SEL-1:0]),
.flogtanh( Id40a7ca1cde7a70cc13e752e19132808),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I915054f2fbb8b93516d8748a3e3e29e2 = (I4a0a8b28429b708363458c74230b0fc2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id40a7ca1cde7a70cc13e752e19132808;


Ic3da32f100a43f826b89a492544e7812 I8377ea96a183b52f5f45dff233e27c13 (
.flogtanh_sel( If585e4075ac1740f3b141ae6a50200f7[flogtanh_SEL-1:0]),
.flogtanh( If7274be2bcc8b2a235c3538db5506d90),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If257757fa31c2f4cc9ec322e4ecccf83 = (If585e4075ac1740f3b141ae6a50200f7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If7274be2bcc8b2a235c3538db5506d90;


Ic3da32f100a43f826b89a492544e7812 I8f0022371d98c4d87d0810697a286dbd (
.flogtanh_sel( Ie1a68cf09bb21a1629369fde87f51bea[flogtanh_SEL-1:0]),
.flogtanh( I3e611982ec9ff6437f22e11b2552693a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If91268e2b84df18785cd6a53e53eb4e9 = (Ie1a68cf09bb21a1629369fde87f51bea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3e611982ec9ff6437f22e11b2552693a;


Ic3da32f100a43f826b89a492544e7812 Id115eead151f333caac671bc2246405c (
.flogtanh_sel( I72b8547125d0ad6c1ad39a68b55c818c[flogtanh_SEL-1:0]),
.flogtanh( I8fcf0a468234f365c33059e26b9f5821),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia072f1d679429d3c3180f8eb67fc7dd7 = (I72b8547125d0ad6c1ad39a68b55c818c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8fcf0a468234f365c33059e26b9f5821;


Ic3da32f100a43f826b89a492544e7812 I249aa48ac54bb2cefcb82f59ae1a5589 (
.flogtanh_sel( Ie14ba4a8657740f9a8d057258db2cb09[flogtanh_SEL-1:0]),
.flogtanh( I3f80250ee19e8250898f2bcc055c2e5b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I91a8168d3b087ab3891cd6d479427b95 = (Ie14ba4a8657740f9a8d057258db2cb09[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3f80250ee19e8250898f2bcc055c2e5b;


Ic3da32f100a43f826b89a492544e7812 Id7a739526603a60ea5134d57b191e876 (
.flogtanh_sel( I27490a69fb2a1f6f298639254c37cf9e[flogtanh_SEL-1:0]),
.flogtanh( I06b3652935db14aaa057f0cf3cffef66),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id1dce8c1542f1279badb381aca3c9b51 = (I27490a69fb2a1f6f298639254c37cf9e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I06b3652935db14aaa057f0cf3cffef66;


Ic3da32f100a43f826b89a492544e7812 I8d6ad838171c25056f78ff7b6050a4f5 (
.flogtanh_sel( I49b9c212fbe74a5dd8b087e417296186[flogtanh_SEL-1:0]),
.flogtanh( Ib01d30e88a3a1fcb204246baafeb47c8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8983f003c30a218543f39f5bbcd9a25c = (I49b9c212fbe74a5dd8b087e417296186[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib01d30e88a3a1fcb204246baafeb47c8;


Ic3da32f100a43f826b89a492544e7812 I695ea24b9833ec81c2700667d6c9afff (
.flogtanh_sel( I0a8e6f5cc8b6ea599b7605abe6479bec[flogtanh_SEL-1:0]),
.flogtanh( I9f688c58878405d1d2865ddc40659c2b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id1b5c33bc63f75561b7cce6fc0981c69 = (I0a8e6f5cc8b6ea599b7605abe6479bec[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f688c58878405d1d2865ddc40659c2b;


Ic3da32f100a43f826b89a492544e7812 Ic5a3e4b327f2c57a11532341580e737d (
.flogtanh_sel( Ib6d94b34d3886717e4016fec196f277f[flogtanh_SEL-1:0]),
.flogtanh( Ic9c77123914f831cee5bc4586b6a2a8b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I003f95fb8f2027efa41a1936e8b53986 = (Ib6d94b34d3886717e4016fec196f277f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic9c77123914f831cee5bc4586b6a2a8b;


Ic3da32f100a43f826b89a492544e7812 If58650b220f1aa2f30645fddcb1fb11f (
.flogtanh_sel( Id7e53d36da7171e036ebfc984dbcea6e[flogtanh_SEL-1:0]),
.flogtanh( Ifd42760504e0f106eb9061d9b9a2d18a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie16dc913f571ae73ce03d755077345a9 = (Id7e53d36da7171e036ebfc984dbcea6e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifd42760504e0f106eb9061d9b9a2d18a;


Ic3da32f100a43f826b89a492544e7812 I556226325c13e5f4e8eae7e44ad07672 (
.flogtanh_sel( I2ec254d80fd0683d782302cf3839559b[flogtanh_SEL-1:0]),
.flogtanh( I452794105cca79653f5509dac3794327),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I86e53eed5b857c439039238bb486067c = (I2ec254d80fd0683d782302cf3839559b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I452794105cca79653f5509dac3794327;


Ic3da32f100a43f826b89a492544e7812 I5945efcaa4e3b34c8355cf891628005e (
.flogtanh_sel( Ibbedaef61051d5df82cd6d55e05c80da[flogtanh_SEL-1:0]),
.flogtanh( I33431ed9c549f5525adfa5d45fbc7653),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I89433799cfa534afd66e8d6b9f1b62b9 = (Ibbedaef61051d5df82cd6d55e05c80da[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I33431ed9c549f5525adfa5d45fbc7653;


Ic3da32f100a43f826b89a492544e7812 I26e43752cc552ec07af0c5d30d07ff1c (
.flogtanh_sel( I501336bb7ba172c05dd5840036e6228c[flogtanh_SEL-1:0]),
.flogtanh( I4b8b4fd334b176cb449ad0296ebff4c8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I80f2e8f6743e28e86e4d85b295e2f768 = (I501336bb7ba172c05dd5840036e6228c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4b8b4fd334b176cb449ad0296ebff4c8;


Ic3da32f100a43f826b89a492544e7812 I5908a81d7dc254c7494055dc4e1009a8 (
.flogtanh_sel( I8e5c4c6c63e42054359cee697cc0d026[flogtanh_SEL-1:0]),
.flogtanh( I66e7dacba9dbfb14e9a71b9d57229880),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1391018fb93372ccc2fcc08700e38b65 = (I8e5c4c6c63e42054359cee697cc0d026[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I66e7dacba9dbfb14e9a71b9d57229880;


Ic3da32f100a43f826b89a492544e7812 I08c4e21da618ed476ce198f617ab1037 (
.flogtanh_sel( Id3daa6db921871b752bf92366446afcc[flogtanh_SEL-1:0]),
.flogtanh( If3a842c52c8c0b2fd24ef265e8cfe330),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8fd26d47ecd4cdd08294cf6133468d17 = (Id3daa6db921871b752bf92366446afcc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If3a842c52c8c0b2fd24ef265e8cfe330;


Ic3da32f100a43f826b89a492544e7812 Id4908ceaa69811b0701028333bf95f29 (
.flogtanh_sel( Id8367ec60787bfad0da8aa76c6ed8ddb[flogtanh_SEL-1:0]),
.flogtanh( I0f3aea4265966e7bc673d3a08ad1c2e4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7097c9518bb3351818b96f31ed49c6d3 = (Id8367ec60787bfad0da8aa76c6ed8ddb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0f3aea4265966e7bc673d3a08ad1c2e4;


Ic3da32f100a43f826b89a492544e7812 I431e1976feff5d3ce21ca3752889e789 (
.flogtanh_sel( I533649312ec995f1f9e514c59a8675b1[flogtanh_SEL-1:0]),
.flogtanh( Ia9de78211d220e68835ff757eb75d919),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id683d693cd50645c3d6d657aa1c8bdb2 = (I533649312ec995f1f9e514c59a8675b1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia9de78211d220e68835ff757eb75d919;


Ic3da32f100a43f826b89a492544e7812 I5bb1267e5f11b9a4c5e016687956a2f2 (
.flogtanh_sel( I0621d0b2c83e70b4afd65eb9dca4b514[flogtanh_SEL-1:0]),
.flogtanh( I2c1c31b8bda73b145cdf74b18bc46a4d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I88bd8012c93dd9e2ed52ea5e9b8b0004 = (I0621d0b2c83e70b4afd65eb9dca4b514[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2c1c31b8bda73b145cdf74b18bc46a4d;


Ic3da32f100a43f826b89a492544e7812 Idde7213ca7df10e15005410ced8b12d7 (
.flogtanh_sel( I2ae01892a3cd0432618d7280b31daddb[flogtanh_SEL-1:0]),
.flogtanh( I300a84deada851e18835d6af55c5e2a3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia8d3667adc34b2b50acf7edb970538d8 = (I2ae01892a3cd0432618d7280b31daddb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I300a84deada851e18835d6af55c5e2a3;


Ic3da32f100a43f826b89a492544e7812 Ideb80dfeff3fee14ce62c76ea51ff4cb (
.flogtanh_sel( I5ed8a2f30bd2ea269341c2267ae3fe83[flogtanh_SEL-1:0]),
.flogtanh( I1fc6745ba86be641dc9bdac044c19519),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3f0bba472e912f11dea8e788fbc1cb63 = (I5ed8a2f30bd2ea269341c2267ae3fe83[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1fc6745ba86be641dc9bdac044c19519;


Ic3da32f100a43f826b89a492544e7812 Ibe707c5b40237213c8941856a92075c1 (
.flogtanh_sel( I2c819e7f62c0dc0aac650074b203163b[flogtanh_SEL-1:0]),
.flogtanh( I2791cc5f69dd0e7f306760048c759af7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6dc671e73b4e9c70cabfdeaac2e5c40b = (I2c819e7f62c0dc0aac650074b203163b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2791cc5f69dd0e7f306760048c759af7;


Ic3da32f100a43f826b89a492544e7812 I29b3b56d98b2e8ba2f00e6415da9ad0f (
.flogtanh_sel( I30e20b58913d6fbe5817e1956ba8e570[flogtanh_SEL-1:0]),
.flogtanh( Ie8157cde860052619820431f87e13c83),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia6255a136d5f36ea6cba654bd5823850 = (I30e20b58913d6fbe5817e1956ba8e570[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie8157cde860052619820431f87e13c83;


Ic3da32f100a43f826b89a492544e7812 I89e5718376d68fc5046b3352835a043b (
.flogtanh_sel( I1b922bed7f3c4a6705f3ce7a885a68cd[flogtanh_SEL-1:0]),
.flogtanh( I9059b74a8f3cf2e4905756cc9c71597f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2b9584392ef9a7828ff57bd4c522a302 = (I1b922bed7f3c4a6705f3ce7a885a68cd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9059b74a8f3cf2e4905756cc9c71597f;


Ic3da32f100a43f826b89a492544e7812 I844c5af5dac16f69bea6678d32514674 (
.flogtanh_sel( I2f65f0917713ecc8585392d3b557c1bf[flogtanh_SEL-1:0]),
.flogtanh( I99584eabd3cbd2546c85f474afa6fabb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6c1235e88ae444a96ea64fd1bfd04d8f = (I2f65f0917713ecc8585392d3b557c1bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I99584eabd3cbd2546c85f474afa6fabb;


Ic3da32f100a43f826b89a492544e7812 I0007b912587020b21a5db1485f1dcbb7 (
.flogtanh_sel( I3301533e7d9e527118a67c462f1b4357[flogtanh_SEL-1:0]),
.flogtanh( I047abade6abf10a65a5b835ac725fa7c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id09b8242c22851fb960d55222fe733d4 = (I3301533e7d9e527118a67c462f1b4357[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I047abade6abf10a65a5b835ac725fa7c;


Ic3da32f100a43f826b89a492544e7812 I41f5da9e92bb6340e65d2ddbf1c80d73 (
.flogtanh_sel( I52a88bdb1f03da82730f7579b7b5305d[flogtanh_SEL-1:0]),
.flogtanh( Icf7ab1d1113bc44358c56a56fca7caf9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie355fa27abbc41291eaf08f2cf9a6ff7 = (I52a88bdb1f03da82730f7579b7b5305d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icf7ab1d1113bc44358c56a56fca7caf9;


Ic3da32f100a43f826b89a492544e7812 I6f39119549e922a0cc32c68620a366e5 (
.flogtanh_sel( I644c730662b3725d26cd46fb46106104[flogtanh_SEL-1:0]),
.flogtanh( I4d24650be7a1088c2310d93000d6392a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I566224393f6bb27bfd8b0b0d6b8e53d6 = (I644c730662b3725d26cd46fb46106104[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4d24650be7a1088c2310d93000d6392a;


Ic3da32f100a43f826b89a492544e7812 Ifb2f9f03ebebe325c5a41668f27caf99 (
.flogtanh_sel( I3da3e36c76c4123bec6879bccb39e933[flogtanh_SEL-1:0]),
.flogtanh( Ic3aea8ebb8eab44a92e7d7d950e1a917),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8fcad6e7d5ffc9f79eaaf634f6fe8cda = (I3da3e36c76c4123bec6879bccb39e933[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic3aea8ebb8eab44a92e7d7d950e1a917;


Ic3da32f100a43f826b89a492544e7812 Iacfb3765fecc5929f30cdfbeacf10db6 (
.flogtanh_sel( Iebde55cddc8170f7dd8855ea55eff0ce[flogtanh_SEL-1:0]),
.flogtanh( I82af0956870500474eac2505bbf15e35),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6f0f74dcc830fdcb0af9df75a2b722f7 = (Iebde55cddc8170f7dd8855ea55eff0ce[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I82af0956870500474eac2505bbf15e35;


Ic3da32f100a43f826b89a492544e7812 I65f19cf8bc0deff06a3691d818ff1fab (
.flogtanh_sel( Ie673e2d92a7090b2fa1c5e14a2e03be3[flogtanh_SEL-1:0]),
.flogtanh( I2d8a8efaa0179340bf5d3ebbd4c11831),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idd95fd099dd2b53c46d02f09575b8032 = (Ie673e2d92a7090b2fa1c5e14a2e03be3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2d8a8efaa0179340bf5d3ebbd4c11831;


Ic3da32f100a43f826b89a492544e7812 I3871f6c8800fbc4edc60686de9107100 (
.flogtanh_sel( If90afe75714f8660ad0eb9f9ea06cd6b[flogtanh_SEL-1:0]),
.flogtanh( I32ff895ff659ec448270067f76e97a90),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0f277bc88d46a4e6e9f1f2c410b503fd = (If90afe75714f8660ad0eb9f9ea06cd6b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I32ff895ff659ec448270067f76e97a90;


Ic3da32f100a43f826b89a492544e7812 I0d9e31b2ee6b243e49354cde278f0362 (
.flogtanh_sel( Ifd96e3a6e0050c30a4308328cfecb21f[flogtanh_SEL-1:0]),
.flogtanh( I15a7fd79aeb5eed24b1c7be3d48296e0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I66b92f1de2cf408c3af53b161a6ffa60 = (Ifd96e3a6e0050c30a4308328cfecb21f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I15a7fd79aeb5eed24b1c7be3d48296e0;


Ic3da32f100a43f826b89a492544e7812 Iddffa69325221e415b4e93fbafce33b9 (
.flogtanh_sel( I68b92cc2d83e9a718edd2aea82314016[flogtanh_SEL-1:0]),
.flogtanh( I12f311f2311e26320a178d6fec95d9d0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id28d9545e8d20ac080fbac5e345692da = (I68b92cc2d83e9a718edd2aea82314016[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I12f311f2311e26320a178d6fec95d9d0;


Ic3da32f100a43f826b89a492544e7812 I6953819e3f7ed90649124e21a06eb08b (
.flogtanh_sel( I6bdbb92363f0e072ed04654e9aad17a5[flogtanh_SEL-1:0]),
.flogtanh( I2b8ce30d1338ad506e4996d2dd1dc11a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4a5cfd6ebd47cda4fa2e06ba9ad6e5b2 = (I6bdbb92363f0e072ed04654e9aad17a5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2b8ce30d1338ad506e4996d2dd1dc11a;


Ic3da32f100a43f826b89a492544e7812 I144a1f3e4197275d0956b9becba5a51a (
.flogtanh_sel( I87a4267db59b97ef1b9bca8743cb0322[flogtanh_SEL-1:0]),
.flogtanh( Ic2b65e7bd42e94f2ad8b6506a6fce7af),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I62bda8dc70e0b5eb38abe094bbe92fc6 = (I87a4267db59b97ef1b9bca8743cb0322[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic2b65e7bd42e94f2ad8b6506a6fce7af;


Ic3da32f100a43f826b89a492544e7812 I2add9cddab0895bf0e7d01fea3eef533 (
.flogtanh_sel( I44eacb2bea725efab7c0dd560279f0f8[flogtanh_SEL-1:0]),
.flogtanh( I0f54a697ea3e2bbf90354c9a6173fb80),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I223b05d94c09b095d1988df121aa5e37 = (I44eacb2bea725efab7c0dd560279f0f8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0f54a697ea3e2bbf90354c9a6173fb80;


Ic3da32f100a43f826b89a492544e7812 Iaa70a21eb0f3ca1e51d63f9ff8d3b40a (
.flogtanh_sel( I87a2736466c5ee62b7cc55f17e715ffa[flogtanh_SEL-1:0]),
.flogtanh( I6a6c0f8e4399c21285d66ddc0f1f70c0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5f73e5faf1aca83ee0a415c9ac4a1b9a = (I87a2736466c5ee62b7cc55f17e715ffa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6a6c0f8e4399c21285d66ddc0f1f70c0;


Ic3da32f100a43f826b89a492544e7812 I50003562d145e8a896129b6585b3cc9f (
.flogtanh_sel( I7a66c7713ba126fdc24940cd92f7e10b[flogtanh_SEL-1:0]),
.flogtanh( Ibfcdfc01f09bcff031e359394947efef),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I75f9d3a41019dca3044a1c2cf7069662 = (I7a66c7713ba126fdc24940cd92f7e10b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibfcdfc01f09bcff031e359394947efef;


Ic3da32f100a43f826b89a492544e7812 Ibbf69218236c464b42dce0698c095c6b (
.flogtanh_sel( I1f11c579f34c41aade41c53f53468057[flogtanh_SEL-1:0]),
.flogtanh( I8efd478f1ae2ea6090774e1ed3bd7b28),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I820fa56328e3919970dd64adb1d4d8e7 = (I1f11c579f34c41aade41c53f53468057[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8efd478f1ae2ea6090774e1ed3bd7b28;


Ic3da32f100a43f826b89a492544e7812 Ie0415709fdff5c060ab931ba2565a70d (
.flogtanh_sel( I651a438f70583d476ae10f066e035435[flogtanh_SEL-1:0]),
.flogtanh( I502d3210c60c82ca682d8e2168d54be0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I05eadf11cdc6c2f2b021e33f2438fa49 = (I651a438f70583d476ae10f066e035435[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I502d3210c60c82ca682d8e2168d54be0;


Ic3da32f100a43f826b89a492544e7812 I85165873bd6afdef91d39b7b974764c8 (
.flogtanh_sel( Ibdf17fa73794c846e15fe0a915b071e5[flogtanh_SEL-1:0]),
.flogtanh( I337d74c3c773a358a936806f751c1117),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2c487770d606451440eecf358202db32 = (Ibdf17fa73794c846e15fe0a915b071e5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I337d74c3c773a358a936806f751c1117;


Ic3da32f100a43f826b89a492544e7812 I24018d3b466c111ae047548bf961ef5b (
.flogtanh_sel( I76d3221fbcefc0ee08655f7ba4919f3c[flogtanh_SEL-1:0]),
.flogtanh( Ia494fdbd70bff11510eb685f3b5d0aae),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I082aa8c413d7ef8f054b1c2857cbe39f = (I76d3221fbcefc0ee08655f7ba4919f3c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia494fdbd70bff11510eb685f3b5d0aae;


Ic3da32f100a43f826b89a492544e7812 Iff069ca9a50cf40acf0d2efc56337fc5 (
.flogtanh_sel( I3458f69c90ea8b20b3d1f67e9a13ec2e[flogtanh_SEL-1:0]),
.flogtanh( I547f7a4c3801c1caa4587c9aef397652),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I420e2c5a8745133f6263a71b458f1e2f = (I3458f69c90ea8b20b3d1f67e9a13ec2e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I547f7a4c3801c1caa4587c9aef397652;


Ic3da32f100a43f826b89a492544e7812 Iffcb8b2b0a0b8934faa0724bc37d5869 (
.flogtanh_sel( Ia2d6e9e1e92a30c7028af50ddfbb9bf9[flogtanh_SEL-1:0]),
.flogtanh( I8009d84fd826dd21eb7091744792f4a7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4b8d520ee88fd39d83a16432e962f731 = (Ia2d6e9e1e92a30c7028af50ddfbb9bf9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8009d84fd826dd21eb7091744792f4a7;


Ic3da32f100a43f826b89a492544e7812 I38ff7e3b1a8cee39d465c440a14bc20d (
.flogtanh_sel( I66c91b5133d9812a03daecc0b14211f8[flogtanh_SEL-1:0]),
.flogtanh( If724b1c92350989910925d275353e544),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia3f7f07ddb09ea33218afe14281ac3c6 = (I66c91b5133d9812a03daecc0b14211f8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If724b1c92350989910925d275353e544;


Ic3da32f100a43f826b89a492544e7812 Ief4f8b2268e627243f72af96ea365b75 (
.flogtanh_sel( Ifb5986949e88167526d9fcfe07b417ca[flogtanh_SEL-1:0]),
.flogtanh( I26f4a180e992f5de04bc047f539bcb48),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I25aefb53f59a00abe88b9dcf6be6907a = (Ifb5986949e88167526d9fcfe07b417ca[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I26f4a180e992f5de04bc047f539bcb48;


Ic3da32f100a43f826b89a492544e7812 Ia9f8d88326fd0e2d4df547de180c8c83 (
.flogtanh_sel( Iedada801ca6cd173ee523ef335e91ff6[flogtanh_SEL-1:0]),
.flogtanh( I83ca10d71caf5ac98fef3d45d228be8e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I22c3140a8db02352d2e2a2a11eeba117 = (Iedada801ca6cd173ee523ef335e91ff6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I83ca10d71caf5ac98fef3d45d228be8e;


Ic3da32f100a43f826b89a492544e7812 I5eb5a8692051256ef289026a6361ba1e (
.flogtanh_sel( I4e2722e547586da7565b2d91a7fc91e7[flogtanh_SEL-1:0]),
.flogtanh( Ib8407faa17d1e96cd317c65459c4fa71),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I954dd66f60316803a8f13a39c460a39a = (I4e2722e547586da7565b2d91a7fc91e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib8407faa17d1e96cd317c65459c4fa71;


Ic3da32f100a43f826b89a492544e7812 Iacbf6f018b3b1b2820c5263e1606962e (
.flogtanh_sel( Ib321a8ceda62c64ab25dc1c718301bda[flogtanh_SEL-1:0]),
.flogtanh( I73829d98e5e2f368c4a2020e3d7814be),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I37b3988d699a1ed42923e3fd1584ecc0 = (Ib321a8ceda62c64ab25dc1c718301bda[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I73829d98e5e2f368c4a2020e3d7814be;


Ic3da32f100a43f826b89a492544e7812 I0091774807a9b33730d198c2715358a2 (
.flogtanh_sel( I58daeebec4873e6c1c07c090ff81235c[flogtanh_SEL-1:0]),
.flogtanh( I9a120c441f8d9ccb617057e042587ba1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If79bc5a35cb55036a367efb88c7d5510 = (I58daeebec4873e6c1c07c090ff81235c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9a120c441f8d9ccb617057e042587ba1;


Ic3da32f100a43f826b89a492544e7812 If0cd9254572357e9af6a7ad69e7160d4 (
.flogtanh_sel( I3f103fbbe49c86c9db46129bd4632cab[flogtanh_SEL-1:0]),
.flogtanh( I8064df8bc33998ad58d460afae699e48),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ideab06dc2448a6950cd1a06a0c90c2c6 = (I3f103fbbe49c86c9db46129bd4632cab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8064df8bc33998ad58d460afae699e48;


Ic3da32f100a43f826b89a492544e7812 I6b80c6ab37f5b005cbdca0c7237a2f63 (
.flogtanh_sel( Id6697ca17f1bd6ddd112951b9d89a8ea[flogtanh_SEL-1:0]),
.flogtanh( If016e079d3b453444558706ef9073233),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1d7d7a68fc53b8be89c4637ac8f29380 = (Id6697ca17f1bd6ddd112951b9d89a8ea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If016e079d3b453444558706ef9073233;


Ic3da32f100a43f826b89a492544e7812 I1b8697cb2079bee1d0ae4d83e3152eac (
.flogtanh_sel( I445ede2983c7470b4418a2ec0cbbd5e1[flogtanh_SEL-1:0]),
.flogtanh( I51cc187d91ee3c480a759104aed41b1b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib34ad1d14978608d1440f59998a31672 = (I445ede2983c7470b4418a2ec0cbbd5e1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I51cc187d91ee3c480a759104aed41b1b;


Ic3da32f100a43f826b89a492544e7812 I62e574584c02081525296f9521df1dd0 (
.flogtanh_sel( I034e56cd77ee400ed81b78177b202930[flogtanh_SEL-1:0]),
.flogtanh( I4b8068a6a866c2424439b2956245ac8d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id081512cd113e4d09df0fb13e443d76b = (I034e56cd77ee400ed81b78177b202930[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4b8068a6a866c2424439b2956245ac8d;


Ic3da32f100a43f826b89a492544e7812 I0c31c19531b2665b9917ec4138a2c321 (
.flogtanh_sel( I08edadbd9366786f96b44268d096b4aa[flogtanh_SEL-1:0]),
.flogtanh( I60513d924016bd300559b7a1bea7f521),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I57a0f8c3710cf8e216d6dc2420f7621c = (I08edadbd9366786f96b44268d096b4aa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I60513d924016bd300559b7a1bea7f521;


Ic3da32f100a43f826b89a492544e7812 I82bc8a5240e5dd2a68fe218564a6c3a7 (
.flogtanh_sel( I8f86a7af86eb04c5df18e09888cdce7b[flogtanh_SEL-1:0]),
.flogtanh( Iec98284ab12724bb63360f29d00f1ecb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaa164a078c8cdaad694a053c9c1e0313 = (I8f86a7af86eb04c5df18e09888cdce7b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iec98284ab12724bb63360f29d00f1ecb;


Ic3da32f100a43f826b89a492544e7812 I167e26920b27dd3e47e116a6bb17fef4 (
.flogtanh_sel( Ic00d037a11f8a27ab34e4daab8c9c2e6[flogtanh_SEL-1:0]),
.flogtanh( I3e3eba8135eb797d0a5e8ac1feefce0c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7eb76b3d17296fdae702d8f820f1428d = (Ic00d037a11f8a27ab34e4daab8c9c2e6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3e3eba8135eb797d0a5e8ac1feefce0c;


Ic3da32f100a43f826b89a492544e7812 I9fed361ab5dce82d062a2216fd7c423c (
.flogtanh_sel( I4d95ceccc6c3ad37f13c98339c59e5c4[flogtanh_SEL-1:0]),
.flogtanh( I6aa98bc7265b8b7c25181a06e75c24c0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I00ecb5e329390023b318a2ceba0df231 = (I4d95ceccc6c3ad37f13c98339c59e5c4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6aa98bc7265b8b7c25181a06e75c24c0;


Ic3da32f100a43f826b89a492544e7812 I2ce031496545060b3d3a9fd71101242a (
.flogtanh_sel( I1ea967d377f462a0e06d7d0d4d95b342[flogtanh_SEL-1:0]),
.flogtanh( I47f9c7018999e1cea25feddbe399e6b7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iea32ebc385c6cfc9212ff37973a0a05d = (I1ea967d377f462a0e06d7d0d4d95b342[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I47f9c7018999e1cea25feddbe399e6b7;


Ic3da32f100a43f826b89a492544e7812 I42725bbb1b731e35d6515a1dab325e2e (
.flogtanh_sel( Ib0feec63123e66bd6ad6935e9b7fa6bf[flogtanh_SEL-1:0]),
.flogtanh( I7224803ba8f0a16a7b2e969fe727bfa1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If845af0d620024f04525244753ba5d18 = (Ib0feec63123e66bd6ad6935e9b7fa6bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7224803ba8f0a16a7b2e969fe727bfa1;


Ic3da32f100a43f826b89a492544e7812 Ibf16dd7e31d580e0d6a40478aa5e5aab (
.flogtanh_sel( I7d120060ddae9ff8f7206b3ef63eda50[flogtanh_SEL-1:0]),
.flogtanh( I65bc4e0d837f94c4301cb2c87e24969c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I08e907b0619bec3ef2cf4cb3779e0794 = (I7d120060ddae9ff8f7206b3ef63eda50[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I65bc4e0d837f94c4301cb2c87e24969c;


Ic3da32f100a43f826b89a492544e7812 I5f2056e011411b04b0a398bb9405539d (
.flogtanh_sel( Ib47f8f72386e2e65a88fbadd3a705225[flogtanh_SEL-1:0]),
.flogtanh( I444f8e61602b8994f7a01f3ebd4ac6ab),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I68e5b12792a86dda0576742831d3b728 = (Ib47f8f72386e2e65a88fbadd3a705225[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I444f8e61602b8994f7a01f3ebd4ac6ab;


Ic3da32f100a43f826b89a492544e7812 I7926aaccdd9186d8ae8feabf86f4ba6e (
.flogtanh_sel( I4e0efc35346e2934f5bb4c34a4bc5f90[flogtanh_SEL-1:0]),
.flogtanh( I86c51ec7ff965132e195835d21c24881),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I72db05084d30d7c59ba1cb06d3b09400 = (I4e0efc35346e2934f5bb4c34a4bc5f90[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I86c51ec7ff965132e195835d21c24881;


Ic3da32f100a43f826b89a492544e7812 Ie562558b900fdb10c62443284b212a0d (
.flogtanh_sel( I3ca1014802f58087e3434a1e0df19c01[flogtanh_SEL-1:0]),
.flogtanh( I07aa1b2db5dedc3230dff10534311a56),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib1f1aef6c0a9291553b62fd555feb2e7 = (I3ca1014802f58087e3434a1e0df19c01[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I07aa1b2db5dedc3230dff10534311a56;


Ic3da32f100a43f826b89a492544e7812 I534db043ec9bced4e4cd89ab8e2c979c (
.flogtanh_sel( I688a3879b7be1544e6f94b4221c03213[flogtanh_SEL-1:0]),
.flogtanh( Ia8809cc89c377e8b4109cdc8976daa54),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib504b808f724ca6032e7c746517cd4fd = (I688a3879b7be1544e6f94b4221c03213[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia8809cc89c377e8b4109cdc8976daa54;


Ic3da32f100a43f826b89a492544e7812 Ie2e9328666f6a9ab4574b027a90c3f4d (
.flogtanh_sel( Ic22988138610c8671ec342f65f34c7ae[flogtanh_SEL-1:0]),
.flogtanh( I7402dc21bfbc0af749dd8fb03c516a50),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia47f7fb27f2d965cfd2989569c257356 = (Ic22988138610c8671ec342f65f34c7ae[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7402dc21bfbc0af749dd8fb03c516a50;


Ic3da32f100a43f826b89a492544e7812 Ib7a4cc99196d24ab8c97d7ed0c36f037 (
.flogtanh_sel( I0b85fdd83569e5cbb7d71eed50cb32fd[flogtanh_SEL-1:0]),
.flogtanh( I8ca06f4250a69dde75889f7a6ba3f456),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If2b17f9e9186542117f43d0dd342326e = (I0b85fdd83569e5cbb7d71eed50cb32fd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8ca06f4250a69dde75889f7a6ba3f456;


Ic3da32f100a43f826b89a492544e7812 If486121eb56046f5f35c266cf308eb47 (
.flogtanh_sel( Idf55390c11e5b41ebc2a28e0af109913[flogtanh_SEL-1:0]),
.flogtanh( Ibab00faeaa6a7be99fa6a239193b92cb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6c4ba0863ab4c8d1a56324a4d89ccbeb = (Idf55390c11e5b41ebc2a28e0af109913[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibab00faeaa6a7be99fa6a239193b92cb;


Ic3da32f100a43f826b89a492544e7812 I78909a9fd4bbca430d67a8206349c75a (
.flogtanh_sel( I6b48935ea25672ee9a42f49eae9e519f[flogtanh_SEL-1:0]),
.flogtanh( I8e44b109466e00487db9dfb7ae225f89),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4dbd1bb8f1641f15e3a4f1e309962811 = (I6b48935ea25672ee9a42f49eae9e519f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8e44b109466e00487db9dfb7ae225f89;


Ic3da32f100a43f826b89a492544e7812 Ie680eb56732b53bd6c339272c65bbd8d (
.flogtanh_sel( I6a9e6c39c20e45773dab7823a7ff9486[flogtanh_SEL-1:0]),
.flogtanh( Ib3e38e46bfa9e1bdc032918269223b32),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I26781ef851ed43c6f88ff1215cddca6b = (I6a9e6c39c20e45773dab7823a7ff9486[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib3e38e46bfa9e1bdc032918269223b32;


Ic3da32f100a43f826b89a492544e7812 I716d5daaa09e44ee38ec699d3a20e73c (
.flogtanh_sel( I42907182010c5889ddb7a700ead16525[flogtanh_SEL-1:0]),
.flogtanh( I659fb1602b9d248940523c14c628ce86),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia349e1f7c10a63ddccb3f300c73b4572 = (I42907182010c5889ddb7a700ead16525[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I659fb1602b9d248940523c14c628ce86;


Ic3da32f100a43f826b89a492544e7812 Ia18623b2774c469fb5ddf3d9fd4a272a (
.flogtanh_sel( Ib6c26f3e3358cc2ed6fbda83eabd4bd3[flogtanh_SEL-1:0]),
.flogtanh( I1a264a901911abed928628d819c162b2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I50c4e1d3a3f63b93bc36b5141226fb3c = (Ib6c26f3e3358cc2ed6fbda83eabd4bd3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1a264a901911abed928628d819c162b2;


Ic3da32f100a43f826b89a492544e7812 I3ff3832352e96aa008336b4504c1d7a0 (
.flogtanh_sel( Ia50d85808790790450f87a5246874b3f[flogtanh_SEL-1:0]),
.flogtanh( I2a53bd293919bc846ab816144b42592a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I12334038c2be8634c47869f397503019 = (Ia50d85808790790450f87a5246874b3f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2a53bd293919bc846ab816144b42592a;


Ic3da32f100a43f826b89a492544e7812 I478b79b5f293cdbc4f3ea64690fda119 (
.flogtanh_sel( Id4a1744702d7808a80bc40697c864765[flogtanh_SEL-1:0]),
.flogtanh( I35ce9e616a3213f2b4ce0597a47f998c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I64692d5168554dfd7ce1c7a046aecf72 = (Id4a1744702d7808a80bc40697c864765[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I35ce9e616a3213f2b4ce0597a47f998c;


Ic3da32f100a43f826b89a492544e7812 I336dbe5b756c3f17e37499b4e99c8c2a (
.flogtanh_sel( I0cf3d2f3e6793a2dcf15949da16ad28d[flogtanh_SEL-1:0]),
.flogtanh( Ic3f28aa77fc84cb8e2fe43bac7ede253),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia4b438844530fff602ea04e72b07db8d = (I0cf3d2f3e6793a2dcf15949da16ad28d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic3f28aa77fc84cb8e2fe43bac7ede253;


Ic3da32f100a43f826b89a492544e7812 Ia2558b16ffc0016f3be46086e0114716 (
.flogtanh_sel( I90bd9107f4c931fa1ccb92998ea8cdeb[flogtanh_SEL-1:0]),
.flogtanh( I7f91c0e606b4082c6aec2e1f111079c5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9574759e112f27778f3645d5d49126b7 = (I90bd9107f4c931fa1ccb92998ea8cdeb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7f91c0e606b4082c6aec2e1f111079c5;


Ic3da32f100a43f826b89a492544e7812 I2c434ceb259b89d6ebfa3631a6e61a05 (
.flogtanh_sel( Ida1c729e6bfcec2c31a92aa9002f2c68[flogtanh_SEL-1:0]),
.flogtanh( I8e0d66c2112193437146e0f503623559),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2ffb7c2ad09bac694ef13ec41e5de327 = (Ida1c729e6bfcec2c31a92aa9002f2c68[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8e0d66c2112193437146e0f503623559;


Ic3da32f100a43f826b89a492544e7812 I3f5ebedbc02e16f3f3d92630e0f7f5ab (
.flogtanh_sel( Ib848feeccd0ea78ebc8ba8368534c3d1[flogtanh_SEL-1:0]),
.flogtanh( Iabe6bf045784762fb6b97be3587fd68d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib190f589f4d663dbc0a3c166a8dcf5fa = (Ib848feeccd0ea78ebc8ba8368534c3d1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iabe6bf045784762fb6b97be3587fd68d;


Ic3da32f100a43f826b89a492544e7812 I99149a651e7e1b07163d0d9d8412ac07 (
.flogtanh_sel( Icc11970bbae3adcfa33a0e5dba3e78f4[flogtanh_SEL-1:0]),
.flogtanh( I11f0fd7033065e1695d846f08d11aed5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I459c59ac61179d74170db53bf45ba89e = (Icc11970bbae3adcfa33a0e5dba3e78f4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I11f0fd7033065e1695d846f08d11aed5;


Ic3da32f100a43f826b89a492544e7812 I2a494d1be114bbdc4dba4baf5f2b509f (
.flogtanh_sel( I86bb4ef4bdd7af8861280ef30fbeeeea[flogtanh_SEL-1:0]),
.flogtanh( Ife1589d99f0764e3757de2a7d8b43008),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie5e432a991aff25577639f1b4ffd594f = (I86bb4ef4bdd7af8861280ef30fbeeeea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ife1589d99f0764e3757de2a7d8b43008;


Ic3da32f100a43f826b89a492544e7812 I0d2a2da6a5771ddd912fd021ece83287 (
.flogtanh_sel( I7e0c259c6c7bacdff5edc44a22e005ba[flogtanh_SEL-1:0]),
.flogtanh( I7cb3f1f2e7f997b861d6c63d55c0f4ca),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I72064a6a84ff956d76a5aa590bbc05a9 = (I7e0c259c6c7bacdff5edc44a22e005ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7cb3f1f2e7f997b861d6c63d55c0f4ca;


Ic3da32f100a43f826b89a492544e7812 I913a65b376473b5c7dae5ba5363fdb5f (
.flogtanh_sel( I897ddba059b27f7ed009b0cb70cfb46f[flogtanh_SEL-1:0]),
.flogtanh( Iae2f185d6338026f3e37696327f214df),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iea74ecbac92e1b8f2ec7ad68d10b8e7d = (I897ddba059b27f7ed009b0cb70cfb46f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iae2f185d6338026f3e37696327f214df;


Ic3da32f100a43f826b89a492544e7812 I9a768e529d163e801f0a14696252c762 (
.flogtanh_sel( I4496243eb0542a514b551b4d09bffd7d[flogtanh_SEL-1:0]),
.flogtanh( I4da8f5b31f5cf7c70bba0cf661d727d8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4f72d0db9fcc358c6fbec9964fbe0bbb = (I4496243eb0542a514b551b4d09bffd7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4da8f5b31f5cf7c70bba0cf661d727d8;


Ic3da32f100a43f826b89a492544e7812 Iaa838d18ba96363e9ec0d600b4dda588 (
.flogtanh_sel( Ic931fb08b2e8441321ebdeed84576a0d[flogtanh_SEL-1:0]),
.flogtanh( I46dd3a6d37d3df901689403a6215b65d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifd958901d2ea2284f506e04a058012fa = (Ic931fb08b2e8441321ebdeed84576a0d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I46dd3a6d37d3df901689403a6215b65d;


Ic3da32f100a43f826b89a492544e7812 I671d9c208058c949f51a066e723dfcd3 (
.flogtanh_sel( Ieb6af5390b98e893ee05a939c16d2ffd[flogtanh_SEL-1:0]),
.flogtanh( I84f43bb1814bdd83a682f7a859cfd611),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie317bbd70b9092b840c0f2713204fb9d = (Ieb6af5390b98e893ee05a939c16d2ffd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I84f43bb1814bdd83a682f7a859cfd611;


Ic3da32f100a43f826b89a492544e7812 I5869a1a085c8e01a2ec070f00f217e66 (
.flogtanh_sel( Ic2a54bad4c5a8885dd24b8687c6db0de[flogtanh_SEL-1:0]),
.flogtanh( I476ea921894e07d3f1d2ff3e7c3b660a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2f9e56d570e72714a06c59aa9e4334c0 = (Ic2a54bad4c5a8885dd24b8687c6db0de[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I476ea921894e07d3f1d2ff3e7c3b660a;


Ic3da32f100a43f826b89a492544e7812 I0b4ce0efef50e77c6bc1452e17257cf1 (
.flogtanh_sel( I6ecbad763d2b48b78a0584beaefc78ee[flogtanh_SEL-1:0]),
.flogtanh( I5cc52764eb8a9961469e1892559ed7ee),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5b53fd45210b92703cb10d583f471ab9 = (I6ecbad763d2b48b78a0584beaefc78ee[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5cc52764eb8a9961469e1892559ed7ee;


Ic3da32f100a43f826b89a492544e7812 I8d0240daf3824abc0b90ac33041d259d (
.flogtanh_sel( I20556d23c873c71c7ebc8a961bf40251[flogtanh_SEL-1:0]),
.flogtanh( I76f68c50b69a7545c0077f5333bfa3e2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8edbe77bacf1975e014faeee6b861980 = (I20556d23c873c71c7ebc8a961bf40251[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I76f68c50b69a7545c0077f5333bfa3e2;


Ic3da32f100a43f826b89a492544e7812 I2cd28720644f1e5529cb04e89d508b53 (
.flogtanh_sel( I79012e6351e6320c22437aa216ea4df1[flogtanh_SEL-1:0]),
.flogtanh( Id0bd4407ef72994435b3794096636553),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I174fcbc2ee01fc55edbc8238e5da7f0c = (I79012e6351e6320c22437aa216ea4df1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id0bd4407ef72994435b3794096636553;


Ic3da32f100a43f826b89a492544e7812 I16b7ce8eacb77c7baa6bfe777b9985d4 (
.flogtanh_sel( Ibf74ab9af877d27c3a6f3881f00ddaf1[flogtanh_SEL-1:0]),
.flogtanh( I0879a96ba0ef5eb523ae807c40c66a63),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id4dc304aef5f35f6ceb91796c278e716 = (Ibf74ab9af877d27c3a6f3881f00ddaf1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0879a96ba0ef5eb523ae807c40c66a63;


Ic3da32f100a43f826b89a492544e7812 I0d4d308354c1ab110438b3ee672b80e5 (
.flogtanh_sel( I843d35db35d7b42a87ce78d3772cec2f[flogtanh_SEL-1:0]),
.flogtanh( I8304ab4dc851d69a7ad7db75ced3eb9e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0cbdfae6f75a639eb591d9c0022f5838 = (I843d35db35d7b42a87ce78d3772cec2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8304ab4dc851d69a7ad7db75ced3eb9e;


Ic3da32f100a43f826b89a492544e7812 I40ade6ae3e353967c3cb23faa09014e2 (
.flogtanh_sel( I2b1398b4bfd374d7221b0a68da28e979[flogtanh_SEL-1:0]),
.flogtanh( I24d773b608ba1ee21855540ee84028da),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I088898ee932a96c14f2f0f568f5455b6 = (I2b1398b4bfd374d7221b0a68da28e979[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I24d773b608ba1ee21855540ee84028da;


Ic3da32f100a43f826b89a492544e7812 I0376f7a762e8efd708830d38a64dce26 (
.flogtanh_sel( I6f615d6e74b0c02f8e4265523ad16404[flogtanh_SEL-1:0]),
.flogtanh( I9458b9a213600ce0c8c1d54d31c8c5c2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ide0abde3644a4fafb436aa59768d016e = (I6f615d6e74b0c02f8e4265523ad16404[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9458b9a213600ce0c8c1d54d31c8c5c2;


Ic3da32f100a43f826b89a492544e7812 Ie232b3917a3ad670e0c8bf8c443327c6 (
.flogtanh_sel( Iae8a98dd4a7cbfbc56c1404b6a2020af[flogtanh_SEL-1:0]),
.flogtanh( Idb6b8e6f2df9b8d96efa93830df86a71),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I08581dc8d42be712cfb36d744f2786e0 = (Iae8a98dd4a7cbfbc56c1404b6a2020af[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idb6b8e6f2df9b8d96efa93830df86a71;


Ic3da32f100a43f826b89a492544e7812 I0b78dbb4e8047b32554e7602dd446e4e (
.flogtanh_sel( Iad53375a54d01c559c74981bf279dfb5[flogtanh_SEL-1:0]),
.flogtanh( I0a8fb8a7a28b364bc8cf49b96fdc66a4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I29fb3830a5fc5922f1ec687a38941e97 = (Iad53375a54d01c559c74981bf279dfb5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0a8fb8a7a28b364bc8cf49b96fdc66a4;


Ic3da32f100a43f826b89a492544e7812 I2d5b32b0396ccf16f181dac6de312612 (
.flogtanh_sel( I5db1307f922e0c742d7d9f3a79a4a4f3[flogtanh_SEL-1:0]),
.flogtanh( I938f8896ddbf95751aea2b327f5d40f0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I715d59fb27e519a9b76bdd8b5139a619 = (I5db1307f922e0c742d7d9f3a79a4a4f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I938f8896ddbf95751aea2b327f5d40f0;


Ic3da32f100a43f826b89a492544e7812 Ifba9b8b58b0cc72cc74bd41051b9a77b (
.flogtanh_sel( I9f78172ed5bf73752196f9a8810005f3[flogtanh_SEL-1:0]),
.flogtanh( Ib5b964583d3ef33b47643ca212bc0ada),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibe6a876a041198a581c95457a7d1fcf8 = (I9f78172ed5bf73752196f9a8810005f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib5b964583d3ef33b47643ca212bc0ada;


Ic3da32f100a43f826b89a492544e7812 I3e4e7e8ebe409db10c9bd3830b1bc05c (
.flogtanh_sel( If85a22d670d47f491dd7568d0453ba1d[flogtanh_SEL-1:0]),
.flogtanh( I4bae2a264af742ffe7be73f9a1129efe),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iec078a95a69b081cfb5e987ba9c5a613 = (If85a22d670d47f491dd7568d0453ba1d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4bae2a264af742ffe7be73f9a1129efe;


Ic3da32f100a43f826b89a492544e7812 I873553498a2422d54b3265dacc59d21b (
.flogtanh_sel( Ib9e529170b2896e930a839295796fd31[flogtanh_SEL-1:0]),
.flogtanh( I041c1a7ef6128c7a1a8f8593d4401f1b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0e8f3f56bce3be1ee4d5f780a2f2a9fe = (Ib9e529170b2896e930a839295796fd31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I041c1a7ef6128c7a1a8f8593d4401f1b;


Ic3da32f100a43f826b89a492544e7812 Iff42f3f1b188bddfbe4d1767f884b694 (
.flogtanh_sel( Ib7af536846bac40c1f221d1f72c6c25c[flogtanh_SEL-1:0]),
.flogtanh( I22c6d2c87ef183ef45805a7c99a7e473),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia73cacadbf80c0701a5b5b430c0d5c98 = (Ib7af536846bac40c1f221d1f72c6c25c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I22c6d2c87ef183ef45805a7c99a7e473;


Ic3da32f100a43f826b89a492544e7812 I342479741035bb20f2751eabb645b1a3 (
.flogtanh_sel( Ib0eb61a2cb831dd35ce9850994e7c2da[flogtanh_SEL-1:0]),
.flogtanh( I45fef5261954fc84be265f39eb8f9647),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic634d26fc09589a29a160e4efb5613a8 = (Ib0eb61a2cb831dd35ce9850994e7c2da[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I45fef5261954fc84be265f39eb8f9647;


Ic3da32f100a43f826b89a492544e7812 Icd8e0b5b7b99f5bef0f6e7ef36f9d383 (
.flogtanh_sel( I89d338f59960af7a47595d6afa206abc[flogtanh_SEL-1:0]),
.flogtanh( I3b292cf842e3a7ca9e6d0c4ab345446f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie1374cac341cf353b1863dae9f544e8b = (I89d338f59960af7a47595d6afa206abc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3b292cf842e3a7ca9e6d0c4ab345446f;


Ic3da32f100a43f826b89a492544e7812 I7dc03977d6d0cb6123ddd123dcf76338 (
.flogtanh_sel( Ib3c1176eb8991e3e85855a9fe845c303[flogtanh_SEL-1:0]),
.flogtanh( Ie7bff678d39738eb49b599772586210a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia07447985347e9a7f3739bd98867cdfb = (Ib3c1176eb8991e3e85855a9fe845c303[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie7bff678d39738eb49b599772586210a;


Ic3da32f100a43f826b89a492544e7812 Ifbabcd4c164db768beed91f6203e590b (
.flogtanh_sel( I93073d05d509b821a743998cf32c58ee[flogtanh_SEL-1:0]),
.flogtanh( Ib9d80aab3818d682b54122974fa3a424),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2121318f589878b4a9260625f97de518 = (I93073d05d509b821a743998cf32c58ee[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib9d80aab3818d682b54122974fa3a424;


Ic3da32f100a43f826b89a492544e7812 I693deabd302d69a1bca4216b0172b7ef (
.flogtanh_sel( Iab6dac1909c1564c3890ffecc13418df[flogtanh_SEL-1:0]),
.flogtanh( Iaa05186a94ba0559ab57ced9202ccefb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibd8424c228f87f85df3da6204edff2b5 = (Iab6dac1909c1564c3890ffecc13418df[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaa05186a94ba0559ab57ced9202ccefb;


Ic3da32f100a43f826b89a492544e7812 Iecd6b9565c414d2ebe2253ac59dac257 (
.flogtanh_sel( I1b75eeb29167a171d89f6e67039436d5[flogtanh_SEL-1:0]),
.flogtanh( I506f39735c3743b3705980c73295c035),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8a7fb51566bf215af214cd2fb5209974 = (I1b75eeb29167a171d89f6e67039436d5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I506f39735c3743b3705980c73295c035;


Ic3da32f100a43f826b89a492544e7812 Ided860652e11465175045394b3dc2968 (
.flogtanh_sel( I3a31adc52a1405555017b2ddf219b407[flogtanh_SEL-1:0]),
.flogtanh( I8f16ead6735608b15b364b9af9b3a22a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7c0f872988488ac69815d288885dfd2f = (I3a31adc52a1405555017b2ddf219b407[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8f16ead6735608b15b364b9af9b3a22a;


Ic3da32f100a43f826b89a492544e7812 I8e9a30125869fa8591b0140843744e39 (
.flogtanh_sel( Iaadba89c6a370240fc0758029f7d8db0[flogtanh_SEL-1:0]),
.flogtanh( Id07af023803badc88c51b891cad1b7e5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3521b10b97b0e74888ce385cfc772945 = (Iaadba89c6a370240fc0758029f7d8db0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id07af023803badc88c51b891cad1b7e5;


Ic3da32f100a43f826b89a492544e7812 I140f82b37ecf788cfb0e8b5f8b2b1f10 (
.flogtanh_sel( I4f4a64fb3ced7d9f7ee4513178e9655a[flogtanh_SEL-1:0]),
.flogtanh( Iecb522fa10764b2c0c044be6c1ca807d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I58f0b81a46549cab8e74ecbc285df23a = (I4f4a64fb3ced7d9f7ee4513178e9655a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iecb522fa10764b2c0c044be6c1ca807d;


Ic3da32f100a43f826b89a492544e7812 Ifc01a716b72e1be7c9c752becef15cd7 (
.flogtanh_sel( I0c76ca58f69c91758e755cd581241284[flogtanh_SEL-1:0]),
.flogtanh( I58b9a09be96353ba6c18f310e1987742),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7095040b38bf9d6b5229c11d2a0d7c57 = (I0c76ca58f69c91758e755cd581241284[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I58b9a09be96353ba6c18f310e1987742;


Ic3da32f100a43f826b89a492544e7812 I6b591e575b56dba4bf43107c5b498a9d (
.flogtanh_sel( I2312bce18958346149c868846e04643b[flogtanh_SEL-1:0]),
.flogtanh( I86ced95bff4327e4ab07338663f82029),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I675ab6c4fb93b006f3fcafc985fbc405 = (I2312bce18958346149c868846e04643b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I86ced95bff4327e4ab07338663f82029;


Ic3da32f100a43f826b89a492544e7812 I24f2539727ade2e7e37c94d1544aced2 (
.flogtanh_sel( I3e154098cb0a48f1c23234f46613f406[flogtanh_SEL-1:0]),
.flogtanh( Ia802328754db2d72d6ec8e12a79b2341),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I239a992ebb62899120a74b1c9e6cc4b4 = (I3e154098cb0a48f1c23234f46613f406[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia802328754db2d72d6ec8e12a79b2341;


Ic3da32f100a43f826b89a492544e7812 I93fd9f3656565455fafd170b68223409 (
.flogtanh_sel( I1645c1c588bcbf15dd62d47e08b8e139[flogtanh_SEL-1:0]),
.flogtanh( I5b5a9fa50a6e4c7e07017249e5dee137),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I927c870d09285dcb47e6d399f319471e = (I1645c1c588bcbf15dd62d47e08b8e139[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5b5a9fa50a6e4c7e07017249e5dee137;


Ic3da32f100a43f826b89a492544e7812 I69b5ca5e88e19dd32779cb7935f5f86f (
.flogtanh_sel( I4c25de66590e1745d37112e08d8c8e2c[flogtanh_SEL-1:0]),
.flogtanh( I73ef262450353dfcfabe3051ab0006f9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie23ed3ee61f468f59f2baf661cb7f85d = (I4c25de66590e1745d37112e08d8c8e2c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I73ef262450353dfcfabe3051ab0006f9;


Ic3da32f100a43f826b89a492544e7812 I18ef26b96443ee652955845b9caaf007 (
.flogtanh_sel( Ia03092ac621b8dd1c206fea1e8b0215f[flogtanh_SEL-1:0]),
.flogtanh( I959c5d62629333d1d60766a6d935ae4a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I68e58664be09261e5a80d6f8ecdd1b60 = (Ia03092ac621b8dd1c206fea1e8b0215f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I959c5d62629333d1d60766a6d935ae4a;


Ic3da32f100a43f826b89a492544e7812 I35a35f4e0d7f5fc1bb8fb8cc1008d939 (
.flogtanh_sel( I5c9bdb033436dc9f6069baca31f24c2d[flogtanh_SEL-1:0]),
.flogtanh( I659d579ea5b5d24ef0ccbb8160dfe2ae),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id2808e0f40992c79ead4da7c734e5b79 = (I5c9bdb033436dc9f6069baca31f24c2d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I659d579ea5b5d24ef0ccbb8160dfe2ae;


Ic3da32f100a43f826b89a492544e7812 Ic1a6258e1cb28cc62901bfd08f870891 (
.flogtanh_sel( I8f07cf4865480f18ad6945974ec2231c[flogtanh_SEL-1:0]),
.flogtanh( Icae3ba8a84ee6ee051a3caf210f47b51),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icb2b390266bff241a688961136db0f51 = (I8f07cf4865480f18ad6945974ec2231c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icae3ba8a84ee6ee051a3caf210f47b51;


Ic3da32f100a43f826b89a492544e7812 I17a1a725957eb14db657229438e010be (
.flogtanh_sel( I4a7119e8862fe4a6a4100dd9ac67dd24[flogtanh_SEL-1:0]),
.flogtanh( I92a005abe2d27beb2949fe29c0d8bc65),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I54cfd68212d97a2cc8241ef429429453 = (I4a7119e8862fe4a6a4100dd9ac67dd24[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I92a005abe2d27beb2949fe29c0d8bc65;


Ic3da32f100a43f826b89a492544e7812 I1cace2c01ed0dc98e0c2023d1bd1e40d (
.flogtanh_sel( Id78fcfc6724a05f46d44d7c3e7d0c756[flogtanh_SEL-1:0]),
.flogtanh( I28fb1164936618d653aa7bf06c03b38f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8d4e3962525c424786ae822a6981a5e6 = (Id78fcfc6724a05f46d44d7c3e7d0c756[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I28fb1164936618d653aa7bf06c03b38f;


Ic3da32f100a43f826b89a492544e7812 I5d881507a603040f0a52c38593fdc025 (
.flogtanh_sel( I7cbd9d619623cbabf8ed6b1fece8f012[flogtanh_SEL-1:0]),
.flogtanh( I8720bdf2c91f113b39aa5b6f82421feb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1a5f22b4e326d1684c0a8c7a7e754ab4 = (I7cbd9d619623cbabf8ed6b1fece8f012[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8720bdf2c91f113b39aa5b6f82421feb;


Ic3da32f100a43f826b89a492544e7812 Id78b9db28e07ea13fb557951fc97e5e1 (
.flogtanh_sel( I58951165d251e370b0f3b3fb537aed18[flogtanh_SEL-1:0]),
.flogtanh( I07320e5fb3beddb93ae325a98c5e3782),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8c2e0c83a8204d6b21e0e3e458d56f05 = (I58951165d251e370b0f3b3fb537aed18[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I07320e5fb3beddb93ae325a98c5e3782;


Ic3da32f100a43f826b89a492544e7812 I8cf7cf89ca1b68dc37dbd3578061e2d7 (
.flogtanh_sel( I21daac106f526d84cb8fa5239c19499d[flogtanh_SEL-1:0]),
.flogtanh( Ib8b29bc86ad9c07d7ae5b358f66cb9ba),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie0622ff815747e4a9f368c74787026ec = (I21daac106f526d84cb8fa5239c19499d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib8b29bc86ad9c07d7ae5b358f66cb9ba;


Ic3da32f100a43f826b89a492544e7812 I037169c21915407665840871e00e4e5e (
.flogtanh_sel( I178029cec3a5d6141abdfa91b91fdbf4[flogtanh_SEL-1:0]),
.flogtanh( I8e2ed2040f5bf8ea125e5b953cf89300),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5ffed139764d90825b9f2eddacd0eddc = (I178029cec3a5d6141abdfa91b91fdbf4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8e2ed2040f5bf8ea125e5b953cf89300;


Ic3da32f100a43f826b89a492544e7812 I2bbccb53115e379bbaba76acd24bda1f (
.flogtanh_sel( I96dfb2efbb55a644616e3474ed07c364[flogtanh_SEL-1:0]),
.flogtanh( I4ad3a5b591cd6b13de04897fbbd068ec),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5a3297f48e1045273db6522744582b05 = (I96dfb2efbb55a644616e3474ed07c364[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4ad3a5b591cd6b13de04897fbbd068ec;


Ic3da32f100a43f826b89a492544e7812 I50a053c0231be5a1634602c4794dfc69 (
.flogtanh_sel( I7a17d8f0e2d16c441044db68ee037731[flogtanh_SEL-1:0]),
.flogtanh( If5208f94e99b0e7ff353c048b55ad7ba),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9858bb2a3cc458aca5bf7eb077ee55dd = (I7a17d8f0e2d16c441044db68ee037731[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If5208f94e99b0e7ff353c048b55ad7ba;


Ic3da32f100a43f826b89a492544e7812 I8403de216283749679bd1d87db013c9f (
.flogtanh_sel( I2ced9bb3ae6bdc5b5ef2865fb46abf07[flogtanh_SEL-1:0]),
.flogtanh( I66106fad536bb49418e7d09e3f4221ac),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6e7e27bb176196e4493bf9c45ca19719 = (I2ced9bb3ae6bdc5b5ef2865fb46abf07[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I66106fad536bb49418e7d09e3f4221ac;


Ic3da32f100a43f826b89a492544e7812 I445dbab6081152c2547362d6edda0f9d (
.flogtanh_sel( I89a93384020d93cf4d26b3902e06cd9e[flogtanh_SEL-1:0]),
.flogtanh( I6af88c096ca3af849bbedb15b2ac7153),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4cff1804df738cbf4f940c775236df9c = (I89a93384020d93cf4d26b3902e06cd9e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6af88c096ca3af849bbedb15b2ac7153;


Ic3da32f100a43f826b89a492544e7812 I664c35dbfcf6d39b6b76c6070c7a740f (
.flogtanh_sel( Ibbb47d29b9a45559c13ffa3b046c66f5[flogtanh_SEL-1:0]),
.flogtanh( I15d6e1e431457b954b5f86cd4fb16a77),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0c1e22375d5e023c24519901b92eceb5 = (Ibbb47d29b9a45559c13ffa3b046c66f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I15d6e1e431457b954b5f86cd4fb16a77;


Ic3da32f100a43f826b89a492544e7812 I336a4543ebe1b9014e0a3422d93939ce (
.flogtanh_sel( I0034177eb1049577a3578b371527f34b[flogtanh_SEL-1:0]),
.flogtanh( Ifd67d6dec292171610a805560d7cb9a0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ida5b16851dc06534844a0b037d74feb3 = (I0034177eb1049577a3578b371527f34b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifd67d6dec292171610a805560d7cb9a0;


Ic3da32f100a43f826b89a492544e7812 Ibb6ecd70a6ef7e136ba0656a1e13795f (
.flogtanh_sel( I22d9ea7bb5a1a3405bcd04b9af40fa62[flogtanh_SEL-1:0]),
.flogtanh( I681c4ec303ff366746d35234fe5a1ff4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iac3cb5b4481687fcf430c8bf52cfb74d = (I22d9ea7bb5a1a3405bcd04b9af40fa62[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I681c4ec303ff366746d35234fe5a1ff4;


Ic3da32f100a43f826b89a492544e7812 I66446889f5308ddf7fcfa1c51cb11b2a (
.flogtanh_sel( I8a632e7a911bf5726fee587189cb6f16[flogtanh_SEL-1:0]),
.flogtanh( I5df2eac3ace0bcef9e48b0850d975cce),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia1499972c4995268acd828c1289f353d = (I8a632e7a911bf5726fee587189cb6f16[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5df2eac3ace0bcef9e48b0850d975cce;


Ic3da32f100a43f826b89a492544e7812 I51b1fb49194b03138c35f709755a229f (
.flogtanh_sel( I3765afc490b34e8a310998a4ebcff8cb[flogtanh_SEL-1:0]),
.flogtanh( Icf6f5254160a82036c4ba0367e8f0404),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie559401a3a913400dc5e3e5641297fa6 = (I3765afc490b34e8a310998a4ebcff8cb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icf6f5254160a82036c4ba0367e8f0404;


Ic3da32f100a43f826b89a492544e7812 Ie36d9c4c51fcd919dabd8762784eab27 (
.flogtanh_sel( I7607e800ae46a96e016b303120da4247[flogtanh_SEL-1:0]),
.flogtanh( If1de12bbb90e49cc1b28eafc2aa551e5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie0667fbe76244eaec0b155d69dcc9447 = (I7607e800ae46a96e016b303120da4247[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If1de12bbb90e49cc1b28eafc2aa551e5;


Ic3da32f100a43f826b89a492544e7812 Id1d58ca8250befaf9188d985d342eed4 (
.flogtanh_sel( I29b2f1fddee5e32f217d25410bcfce4f[flogtanh_SEL-1:0]),
.flogtanh( Ibf9f7f1f6a759af21ac82d6e6ff7df43),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1d0f031e8ae9c0335d501d1565118220 = (I29b2f1fddee5e32f217d25410bcfce4f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibf9f7f1f6a759af21ac82d6e6ff7df43;


Ic3da32f100a43f826b89a492544e7812 I923303497e7d4bad25127787f325d38e (
.flogtanh_sel( Iba5f8a31a81f6aa06f5e38c03dc6db54[flogtanh_SEL-1:0]),
.flogtanh( Ie44bc9632854c4c2077bcec5f46d29ad),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie2c801b2de066c3218d7312615b7bfda = (Iba5f8a31a81f6aa06f5e38c03dc6db54[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie44bc9632854c4c2077bcec5f46d29ad;


Ic3da32f100a43f826b89a492544e7812 Icd41893ab6ca9a98a6a074b94031b531 (
.flogtanh_sel( Ifcb5c907ad503331317599e4e0ce7be8[flogtanh_SEL-1:0]),
.flogtanh( I97ae894cd928e17cad4c4631aec2c7a0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I64c4bb0d40d80ec52aab61ce46954f43 = (Ifcb5c907ad503331317599e4e0ce7be8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I97ae894cd928e17cad4c4631aec2c7a0;


Ic3da32f100a43f826b89a492544e7812 Id3564b6edcf9a0f7774eadcf5bb1a351 (
.flogtanh_sel( I62d6f2ab4ec8b6ecfa544ad4d90eb30b[flogtanh_SEL-1:0]),
.flogtanh( I500a903104b4b532b3c07d1640e80b55),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I512f57a40c7c8cb2f040bdde73e44ca3 = (I62d6f2ab4ec8b6ecfa544ad4d90eb30b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I500a903104b4b532b3c07d1640e80b55;


Ic3da32f100a43f826b89a492544e7812 I612477e72ad9148a39f41bbbc9e66388 (
.flogtanh_sel( Ide65414c51b3cb182c0f2f238903d60a[flogtanh_SEL-1:0]),
.flogtanh( I1d3ae54c8fa3d87a39e3a51018a20727),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id60cbf534604e5dba988050ef5abe625 = (Ide65414c51b3cb182c0f2f238903d60a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1d3ae54c8fa3d87a39e3a51018a20727;


Ic3da32f100a43f826b89a492544e7812 If3b251847164b3a628df40b0cc0fb0bf (
.flogtanh_sel( I03a8dc2288eaeb619e746990e20cc868[flogtanh_SEL-1:0]),
.flogtanh( I23d3b6da58b66185ddb3c5eae0f68dae),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I37998a91d20db2248ebdd8e661d42f70 = (I03a8dc2288eaeb619e746990e20cc868[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I23d3b6da58b66185ddb3c5eae0f68dae;


Ic3da32f100a43f826b89a492544e7812 I259bfae820c96dc73e3aeebcf07abc30 (
.flogtanh_sel( Id81c1b44d16ddbcd466382c60fe84986[flogtanh_SEL-1:0]),
.flogtanh( I88b1352db9aa35be019bc0f345c7131e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib65ff82aff398f6ff7ba711a36f41ee4 = (Id81c1b44d16ddbcd466382c60fe84986[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I88b1352db9aa35be019bc0f345c7131e;


Ic3da32f100a43f826b89a492544e7812 I381aa14f5aa2bf8501fbf80bee931cc5 (
.flogtanh_sel( I503d72f4a2fd20dbf35aa27321d2ede7[flogtanh_SEL-1:0]),
.flogtanh( I1115071c073981f4db4917844fb12a73),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3d1dd8b9c7c6d3913f7ac369ad7e625c = (I503d72f4a2fd20dbf35aa27321d2ede7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1115071c073981f4db4917844fb12a73;


Ic3da32f100a43f826b89a492544e7812 Ib2df341e0d57303f2090d58b2c003043 (
.flogtanh_sel( Id6595a4cf33062d1f05cbcee2d0685f1[flogtanh_SEL-1:0]),
.flogtanh( Ia9e4e593fd82657c81aeea8fbcd1194b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I097722547450582dc5776bdaff914741 = (Id6595a4cf33062d1f05cbcee2d0685f1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia9e4e593fd82657c81aeea8fbcd1194b;


Ic3da32f100a43f826b89a492544e7812 Ie608e1662710e3bf50e77976d124d5a2 (
.flogtanh_sel( I83ebdd7331ca8fbcf5250851b346c0b0[flogtanh_SEL-1:0]),
.flogtanh( I22300986ed621a97a6dac1f3b4d59b8e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id4a213e494f9c9be0fd1a307e87c756a = (I83ebdd7331ca8fbcf5250851b346c0b0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I22300986ed621a97a6dac1f3b4d59b8e;


Ic3da32f100a43f826b89a492544e7812 Ifa74b9ea0dc984201251de4556d1914c (
.flogtanh_sel( I7f6ea26cdfe5986065e7b5aa6842cc1c[flogtanh_SEL-1:0]),
.flogtanh( Icc08ab7c64b40e53278a93f4ae0f9209),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I21594c8b0169efd7c2aa6cbc31f4a901 = (I7f6ea26cdfe5986065e7b5aa6842cc1c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icc08ab7c64b40e53278a93f4ae0f9209;


Ic3da32f100a43f826b89a492544e7812 I953a8f5d42f964efd7360912c7108300 (
.flogtanh_sel( Idab1ec32c20f93c4cc1acb38158f92d5[flogtanh_SEL-1:0]),
.flogtanh( I8cc9f5531f2675b3058df110912551b6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I15022e1b349eee259d3567837283dbf6 = (Idab1ec32c20f93c4cc1acb38158f92d5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8cc9f5531f2675b3058df110912551b6;


Ic3da32f100a43f826b89a492544e7812 I2416bd8b90c2f46a7b265b18c6f4c12f (
.flogtanh_sel( I0738add83419502e73674ded2f1ad6c7[flogtanh_SEL-1:0]),
.flogtanh( Icdba6332ba9ea91ffefd690150fba09f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1070940dc2ef6e8ee3d1227ec9ff3162 = (I0738add83419502e73674ded2f1ad6c7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icdba6332ba9ea91ffefd690150fba09f;


Ic3da32f100a43f826b89a492544e7812 I9b821269f3d41a016ed696f17d34b1bd (
.flogtanh_sel( I6c93e63a8e5a2dbd598f1565c7323b39[flogtanh_SEL-1:0]),
.flogtanh( Idaef789d04cd5c6291dae88f616460e6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8922cc37cde6ba132f632743113e42af = (I6c93e63a8e5a2dbd598f1565c7323b39[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idaef789d04cd5c6291dae88f616460e6;


Ic3da32f100a43f826b89a492544e7812 Icbaf905be551871493ffac5a7daacc0e (
.flogtanh_sel( I4aa57a9d46371f1680d5f95596f60b5d[flogtanh_SEL-1:0]),
.flogtanh( I016cb9c8307b28a7cabf9a91e8da03d6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia66c399023e500ed67197dcf236f5d42 = (I4aa57a9d46371f1680d5f95596f60b5d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I016cb9c8307b28a7cabf9a91e8da03d6;


Ic3da32f100a43f826b89a492544e7812 I56d0d1fe5a3d0bd8c5534139cafb2954 (
.flogtanh_sel( I5369a7203b78951a3c006c2d3b22507c[flogtanh_SEL-1:0]),
.flogtanh( I54517f62dd6f2e7de7d522dfc506383e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1171dc208d5db1024dc3f09a90c78ca0 = (I5369a7203b78951a3c006c2d3b22507c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I54517f62dd6f2e7de7d522dfc506383e;


Ic3da32f100a43f826b89a492544e7812 I32977d796f3fb2c52e4bd90f1daf35a5 (
.flogtanh_sel( Ie72a79a6966cf198687b7c8a8bcdeb13[flogtanh_SEL-1:0]),
.flogtanh( I6b0c1ef6f0a94adaf62425829edf28dd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic28b148967a5b3d05409976fa9001ac8 = (Ie72a79a6966cf198687b7c8a8bcdeb13[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6b0c1ef6f0a94adaf62425829edf28dd;


Ic3da32f100a43f826b89a492544e7812 I1d01b61d41838e56f7a37538f8dc10af (
.flogtanh_sel( Ie917ae4c44ab0f9c2f1747ff0d2a754e[flogtanh_SEL-1:0]),
.flogtanh( I067ce754b1084de762c33b295f2f47b2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I79fe46308b93fbb24245fe1c75edf4a5 = (Ie917ae4c44ab0f9c2f1747ff0d2a754e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I067ce754b1084de762c33b295f2f47b2;


Ic3da32f100a43f826b89a492544e7812 I222d8e31c344ea83aa17b2d4105f8f77 (
.flogtanh_sel( I0b1a31ccb34a742552c11b1945e23dd8[flogtanh_SEL-1:0]),
.flogtanh( Ib2fe88cfe23c363993dfcb7722c4fef0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3bfcd63e92f1949234ab1d2701dbb499 = (I0b1a31ccb34a742552c11b1945e23dd8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib2fe88cfe23c363993dfcb7722c4fef0;


Ic3da32f100a43f826b89a492544e7812 Ie048f388e3db01938d09f49f6a460f4b (
.flogtanh_sel( I9a65a845cf2eced39050e8481665f557[flogtanh_SEL-1:0]),
.flogtanh( I71f836227a1f7f81500a6c980c06f1f7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5e2331edf6e881e9f3a8c47eebda0ac4 = (I9a65a845cf2eced39050e8481665f557[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I71f836227a1f7f81500a6c980c06f1f7;


Ic3da32f100a43f826b89a492544e7812 Ic10cddd3acf48fdb75a352de8320a907 (
.flogtanh_sel( I3b402b35d38a9fde312c89b82297c1a5[flogtanh_SEL-1:0]),
.flogtanh( I6faf34757a61a0b64e61ba059aca33fa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4b66c202450986ef0df05e979cc8bc7f = (I3b402b35d38a9fde312c89b82297c1a5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6faf34757a61a0b64e61ba059aca33fa;


Ic3da32f100a43f826b89a492544e7812 I888c37eb7d1083080b4bf6e88617fced (
.flogtanh_sel( I309fa33562370e339c19e2377e6a6a7a[flogtanh_SEL-1:0]),
.flogtanh( Ib1821b79b79aadf1486fe1e2df2f297c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I737daf208eccf95feb3192897586cdce = (I309fa33562370e339c19e2377e6a6a7a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib1821b79b79aadf1486fe1e2df2f297c;


Ic3da32f100a43f826b89a492544e7812 Ief4101d2dfa58fad383a902976f3eaed (
.flogtanh_sel( I7d06aed81222a030837cad2074c68e19[flogtanh_SEL-1:0]),
.flogtanh( I84daf07d3f3790c691b9192f7e2018c1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I29c8133231cfda17668bbe7b692bdfe2 = (I7d06aed81222a030837cad2074c68e19[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I84daf07d3f3790c691b9192f7e2018c1;


Ic3da32f100a43f826b89a492544e7812 I52c6aa1b039e877d4290df8c20627089 (
.flogtanh_sel( I835cc6af0cd8189035f2441c2e0d3100[flogtanh_SEL-1:0]),
.flogtanh( Ib4b3ed1f9d1dee96a3ec846424412e2f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id9d56f09595e80d66c2ac300f7d1d972 = (I835cc6af0cd8189035f2441c2e0d3100[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib4b3ed1f9d1dee96a3ec846424412e2f;


Ic3da32f100a43f826b89a492544e7812 I75786410afa3d66a24ba0809669b22bf (
.flogtanh_sel( If6f768d12f04087246a0d65de1aef99b[flogtanh_SEL-1:0]),
.flogtanh( Ibe73f00bb6f1494ede2e6f11f5e7d3f8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I97e89a2ee18d2688d7c1a640318a1e0d = (If6f768d12f04087246a0d65de1aef99b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibe73f00bb6f1494ede2e6f11f5e7d3f8;


Ic3da32f100a43f826b89a492544e7812 Ie2ea63b2ecd4e5c1294f6dbd58197511 (
.flogtanh_sel( Ie4b180e1e2cadb865b0eaf6509f99dbb[flogtanh_SEL-1:0]),
.flogtanh( I1542461b996a466d7d3d50bb48ebd690),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ife123bf57fe693dabe6aeaa236c4e058 = (Ie4b180e1e2cadb865b0eaf6509f99dbb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1542461b996a466d7d3d50bb48ebd690;


Ic3da32f100a43f826b89a492544e7812 Id0dd3399358a3205792c76d3a0050b4d (
.flogtanh_sel( Ie329a11fc3f6f59f6f1790612fde3250[flogtanh_SEL-1:0]),
.flogtanh( If97a5a2c523f51c5881496c5dc8ad11e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0c0d844fe3b7d35c1ed6bd7cc4e0dc24 = (Ie329a11fc3f6f59f6f1790612fde3250[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If97a5a2c523f51c5881496c5dc8ad11e;


Ic3da32f100a43f826b89a492544e7812 I10a273eee04903171448f3c3fb799465 (
.flogtanh_sel( Idb7ddbee4076f7bf49177e69f5e4d112[flogtanh_SEL-1:0]),
.flogtanh( Ie19ea558cf2a95ca0c8ae769a809d908),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2d9632ae6a0f3ba44c3da8f56ba3fedf = (Idb7ddbee4076f7bf49177e69f5e4d112[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie19ea558cf2a95ca0c8ae769a809d908;


Ic3da32f100a43f826b89a492544e7812 I9a549a2f5bb9adb242cb0037670c296e (
.flogtanh_sel( I614d66a7dca2d08efdfdc157ca803d5c[flogtanh_SEL-1:0]),
.flogtanh( I6532e6299b8c1fdf7f61b3a44b61c35c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I38cc7b117c0bcd5e3060cd370d710d7e = (I614d66a7dca2d08efdfdc157ca803d5c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6532e6299b8c1fdf7f61b3a44b61c35c;


Ic3da32f100a43f826b89a492544e7812 I76fee3100eb2fb8017468ff03ced2e3b (
.flogtanh_sel( Iea16eb0ab70ebb1bc47ae55e11ced62d[flogtanh_SEL-1:0]),
.flogtanh( Ic7102fb8b5df222fff6151e8794bec3c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I793ddbf6a5d026a57ab72984ca19deac = (Iea16eb0ab70ebb1bc47ae55e11ced62d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic7102fb8b5df222fff6151e8794bec3c;


Ic3da32f100a43f826b89a492544e7812 I00ffce2f0d8f51b004cfe67e14914952 (
.flogtanh_sel( Ifa8db43284d5bbebaed4f72d65cf9f92[flogtanh_SEL-1:0]),
.flogtanh( I1f97ea0e7bf46382824cbffc3e94e9df),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I79458089b042e181e37cc44c06d08681 = (Ifa8db43284d5bbebaed4f72d65cf9f92[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1f97ea0e7bf46382824cbffc3e94e9df;


Ic3da32f100a43f826b89a492544e7812 If37cd2d436809a4da71f11b87ee52c8c (
.flogtanh_sel( I365d9f3e8b2a9890427f07386deeb093[flogtanh_SEL-1:0]),
.flogtanh( I801dfe17655932ad8fe9702cbaad270f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I42460fae0acff25fa2b829e39ddcc4fd = (I365d9f3e8b2a9890427f07386deeb093[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I801dfe17655932ad8fe9702cbaad270f;


Ic3da32f100a43f826b89a492544e7812 Ia7c27f8ea615378bc01b8abb21e6cb45 (
.flogtanh_sel( I466aaa0b6cde2ade1901797b8c11e32c[flogtanh_SEL-1:0]),
.flogtanh( Idbd834f0c907b233a8eff58eaca28863),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id3670a6f05d40ab69624544de92b9c64 = (I466aaa0b6cde2ade1901797b8c11e32c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idbd834f0c907b233a8eff58eaca28863;


Ic3da32f100a43f826b89a492544e7812 Idc8d80e360d1f16f4395231495a54596 (
.flogtanh_sel( I7057e329a65ab240ed6cfa824307af65[flogtanh_SEL-1:0]),
.flogtanh( Ic69e0c34630bde15f4172714bc3d92be),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I81800fb49855a4fd2737faa07ff15d29 = (I7057e329a65ab240ed6cfa824307af65[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic69e0c34630bde15f4172714bc3d92be;


Ic3da32f100a43f826b89a492544e7812 I781ff1146cb02b6b7df07b79e6cac075 (
.flogtanh_sel( I624e50e3457d33d12680eaf8e7c34aa3[flogtanh_SEL-1:0]),
.flogtanh( I465a735c8e94ddbfdbaeb2a7652e481e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibfe325e48511372569e0d98d9c4e70e3 = (I624e50e3457d33d12680eaf8e7c34aa3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I465a735c8e94ddbfdbaeb2a7652e481e;


Ic3da32f100a43f826b89a492544e7812 I26fc142459c21e0ed803186ded96a08d (
.flogtanh_sel( I9f356fd6820c33fdb5baff05a781e192[flogtanh_SEL-1:0]),
.flogtanh( Id1c6a3f52dd7972f47cbd8103ace643f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I326660e98f61bb2ced4c23c7bcc9324a = (I9f356fd6820c33fdb5baff05a781e192[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id1c6a3f52dd7972f47cbd8103ace643f;


Ic3da32f100a43f826b89a492544e7812 I937f12d376dc1726882b2584c8bcbd93 (
.flogtanh_sel( I39b9c7c664fe7017731877d145d55b44[flogtanh_SEL-1:0]),
.flogtanh( I26b9e2d073b20376980662c249bf9d43),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic6fa98631d742b27f252fe7c95caef55 = (I39b9c7c664fe7017731877d145d55b44[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I26b9e2d073b20376980662c249bf9d43;


Ic3da32f100a43f826b89a492544e7812 Id4c953a4b226f9ba8424dd45e5142a61 (
.flogtanh_sel( Ic62ffbb9e58e0d08b0dec24bba1dc6f2[flogtanh_SEL-1:0]),
.flogtanh( Id4cc1b15055941d401ded6ff8b777461),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iab6d0f72579687407e029c630b107f7d = (Ic62ffbb9e58e0d08b0dec24bba1dc6f2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id4cc1b15055941d401ded6ff8b777461;


Ic3da32f100a43f826b89a492544e7812 I4b42f38a25461aecd6a4c343a01d8eb6 (
.flogtanh_sel( I8da2a532288fb817e7dc0cb7b4e3761c[flogtanh_SEL-1:0]),
.flogtanh( I064bd1f4b7fa40b2cae3ea361edf9167),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I19eae741ef89baa1a64c403fb29f14f4 = (I8da2a532288fb817e7dc0cb7b4e3761c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I064bd1f4b7fa40b2cae3ea361edf9167;


Ic3da32f100a43f826b89a492544e7812 I115e7b1ec42d65d6045f89cb45a5222a (
.flogtanh_sel( I6a6e559f5c98f846014e8107fea5a5d9[flogtanh_SEL-1:0]),
.flogtanh( I4b5aadc25b0ed6811a665b33d6c4ae2a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I749b9c345f23aae03c595a2c76126ecb = (I6a6e559f5c98f846014e8107fea5a5d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4b5aadc25b0ed6811a665b33d6c4ae2a;


Ic3da32f100a43f826b89a492544e7812 Ib63f47bf1685620b745ca23bad903f43 (
.flogtanh_sel( Ibef9219f577b1a62dfdd77296fbfb24d[flogtanh_SEL-1:0]),
.flogtanh( Ic883bcc70572a237ba0e3d465337bc59),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idc77c7d5123717fc2596a51d904c6d82 = (Ibef9219f577b1a62dfdd77296fbfb24d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic883bcc70572a237ba0e3d465337bc59;


Ic3da32f100a43f826b89a492544e7812 I60bbb4067a4a56df7f17b07664551caf (
.flogtanh_sel( I52e6688b5bfff75529d18e20b22832ce[flogtanh_SEL-1:0]),
.flogtanh( I7181ab1d663b0cbe30861e29fc3f8532),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I779da979707d9712c1626d6025f97599 = (I52e6688b5bfff75529d18e20b22832ce[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7181ab1d663b0cbe30861e29fc3f8532;


Ic3da32f100a43f826b89a492544e7812 I48a65e645eaf9a7c0ad70056a3395bfd (
.flogtanh_sel( Iff22c49354eefca0ea3c5959c14b782c[flogtanh_SEL-1:0]),
.flogtanh( Id3fbb6d083344684de89d99c040b2100),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I97aede8502e443f98938487a5a5c072c = (Iff22c49354eefca0ea3c5959c14b782c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id3fbb6d083344684de89d99c040b2100;


Ic3da32f100a43f826b89a492544e7812 Ic0867b8887815ddada5f9b588f33e224 (
.flogtanh_sel( Ie5377bbdb4111ed00356d5b7737102f3[flogtanh_SEL-1:0]),
.flogtanh( Iee8d139aa5a8ae046f5019abecdbc3c4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie7820d1a242bc28c19ec32d2c91e47b7 = (Ie5377bbdb4111ed00356d5b7737102f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iee8d139aa5a8ae046f5019abecdbc3c4;


Ic3da32f100a43f826b89a492544e7812 Ic27807394fb38478169390b0ee5f7ecf (
.flogtanh_sel( I55bf0f3379a8c44634b8f0a3d06c049e[flogtanh_SEL-1:0]),
.flogtanh( Idc0bfe36a3a9b3006a04d5dfc31b8107),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I82a14e1ee4723e7d9a13c1f2b8b13691 = (I55bf0f3379a8c44634b8f0a3d06c049e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idc0bfe36a3a9b3006a04d5dfc31b8107;


Ic3da32f100a43f826b89a492544e7812 I096dfe35256cf811f9dd6567507148e5 (
.flogtanh_sel( I9bc9541607f4f6aedb686cdde297bcda[flogtanh_SEL-1:0]),
.flogtanh( Ia2462ec52aaccc97597d1dfc2e33b7e2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I77a94cd9186ca546ca9664942ea3537f = (I9bc9541607f4f6aedb686cdde297bcda[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia2462ec52aaccc97597d1dfc2e33b7e2;


Ic3da32f100a43f826b89a492544e7812 Ie9219c63bbd2b4fc7cab8412da065967 (
.flogtanh_sel( Ia4620554fbb1d81a71a15a846e4be2f5[flogtanh_SEL-1:0]),
.flogtanh( I8048bbe27b49b9d248fee919be6dc977),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3c0ddec25c53c166d30eb78d4518840e = (Ia4620554fbb1d81a71a15a846e4be2f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8048bbe27b49b9d248fee919be6dc977;


Ic3da32f100a43f826b89a492544e7812 I299c813aea4c80a074ac238e6991ddef (
.flogtanh_sel( Ibb31b35388ba8ba2ecf98449308ee67d[flogtanh_SEL-1:0]),
.flogtanh( I838d1cc5e9ca5058c25223ec53d9c34f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I98bbe3b75958f10195dee6460cf2aca6 = (Ibb31b35388ba8ba2ecf98449308ee67d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I838d1cc5e9ca5058c25223ec53d9c34f;


Ic3da32f100a43f826b89a492544e7812 Iadc01acc68bf451895eb7a0963a9a47e (
.flogtanh_sel( Ia20410fb3d56587f89a54c00b943b305[flogtanh_SEL-1:0]),
.flogtanh( Id9e5147e089e6e52ef2a687d76534f16),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If6d436031f68ef587750c5c1dfcfffc2 = (Ia20410fb3d56587f89a54c00b943b305[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id9e5147e089e6e52ef2a687d76534f16;


Ic3da32f100a43f826b89a492544e7812 Ia1bc252746e06f4950ce0dfc564540f0 (
.flogtanh_sel( I9d268f3da12e35b9a4229b7340c0f018[flogtanh_SEL-1:0]),
.flogtanh( Ia043941abbcf10c16f086fe8d61dd456),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I461398638cb8280f1779915298540b00 = (I9d268f3da12e35b9a4229b7340c0f018[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia043941abbcf10c16f086fe8d61dd456;


Ic3da32f100a43f826b89a492544e7812 I7055c77cbcbf7ce4ec695e1f5510a551 (
.flogtanh_sel( I2fce29bd666082eedb2fb3ec8b5ae4dd[flogtanh_SEL-1:0]),
.flogtanh( I625ab32380498dfbf9d3290c2053bf3d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I20c65000bbc10299168af7390776a03c = (I2fce29bd666082eedb2fb3ec8b5ae4dd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I625ab32380498dfbf9d3290c2053bf3d;


Ic3da32f100a43f826b89a492544e7812 I1d1416314ed79dda4691239a19f2195c (
.flogtanh_sel( Ia1e8b61e2579a90f5c88ded11c7322c2[flogtanh_SEL-1:0]),
.flogtanh( I903f7844e55d1cd6969352490c275c8e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia840e19ca36795a50ab1a6e6a1729edb = (Ia1e8b61e2579a90f5c88ded11c7322c2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I903f7844e55d1cd6969352490c275c8e;


Ic3da32f100a43f826b89a492544e7812 Ie83447e6dac9967cb1c08a32e4a89122 (
.flogtanh_sel( I8cf3718ba65b7fed72e3955f190e34d1[flogtanh_SEL-1:0]),
.flogtanh( Ie5951bc919195ba594fe87375ad41269),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7d98d1e5f07fccff5f20eaca6363c700 = (I8cf3718ba65b7fed72e3955f190e34d1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie5951bc919195ba594fe87375ad41269;


Ic3da32f100a43f826b89a492544e7812 I889a7e9ca2e0a8b764172da4b7549bb3 (
.flogtanh_sel( I7e802d300af54d394b4ee041798c0513[flogtanh_SEL-1:0]),
.flogtanh( Ieeed8d4eebc0adea7ee0af6a5dbe045c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I97a75b8625ae2a143cf364790ae77753 = (I7e802d300af54d394b4ee041798c0513[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieeed8d4eebc0adea7ee0af6a5dbe045c;


Ic3da32f100a43f826b89a492544e7812 I50c58df3227a67ff685f2ab4c174c78a (
.flogtanh_sel( Id4fd5a4b97cfa1e176a26f3a823c5516[flogtanh_SEL-1:0]),
.flogtanh( I266cd5f0a56cd5171da8d59df0042d5d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idbea892c8109117f90b453efe8ae25af = (Id4fd5a4b97cfa1e176a26f3a823c5516[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I266cd5f0a56cd5171da8d59df0042d5d;


Ic3da32f100a43f826b89a492544e7812 I4e2205ceebfb931e0cbbe883995f1dbe (
.flogtanh_sel( Icbf8d4e75fc66c05eb49c5075696fb07[flogtanh_SEL-1:0]),
.flogtanh( Ie5a57c603ad520441bc5819c81fb877f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icfc1c6d96a3598af73e99a350c387d72 = (Icbf8d4e75fc66c05eb49c5075696fb07[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie5a57c603ad520441bc5819c81fb877f;


Ic3da32f100a43f826b89a492544e7812 I556bd49f54bed7f02f4fa70fd722d330 (
.flogtanh_sel( I746a7e90adb2f213b75ae12a161aca0d[flogtanh_SEL-1:0]),
.flogtanh( I17ac503f4f952f9e2fcdea3f955cc1a9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I523e9b6f828ec7f166750112f8a3f676 = (I746a7e90adb2f213b75ae12a161aca0d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I17ac503f4f952f9e2fcdea3f955cc1a9;


Ic3da32f100a43f826b89a492544e7812 Ia4885673c36273845149a44316d5f87b (
.flogtanh_sel( Icb1029aaaaed8c698862ea9c5e22132c[flogtanh_SEL-1:0]),
.flogtanh( Id8b704aada09411d5f5153d088c1c613),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I79259217f63b2f6263552c434d0e5c93 = (Icb1029aaaaed8c698862ea9c5e22132c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id8b704aada09411d5f5153d088c1c613;


Ic3da32f100a43f826b89a492544e7812 I8a21b374c9d389b17e1ff59558b63c10 (
.flogtanh_sel( Ib93ea7028c172373b53cdafecae32a67[flogtanh_SEL-1:0]),
.flogtanh( If64a200b2dac7049b77e5b6bb03b9cc3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice6db5ba70d3c7499df6723a2df56bfe = (Ib93ea7028c172373b53cdafecae32a67[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If64a200b2dac7049b77e5b6bb03b9cc3;


Ic3da32f100a43f826b89a492544e7812 I19a127cc43a3d4342102de60c015561b (
.flogtanh_sel( If9628275b000e418f3903daebfdace92[flogtanh_SEL-1:0]),
.flogtanh( Iee1b48cae01fe51344b8d662ace9c6f1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I28aa517220bf597cf898660f698ef19d = (If9628275b000e418f3903daebfdace92[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iee1b48cae01fe51344b8d662ace9c6f1;


Ic3da32f100a43f826b89a492544e7812 If3cd18d66bfb945556f3bac0d778a01f (
.flogtanh_sel( I830202fb6f08f98c7f71893a881bd555[flogtanh_SEL-1:0]),
.flogtanh( Ic879cd355d61eb021250d62841115a52),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I07048dc5cbe24ff72d24902d572face0 = (I830202fb6f08f98c7f71893a881bd555[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic879cd355d61eb021250d62841115a52;


Ic3da32f100a43f826b89a492544e7812 I6637af7e16dac0b96bafb48078493b27 (
.flogtanh_sel( I6f38bc9359562f57c1603355e9ee312b[flogtanh_SEL-1:0]),
.flogtanh( I46e2d889b9ba7eccad5529200852ca17),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iab3876e5107e3a56b1fafe41e16d9482 = (I6f38bc9359562f57c1603355e9ee312b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I46e2d889b9ba7eccad5529200852ca17;


Ic3da32f100a43f826b89a492544e7812 Ia7fc9b93f27f3463bf877f45aaa993f9 (
.flogtanh_sel( I4701b732d59c26e3790a63c1936f9a24[flogtanh_SEL-1:0]),
.flogtanh( Ia4e080f13520998be95b64eb883f8e32),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I511a55c2f4d6d3727dff5825597f55a9 = (I4701b732d59c26e3790a63c1936f9a24[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia4e080f13520998be95b64eb883f8e32;


Ic3da32f100a43f826b89a492544e7812 I506a2555ca7dd87dd64008bb6efb1590 (
.flogtanh_sel( Ib5d28d8f73d17ab6df6a1291e50c04ab[flogtanh_SEL-1:0]),
.flogtanh( I2ad2ede07f1ffac643211e88bf8ddbd6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2493237a24acdcab8b5bda10e804a5cf = (Ib5d28d8f73d17ab6df6a1291e50c04ab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2ad2ede07f1ffac643211e88bf8ddbd6;


Ic3da32f100a43f826b89a492544e7812 I6941e562ade82b683e5f3b8ad17ccbc7 (
.flogtanh_sel( I81259f391db792339824ad5dd1a0057b[flogtanh_SEL-1:0]),
.flogtanh( I5bc390dc300be5f8bc85f928cca1cd0b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I03829256e357ac17c7ca7cae2f980f41 = (I81259f391db792339824ad5dd1a0057b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5bc390dc300be5f8bc85f928cca1cd0b;


Ic3da32f100a43f826b89a492544e7812 I24b8ce3ca389446adc0feaa7fab6ca27 (
.flogtanh_sel( I6f09ac63effe67a86798b9b4e1690664[flogtanh_SEL-1:0]),
.flogtanh( I3e7efaed64fd3c276e882ab38109d538),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iae32c44b88fe7ddb5d4f19cf8fff3ba6 = (I6f09ac63effe67a86798b9b4e1690664[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3e7efaed64fd3c276e882ab38109d538;


Ic3da32f100a43f826b89a492544e7812 I0af6c221991a0c2c636862815770c96c (
.flogtanh_sel( I370b4b3a0048a93ba374a40e170c75a3[flogtanh_SEL-1:0]),
.flogtanh( Ib4738fe629dbe40eefed821b40ab93c8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3bdc5ba374f85dc61346e4868c41a6bf = (I370b4b3a0048a93ba374a40e170c75a3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib4738fe629dbe40eefed821b40ab93c8;


Ic3da32f100a43f826b89a492544e7812 I522e6f7238a032757ea7b0831259150d (
.flogtanh_sel( I3f8476d0aa0ea2439b67ea1a4adf36c5[flogtanh_SEL-1:0]),
.flogtanh( I30268ed341753c3ab53b65ad43e94923),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I557ef77ce931535467a07a8d70145f55 = (I3f8476d0aa0ea2439b67ea1a4adf36c5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I30268ed341753c3ab53b65ad43e94923;


Ic3da32f100a43f826b89a492544e7812 I3c1298b29a025ebefa8231ab0a5f272e (
.flogtanh_sel( I35b52dba10a8a5b22b518388fecac82d[flogtanh_SEL-1:0]),
.flogtanh( I2f10be9cbe2a935475077c0218031a5a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib4695d4389db72c5ac7e31809072c290 = (I35b52dba10a8a5b22b518388fecac82d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2f10be9cbe2a935475077c0218031a5a;


Ic3da32f100a43f826b89a492544e7812 I7eb710a694aae2d7a7ef26692d166951 (
.flogtanh_sel( Ic7db274ed18e6fdecf30381a31238777[flogtanh_SEL-1:0]),
.flogtanh( I41d598b80334ab12e5f53b2a6c721517),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie81315a3a14a5ef879d8e3f405936365 = (Ic7db274ed18e6fdecf30381a31238777[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41d598b80334ab12e5f53b2a6c721517;


Ic3da32f100a43f826b89a492544e7812 I6a412c77417f42ee1aa6d365136b63f5 (
.flogtanh_sel( I2c4e538a8db759e9799541d9178ec61e[flogtanh_SEL-1:0]),
.flogtanh( I94b3d895ee69e3ab482ff1aa0798c92a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia7520053a7c4a94437c6a780b03a28a5 = (I2c4e538a8db759e9799541d9178ec61e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I94b3d895ee69e3ab482ff1aa0798c92a;


Ic3da32f100a43f826b89a492544e7812 Icb9398effd2fabf7710469815644f351 (
.flogtanh_sel( Ief6d4c3f5ef8663e111ef99347b023f5[flogtanh_SEL-1:0]),
.flogtanh( I24a25d4725db6bcb4732fa21bc861736),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic308a5413f38b96d244cac3b0bc9462c = (Ief6d4c3f5ef8663e111ef99347b023f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I24a25d4725db6bcb4732fa21bc861736;


Ic3da32f100a43f826b89a492544e7812 I27d97e206c939b80017dc8b1fd982b55 (
.flogtanh_sel( Id95e964e5faecb52c72669b0d28a4bf5[flogtanh_SEL-1:0]),
.flogtanh( I1877b73e028c908de9dc734b93cbf8bb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I034fb3850485fae2d1358041a1c41888 = (Id95e964e5faecb52c72669b0d28a4bf5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1877b73e028c908de9dc734b93cbf8bb;


Ic3da32f100a43f826b89a492544e7812 I13829e46ba8fc5b6bbce459cbff9ab9b (
.flogtanh_sel( I0fcef4538102ac6d24aa7090d5405afa[flogtanh_SEL-1:0]),
.flogtanh( Ic99b64430e5dfdabe3634fbddeb41b3c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0e7079db66c15210046b997f319ece89 = (I0fcef4538102ac6d24aa7090d5405afa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic99b64430e5dfdabe3634fbddeb41b3c;


Ic3da32f100a43f826b89a492544e7812 Id99936a0ccafb9ea53b4e461beea6e1d (
.flogtanh_sel( I055019e38eec6badd1739033d43d7d97[flogtanh_SEL-1:0]),
.flogtanh( I3c0ddec6d702a344930fd04f923bb2f1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9a5388f8aa6e9924a309aa8db4c1983b = (I055019e38eec6badd1739033d43d7d97[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3c0ddec6d702a344930fd04f923bb2f1;


Ic3da32f100a43f826b89a492544e7812 I3ebda9889e06310deb71057e4d9da07c (
.flogtanh_sel( I35c20a6e823da77a870b421eef2e0a95[flogtanh_SEL-1:0]),
.flogtanh( I41829e511abe1ddf9b67f899143db19a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ief76663994991118b1899ea4ddf4527d = (I35c20a6e823da77a870b421eef2e0a95[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41829e511abe1ddf9b67f899143db19a;


Ic3da32f100a43f826b89a492544e7812 I8b185066080134fe483f4b004decda7f (
.flogtanh_sel( I32cc12cdacef1a4ef64577e0fa977f46[flogtanh_SEL-1:0]),
.flogtanh( I41961139f5b650e4f4ba5c2eadda6702),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6fb63ea54e492bdbc6d1145affc683e9 = (I32cc12cdacef1a4ef64577e0fa977f46[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41961139f5b650e4f4ba5c2eadda6702;


Ic3da32f100a43f826b89a492544e7812 I4642cdcc784f7b1f6cfdb6a1147e4113 (
.flogtanh_sel( I26b3f2360ca4a8caee61b2f3a3a08267[flogtanh_SEL-1:0]),
.flogtanh( I8ef0ac3bf43f16d2edf5a5045b0eb498),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If83ce1cbe3a73472419520c225b288a6 = (I26b3f2360ca4a8caee61b2f3a3a08267[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8ef0ac3bf43f16d2edf5a5045b0eb498;


Ic3da32f100a43f826b89a492544e7812 Iafcc6c2f2e91f48fe8ec3c769902d9b6 (
.flogtanh_sel( I5ef9b7dc0c63e9ca6a5fb5f7ffa06041[flogtanh_SEL-1:0]),
.flogtanh( I4084e3c9ba635fc4a8d281015bdeb33a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id1df78ab32daf524b77c0431c782f2bf = (I5ef9b7dc0c63e9ca6a5fb5f7ffa06041[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4084e3c9ba635fc4a8d281015bdeb33a;


Ic3da32f100a43f826b89a492544e7812 Ib6f233f249dc9c2e56b42e93e6c3e762 (
.flogtanh_sel( If881473b05090f40a027d7eeee7f7ed9[flogtanh_SEL-1:0]),
.flogtanh( I199a14038a0ff6ac25dab60162f8c6c9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iff142b88493149045fc0de355b767c16 = (If881473b05090f40a027d7eeee7f7ed9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I199a14038a0ff6ac25dab60162f8c6c9;


Ic3da32f100a43f826b89a492544e7812 I121f3fcc436b61efeb0723173ea0ae2c (
.flogtanh_sel( I23bd59ab5b038935301396aaf2acefc1[flogtanh_SEL-1:0]),
.flogtanh( Ic6859263f79d29d5f4896d85367be2bf),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I28c3818247c7c6de11790f6692882b5a = (I23bd59ab5b038935301396aaf2acefc1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic6859263f79d29d5f4896d85367be2bf;


Ic3da32f100a43f826b89a492544e7812 I5a9a39b65842a94cca38b59ae4c4e851 (
.flogtanh_sel( I874386d94dacf84e699d159af1a49836[flogtanh_SEL-1:0]),
.flogtanh( If0af3259e321390fffe518318f0f2545),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib451127b69a0a800332a712af77c6d29 = (I874386d94dacf84e699d159af1a49836[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If0af3259e321390fffe518318f0f2545;


Ic3da32f100a43f826b89a492544e7812 I26f612f5fe48f0048cb12e6ca101489c (
.flogtanh_sel( I95bfe51a759bf4165168e5e3b99d6b34[flogtanh_SEL-1:0]),
.flogtanh( Icafbf36da24f4db99e0ce4eeca6ca338),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3d601db540da359ae4d22f960d3d5af8 = (I95bfe51a759bf4165168e5e3b99d6b34[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icafbf36da24f4db99e0ce4eeca6ca338;


Ic3da32f100a43f826b89a492544e7812 I51f325914c5d23cde8d920113455f649 (
.flogtanh_sel( I4ba5b2f9b7ec0937ecd2c9945cf6de87[flogtanh_SEL-1:0]),
.flogtanh( Ia614303d31afc0ef4f15ec5b43231cd8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2c1f2476efe593829ade470fe8ec2526 = (I4ba5b2f9b7ec0937ecd2c9945cf6de87[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia614303d31afc0ef4f15ec5b43231cd8;


Ic3da32f100a43f826b89a492544e7812 Ic0482656a2c4a41df942eb453675f690 (
.flogtanh_sel( I0b08fb8db0e8a1de3d416907c87fe700[flogtanh_SEL-1:0]),
.flogtanh( I28ff2f86da2016b00bd0c21cbd1b4530),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7e685b06df8a8c2ac351fa9f9b76a81d = (I0b08fb8db0e8a1de3d416907c87fe700[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I28ff2f86da2016b00bd0c21cbd1b4530;


Ic3da32f100a43f826b89a492544e7812 Id7783cf1ec7c6601d6f0e300492d028f (
.flogtanh_sel( Ie030d12e5acf9ef4975a17c83b2481c1[flogtanh_SEL-1:0]),
.flogtanh( I2b8c969c11b4117c96470f4f6ed6963a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1338d211b5d2d409bfe0df76d2ca2701 = (Ie030d12e5acf9ef4975a17c83b2481c1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2b8c969c11b4117c96470f4f6ed6963a;


Ic3da32f100a43f826b89a492544e7812 Idb18f5c32cf359a0203c379c478f8aee (
.flogtanh_sel( Ia7a0e852d3dfcef950804ea0ebb0c80a[flogtanh_SEL-1:0]),
.flogtanh( Iea563639beb7fcb0291b5dc1410951d1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia40dad546d9c852e2fa8942c62a1c1f8 = (Ia7a0e852d3dfcef950804ea0ebb0c80a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iea563639beb7fcb0291b5dc1410951d1;


Ic3da32f100a43f826b89a492544e7812 I65da849c49d4f57f51632d8d12b93a0a (
.flogtanh_sel( Iaa4c38d030eab2b7899399aa0d7886d9[flogtanh_SEL-1:0]),
.flogtanh( Ic1b35046657e23f42199e39343a652a8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0b0dd019d8bd24684403a29aed668b6d = (Iaa4c38d030eab2b7899399aa0d7886d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic1b35046657e23f42199e39343a652a8;


Ic3da32f100a43f826b89a492544e7812 I81e515bf9212a3187e79f2f6cd90f773 (
.flogtanh_sel( Icce7ff1d652d4d9c2be5ecf679059bbe[flogtanh_SEL-1:0]),
.flogtanh( Ie7b26120ee77b43574c1ca171d7ec15f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I66a304016a9adfd85a2abb6f8fd39afc = (Icce7ff1d652d4d9c2be5ecf679059bbe[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie7b26120ee77b43574c1ca171d7ec15f;


Ic3da32f100a43f826b89a492544e7812 Iec265fe8ef7994a35765a896718571ea (
.flogtanh_sel( If816bc5eacaea23443602e575ddf60b8[flogtanh_SEL-1:0]),
.flogtanh( I2ed61ced1577d905da91d97592006ed5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I177be24718c59688752097fe2a4085c4 = (If816bc5eacaea23443602e575ddf60b8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2ed61ced1577d905da91d97592006ed5;


Ic3da32f100a43f826b89a492544e7812 I8566d28aa1617f0caa389da0d165a4b0 (
.flogtanh_sel( I3b224a4ded05446cc5300d430bdd1947[flogtanh_SEL-1:0]),
.flogtanh( I332dc26a52194745d19c4d8468e42864),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7e66a42eb7cdb820cd1297c39f0625e8 = (I3b224a4ded05446cc5300d430bdd1947[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I332dc26a52194745d19c4d8468e42864;


Ic3da32f100a43f826b89a492544e7812 I6bb1c4da921bdcfbf76302d05095a181 (
.flogtanh_sel( Ia5fc5cfb0e52237b407b37a3858fccb5[flogtanh_SEL-1:0]),
.flogtanh( Ibb4fefe05e94e055e86a743c40fb1c5e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If2021f0735c6c5649ebac0d230fda87c = (Ia5fc5cfb0e52237b407b37a3858fccb5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibb4fefe05e94e055e86a743c40fb1c5e;


Ic3da32f100a43f826b89a492544e7812 I262b2147b6af9de68adc9647d8557ed9 (
.flogtanh_sel( I92f8ba6e7f8e9b30fb5b6973eb8fd03e[flogtanh_SEL-1:0]),
.flogtanh( Ia56a76a20d4f11b0e80cbe31820a6977),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie1bf5d97b8f679095d2442bbf9f95608 = (I92f8ba6e7f8e9b30fb5b6973eb8fd03e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia56a76a20d4f11b0e80cbe31820a6977;


Ic3da32f100a43f826b89a492544e7812 I51b828072aab378fe0004e98f00c2428 (
.flogtanh_sel( Icdfa60d2a024dd934f7e6639c6cb2c28[flogtanh_SEL-1:0]),
.flogtanh( I054ebc7f9e3da325ba0c6e329f2ee770),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I632469889d6bb1c268b45fb805467ebd = (Icdfa60d2a024dd934f7e6639c6cb2c28[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I054ebc7f9e3da325ba0c6e329f2ee770;


Ic3da32f100a43f826b89a492544e7812 Id516db9d9b9cdf399c3f4676c3eb2892 (
.flogtanh_sel( Ifff70b976513eaa42b6bd4b80c98611e[flogtanh_SEL-1:0]),
.flogtanh( I3361df26cc86ca8be1653d9376d0c8e0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie230ba3c73808e102eee9e5868595e7c = (Ifff70b976513eaa42b6bd4b80c98611e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3361df26cc86ca8be1653d9376d0c8e0;


Ic3da32f100a43f826b89a492544e7812 Ie2568aa361a3cf5a8fc9a1f5026c4778 (
.flogtanh_sel( Ica12fa8b631b70a6bbe9f6e92bf73ea0[flogtanh_SEL-1:0]),
.flogtanh( I586fbde80f0130c4a6ead49de11efdd9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie1e9326e4eee006ec07abb6bb7d269a5 = (Ica12fa8b631b70a6bbe9f6e92bf73ea0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I586fbde80f0130c4a6ead49de11efdd9;


Ic3da32f100a43f826b89a492544e7812 Id116c201b0363bd0be5816b4f5e83d41 (
.flogtanh_sel( Ie69c255335760f706c644b115887269b[flogtanh_SEL-1:0]),
.flogtanh( Ifa087137c8a6028b13bfa95aba19fc34),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ica4ec1647bdb5a3aad6db6b447bd7995 = (Ie69c255335760f706c644b115887269b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifa087137c8a6028b13bfa95aba19fc34;


Ic3da32f100a43f826b89a492544e7812 Ieac043faee94714c30338260c72e2917 (
.flogtanh_sel( Idb06676b41de19bc86eae34c292183d9[flogtanh_SEL-1:0]),
.flogtanh( I51a3a6c79c488c092394375891775be3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia17295aec0a40c2b46a595dacfede2d5 = (Idb06676b41de19bc86eae34c292183d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I51a3a6c79c488c092394375891775be3;


Ic3da32f100a43f826b89a492544e7812 I4c1b9599327d309a36cdaa2cd380701b (
.flogtanh_sel( Ib21d2306d5ded3406fac754e69a10d20[flogtanh_SEL-1:0]),
.flogtanh( I01a7ebdc760227ee40b85828e28238a9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4c6d3d6fc2d10066a744fdd9405a7902 = (Ib21d2306d5ded3406fac754e69a10d20[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I01a7ebdc760227ee40b85828e28238a9;


Ic3da32f100a43f826b89a492544e7812 If0a567f015e289af7d5a2d4549ea6dbd (
.flogtanh_sel( Ib41d1aa2dcf81879976fb8964cbf6f79[flogtanh_SEL-1:0]),
.flogtanh( Ib3f9e4c05e363069775e5de9d240b3dc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia9c043c5e8873fd13e39cf6bd8136c51 = (Ib41d1aa2dcf81879976fb8964cbf6f79[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib3f9e4c05e363069775e5de9d240b3dc;


Ic3da32f100a43f826b89a492544e7812 I327a176d4b4f634e6d8346b56f014f5a (
.flogtanh_sel( I5f8f5e246f008b8d8c75f72828337bab[flogtanh_SEL-1:0]),
.flogtanh( I18664482dcc1371fa4b915af96070539),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2e802c75c6ce34b05943b678ecbfacb1 = (I5f8f5e246f008b8d8c75f72828337bab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I18664482dcc1371fa4b915af96070539;


Ic3da32f100a43f826b89a492544e7812 I89ab48c6472fa84fd8577017fb6be26c (
.flogtanh_sel( Id6625e78da0e14d2eeb19cc8ac6520e0[flogtanh_SEL-1:0]),
.flogtanh( I6a41c6cf78cb25ad1c47550756449002),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieb3f28762410fb40a0c8a8556b4b3ca0 = (Id6625e78da0e14d2eeb19cc8ac6520e0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6a41c6cf78cb25ad1c47550756449002;


Ic3da32f100a43f826b89a492544e7812 Icd3bf02fa1fed76e992180c026ad3771 (
.flogtanh_sel( I6d9ddc6afa559ac35c042df1a9390ce9[flogtanh_SEL-1:0]),
.flogtanh( Iaf660a97d66e0d7f8e26f65229b7683f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie3e0c0e40c7a67ce7f957e74bd2a895d = (I6d9ddc6afa559ac35c042df1a9390ce9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaf660a97d66e0d7f8e26f65229b7683f;


Ic3da32f100a43f826b89a492544e7812 Iee3d2f745d4715e69e78e2705b1f1204 (
.flogtanh_sel( I9334055c7833676469670372d3c5cc31[flogtanh_SEL-1:0]),
.flogtanh( I7ded197ff64af1bce0e0d85705900a42),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I491f2373b2df19a4c22e1787ef034179 = (I9334055c7833676469670372d3c5cc31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7ded197ff64af1bce0e0d85705900a42;


Ic3da32f100a43f826b89a492544e7812 Ib8378fbe79e7712a8c7fc9f57bac9bac (
.flogtanh_sel( I0c97d772c737c6ff85b584bf69ccaf93[flogtanh_SEL-1:0]),
.flogtanh( I7c06179d5424165f8a805754834fd98c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ief96603d41b4f670d2bbfa3d3875c903 = (I0c97d772c737c6ff85b584bf69ccaf93[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7c06179d5424165f8a805754834fd98c;


Ic3da32f100a43f826b89a492544e7812 Ia85a41c28b364302b42310dc783dafdc (
.flogtanh_sel( Ic6ce97ae85d91dd8a79f3f9d0da375a2[flogtanh_SEL-1:0]),
.flogtanh( Id364f2a517a0f3109564a025ffd8eec3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7a029c27d92754041eb6d605837238dd = (Ic6ce97ae85d91dd8a79f3f9d0da375a2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id364f2a517a0f3109564a025ffd8eec3;


Ic3da32f100a43f826b89a492544e7812 I9cd35c24488c360891a391071ac99236 (
.flogtanh_sel( I83ff9a2750b298b0f7c9b6ce13f574af[flogtanh_SEL-1:0]),
.flogtanh( Ie3ea12584ed3e255073776620d778f06),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I00dad36628d2fa923120fdaa79bf0045 = (I83ff9a2750b298b0f7c9b6ce13f574af[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie3ea12584ed3e255073776620d778f06;


Ic3da32f100a43f826b89a492544e7812 Ibabe30d8e65e61d7d26f161a8322af84 (
.flogtanh_sel( I85699a2a05c343a6a9e828af6d445e9e[flogtanh_SEL-1:0]),
.flogtanh( I38d885c58b4f7333c679b0b5783418df),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3707f68de059df0af5c652fc0478e543 = (I85699a2a05c343a6a9e828af6d445e9e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I38d885c58b4f7333c679b0b5783418df;


Ic3da32f100a43f826b89a492544e7812 Id7eeaf580c8bca664af9ec729ae6448b (
.flogtanh_sel( I51f6e39b24b2554884e381be79f47ff2[flogtanh_SEL-1:0]),
.flogtanh( I69251440f80eb2e177307aec4cb0111f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I94af4b6b9dc11935db54ba872889392d = (I51f6e39b24b2554884e381be79f47ff2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I69251440f80eb2e177307aec4cb0111f;


Ic3da32f100a43f826b89a492544e7812 Id66892f49e9605c15615668db8dac71e (
.flogtanh_sel( I9f65fd05c6929300860c8cbbde5607f2[flogtanh_SEL-1:0]),
.flogtanh( I0a9bcd4a3b79b003b5df8afa0d6b6782),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I38e2dbba093928b874d447362d89b291 = (I9f65fd05c6929300860c8cbbde5607f2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0a9bcd4a3b79b003b5df8afa0d6b6782;


Ic3da32f100a43f826b89a492544e7812 I2eaa9a85d8cd78b7310449d3c95bc0b6 (
.flogtanh_sel( If09761d8f06051d4287ee29ac9c9fa19[flogtanh_SEL-1:0]),
.flogtanh( I36569656996bf98bce33b2d7a4b79def),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia48f0029e9e76386f3dd70aacd9adbfa = (If09761d8f06051d4287ee29ac9c9fa19[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I36569656996bf98bce33b2d7a4b79def;


Ic3da32f100a43f826b89a492544e7812 I2e9b0778263e734d37c98896710cdeab (
.flogtanh_sel( I33bfbe0bcca6d32c86b9576577e3f265[flogtanh_SEL-1:0]),
.flogtanh( I7e408a50d0511909aeb57d5a00535e80),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic2b20168744fafbe15037ed7fa83da72 = (I33bfbe0bcca6d32c86b9576577e3f265[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7e408a50d0511909aeb57d5a00535e80;


Ic3da32f100a43f826b89a492544e7812 I072d1881db0aa7efe8ecc05bb51e8b49 (
.flogtanh_sel( If2921210b1c05ecbf00af3a2bcb96ef4[flogtanh_SEL-1:0]),
.flogtanh( Iacc6f48dd92dc515be06a681cc5b56e9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I62fdc8936121a2707d94cf3bd6e660ac = (If2921210b1c05ecbf00af3a2bcb96ef4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iacc6f48dd92dc515be06a681cc5b56e9;


Ic3da32f100a43f826b89a492544e7812 If2f079694ac286bbb54d894bfaebacd4 (
.flogtanh_sel( Ib074e38e280474a782da831a3e0028b4[flogtanh_SEL-1:0]),
.flogtanh( Icafa051878ad3421c31ed2550ea09945),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia0932b3fd6a5ae6da2bacd2b86ba3a43 = (Ib074e38e280474a782da831a3e0028b4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icafa051878ad3421c31ed2550ea09945;


Ic3da32f100a43f826b89a492544e7812 I22bbcccdd11972432c810c8de5e34cde (
.flogtanh_sel( I507449dde0bc0c8f53a10759436ec731[flogtanh_SEL-1:0]),
.flogtanh( If4e4f2776b1467e4f03bf15ff5f43c04),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9fce6091885f1bb97d29fb1f543b1a38 = (I507449dde0bc0c8f53a10759436ec731[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If4e4f2776b1467e4f03bf15ff5f43c04;


Ic3da32f100a43f826b89a492544e7812 Ibea18c7e11276eab9ad397ede48bfd68 (
.flogtanh_sel( Id55a3e3f2d75baeba71a345fad695c69[flogtanh_SEL-1:0]),
.flogtanh( I9387cd07e38260005bb3e41807d2d794),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib402cdbfaa9900820b85bd625415c547 = (Id55a3e3f2d75baeba71a345fad695c69[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9387cd07e38260005bb3e41807d2d794;


Ic3da32f100a43f826b89a492544e7812 I2d76dfc24db66cc0c6a14cf44327988e (
.flogtanh_sel( I20984f43d22671639a7a178ad15aec04[flogtanh_SEL-1:0]),
.flogtanh( I8bede290f421e6a05e49244f0d1d3d9b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I518a2736384c14c02f27bfa3d8ea7aff = (I20984f43d22671639a7a178ad15aec04[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8bede290f421e6a05e49244f0d1d3d9b;


Ic3da32f100a43f826b89a492544e7812 Ia25af39efe557c4035dc5288c9c70950 (
.flogtanh_sel( I59f88336d6bdd50ded87d353fb5ce3e9[flogtanh_SEL-1:0]),
.flogtanh( I6d8c2489fdeb42411f2e12bfa30752d2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I847cf7ff866f8a666872c12d6b67b1b1 = (I59f88336d6bdd50ded87d353fb5ce3e9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6d8c2489fdeb42411f2e12bfa30752d2;


Ic3da32f100a43f826b89a492544e7812 I4a1cec3f6223dd21367c98754a421dad (
.flogtanh_sel( I488635e3f7ed77ea88199f5bffd4b1d6[flogtanh_SEL-1:0]),
.flogtanh( I082715d1b8943faf11d464087542a83e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9e45e3d7117ce48cdbfc5db8c0ccfcf4 = (I488635e3f7ed77ea88199f5bffd4b1d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I082715d1b8943faf11d464087542a83e;


Ic3da32f100a43f826b89a492544e7812 I319bf3ed0bb8bb73bceb61e61c006e79 (
.flogtanh_sel( Ie6893017d21c050ba10d206854f4a9f4[flogtanh_SEL-1:0]),
.flogtanh( I4de91d9613edc5c4d096b717d9df5de4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I380ff8528cdba4026fac3c4eda8b2c52 = (Ie6893017d21c050ba10d206854f4a9f4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4de91d9613edc5c4d096b717d9df5de4;


Ic3da32f100a43f826b89a492544e7812 I6f4b9e87f3f0c32aa7ec7cb65a324661 (
.flogtanh_sel( Id3f68b4dc0ab60673208b7d2081f3533[flogtanh_SEL-1:0]),
.flogtanh( Ifb2a91a74b87c75592cb046b9bfd9c8b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iee8f9b0654f6f6797f11cae0947e454e = (Id3f68b4dc0ab60673208b7d2081f3533[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifb2a91a74b87c75592cb046b9bfd9c8b;


Ic3da32f100a43f826b89a492544e7812 I6ff351439834adce959f6c0390a19d5c (
.flogtanh_sel( I433756b944e061a824a89bda241e879f[flogtanh_SEL-1:0]),
.flogtanh( Ie21cffaecd7fe37601dcaef49a0d6cc3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie3e54a4700d8d0f6478187e06cb6f85d = (I433756b944e061a824a89bda241e879f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie21cffaecd7fe37601dcaef49a0d6cc3;


Ic3da32f100a43f826b89a492544e7812 I830435fb2e45dcef0eda0dd90c348029 (
.flogtanh_sel( I2eb60a922aa4f7482dd92b9351d53a2d[flogtanh_SEL-1:0]),
.flogtanh( Ia648c9d395ad2727209229807b4224fb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8c0069e8756bcff203ce21ae3170aa42 = (I2eb60a922aa4f7482dd92b9351d53a2d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia648c9d395ad2727209229807b4224fb;


Ic3da32f100a43f826b89a492544e7812 Ide03d1a2b9d28adc0e2cb1c9c838eb32 (
.flogtanh_sel( I0867979e1b159c8ceae548930376f482[flogtanh_SEL-1:0]),
.flogtanh( Ib415da845b88e5a8261beaf88b7ec804),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I856eada207c5006beb8f83f01d5d74c9 = (I0867979e1b159c8ceae548930376f482[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib415da845b88e5a8261beaf88b7ec804;


Ic3da32f100a43f826b89a492544e7812 I234ce778264c8b20f4b608ea9ff0a601 (
.flogtanh_sel( I4accfbeae8a5ee0dbeab23ef3a116145[flogtanh_SEL-1:0]),
.flogtanh( I6dffcf934a74385aa716db9d7fa29ed1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I79a46279070c53678a5af54f661c5821 = (I4accfbeae8a5ee0dbeab23ef3a116145[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6dffcf934a74385aa716db9d7fa29ed1;


Ic3da32f100a43f826b89a492544e7812 Ifb32dc14449c33aacd9e7d2fa3c0e374 (
.flogtanh_sel( Ic7570b0b7c5bef5758f68562ae4c90f6[flogtanh_SEL-1:0]),
.flogtanh( I13383df545ed8620a17a4fc2493cd770),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ica807adc510a2e32580ca77c18ea0b45 = (Ic7570b0b7c5bef5758f68562ae4c90f6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I13383df545ed8620a17a4fc2493cd770;


Ic3da32f100a43f826b89a492544e7812 I862601ed2d128662f621988b2cc7883d (
.flogtanh_sel( Iceadadc4456881fdeea85934a9bf4d6c[flogtanh_SEL-1:0]),
.flogtanh( I87ea43bfae8fad4e4c26741fd2de5b41),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia8094903aed8dd0ce8e9ff459a5287b0 = (Iceadadc4456881fdeea85934a9bf4d6c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I87ea43bfae8fad4e4c26741fd2de5b41;


Ic3da32f100a43f826b89a492544e7812 I57e79f137181e794b470f68ed52d559e (
.flogtanh_sel( I7b2b617ae67424f54961eebce42de77e[flogtanh_SEL-1:0]),
.flogtanh( I6d2022ba184980b8e5bc5edb4f4b0ff3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie018f3003c5f124bddd13c359257bf35 = (I7b2b617ae67424f54961eebce42de77e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6d2022ba184980b8e5bc5edb4f4b0ff3;


Ic3da32f100a43f826b89a492544e7812 Ic2f5c45a433c880b4c64b3f9b8002843 (
.flogtanh_sel( I953f0f8af76f89b2d9ab4abf19fb411d[flogtanh_SEL-1:0]),
.flogtanh( I68f98b68c9a3836d0c7dc152a2d441da),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice18bceb10fec484ffc96155e14c4974 = (I953f0f8af76f89b2d9ab4abf19fb411d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I68f98b68c9a3836d0c7dc152a2d441da;


Ic3da32f100a43f826b89a492544e7812 Id9c0665ceb8e62c7e6f017cb57c8f9d5 (
.flogtanh_sel( I915b4736dcb20f831d02e48f4e79f008[flogtanh_SEL-1:0]),
.flogtanh( I2dc3cec85c37aa943f01df545f952e05),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib484aa64b795f7e36198b800f302164f = (I915b4736dcb20f831d02e48f4e79f008[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2dc3cec85c37aa943f01df545f952e05;


Ic3da32f100a43f826b89a492544e7812 I0383416cc22272ced165deb846f3d355 (
.flogtanh_sel( Ib7eec587348ae1ca1f00c0a3ad10ad27[flogtanh_SEL-1:0]),
.flogtanh( Ieed49c262f87c86b30d94e9842525ab0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icdb143a4ce96029c2441758bf2edd7b0 = (Ib7eec587348ae1ca1f00c0a3ad10ad27[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieed49c262f87c86b30d94e9842525ab0;


Ic3da32f100a43f826b89a492544e7812 I2eb4ba9ff4cfb78040c5aa6eeb7343c9 (
.flogtanh_sel( I001a212686304248c8359e5fc01227c0[flogtanh_SEL-1:0]),
.flogtanh( Ib9ab475010c98fc4e06df5c98944387a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3a76f70ca3bfbcacc6f3342aa71f1912 = (I001a212686304248c8359e5fc01227c0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib9ab475010c98fc4e06df5c98944387a;


Ic3da32f100a43f826b89a492544e7812 I5874aee015469d98ed78c6c67b4eb404 (
.flogtanh_sel( Ibb7554e012c0fc1223c29b759c900666[flogtanh_SEL-1:0]),
.flogtanh( If7c8bdd5bae4a1bffd4bd2c8015bb738),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9470c7ab9634c01bb832c9e4ff5496bf = (Ibb7554e012c0fc1223c29b759c900666[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If7c8bdd5bae4a1bffd4bd2c8015bb738;


Ic3da32f100a43f826b89a492544e7812 I2af67887325023976a5c57088ba3095c (
.flogtanh_sel( I9aeb9c42b54a05be6bf9b7b88b6860ba[flogtanh_SEL-1:0]),
.flogtanh( I6463249144cd032e1c5af9e2987254b3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I218ee96418a4f5d734d3d71685bc09c7 = (I9aeb9c42b54a05be6bf9b7b88b6860ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6463249144cd032e1c5af9e2987254b3;


Ic3da32f100a43f826b89a492544e7812 I26de7d69716f4a0cf26ec60db35b37d8 (
.flogtanh_sel( I6a5a5966965b0790b906c6fda71aef80[flogtanh_SEL-1:0]),
.flogtanh( I5f9e468fc1bc199574d719d866d52dfc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I924514226fdb5bac110a2650bcb2e85f = (I6a5a5966965b0790b906c6fda71aef80[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5f9e468fc1bc199574d719d866d52dfc;


Ic3da32f100a43f826b89a492544e7812 I3e741d7243a368670dd3a241a7a83c71 (
.flogtanh_sel( Ic943083ca65ace6c42d73f4234739a06[flogtanh_SEL-1:0]),
.flogtanh( Ie69f792c606c3162052840dec732ef99),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idc57f37015a48393608e2b026bc7065c = (Ic943083ca65ace6c42d73f4234739a06[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie69f792c606c3162052840dec732ef99;


Ic3da32f100a43f826b89a492544e7812 Id57bee50431a45fb525cfe2a9589af9c (
.flogtanh_sel( Id0b321686d4c39621024cf0dd99822dc[flogtanh_SEL-1:0]),
.flogtanh( If874254c3c6813ff0d5184b574cb613d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I41af7e4c97fc04154fe6de66b82499f5 = (Id0b321686d4c39621024cf0dd99822dc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If874254c3c6813ff0d5184b574cb613d;


Ic3da32f100a43f826b89a492544e7812 I38930a94c726f0e24181ecb0f18c5939 (
.flogtanh_sel( I0839dd3787442f1b79b87e02436bfdce[flogtanh_SEL-1:0]),
.flogtanh( I90969c917df8480d379afef834c1a253),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I972bee4216f8e532e8fa4bd25fbb9c57 = (I0839dd3787442f1b79b87e02436bfdce[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I90969c917df8480d379afef834c1a253;


Ic3da32f100a43f826b89a492544e7812 I820f0f282d105391060a29b9a09d6004 (
.flogtanh_sel( I89e6a9fd97d8aa4dd3b832c3be4697b2[flogtanh_SEL-1:0]),
.flogtanh( I07280ae3417855f994980fbb95696fc6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib303ea0240e7ab5f000dd10e975b2274 = (I89e6a9fd97d8aa4dd3b832c3be4697b2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I07280ae3417855f994980fbb95696fc6;


Ic3da32f100a43f826b89a492544e7812 I2e46fb44deeb7be89b7c248d229311b3 (
.flogtanh_sel( I93d4157f48b132642752220059861e98[flogtanh_SEL-1:0]),
.flogtanh( I852c62fffff0fd7bf06939d75fada3eb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5971253546899e9a82f387d5eabcc7b3 = (I93d4157f48b132642752220059861e98[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I852c62fffff0fd7bf06939d75fada3eb;


Ic3da32f100a43f826b89a492544e7812 I935e5947e5cfaf00fe77699c0f264fdf (
.flogtanh_sel( I8fc4faa2891d7fd3479ac1f788f481dc[flogtanh_SEL-1:0]),
.flogtanh( I9e0a2da5a82f1b509bd502554f4760aa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1fc36e6f738fab96df356979e1e3a612 = (I8fc4faa2891d7fd3479ac1f788f481dc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9e0a2da5a82f1b509bd502554f4760aa;


Ic3da32f100a43f826b89a492544e7812 I1405a927347431cd0456a03e4fdc7733 (
.flogtanh_sel( I440f30e9cb4bc89233b46ea00b4cbeb4[flogtanh_SEL-1:0]),
.flogtanh( I6293c2b405087f14b42b423336f6990c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie2d8c84d8c9a4c8f637068a2ae39fdde = (I440f30e9cb4bc89233b46ea00b4cbeb4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6293c2b405087f14b42b423336f6990c;


Ic3da32f100a43f826b89a492544e7812 Iff5e19522b593de1fc469a3b2d9e2045 (
.flogtanh_sel( I6568bfd8780c11e0b1b049a01f92abd8[flogtanh_SEL-1:0]),
.flogtanh( I70e8d96970e69bc828a6aea5ade3bdd1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I114c595caa67a3f777f087a634130a6d = (I6568bfd8780c11e0b1b049a01f92abd8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I70e8d96970e69bc828a6aea5ade3bdd1;


Ic3da32f100a43f826b89a492544e7812 I7f71fa758d8a6bccb8ee12b838e89e5e (
.flogtanh_sel( Ibf7dc4da07f9955d5d4c7e1f63f1ad68[flogtanh_SEL-1:0]),
.flogtanh( I0380003f741eedb994793c2cb7e6c5c3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idad14b6383b9af54eb35e72ff3d10035 = (Ibf7dc4da07f9955d5d4c7e1f63f1ad68[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0380003f741eedb994793c2cb7e6c5c3;


Ic3da32f100a43f826b89a492544e7812 I4bd026fcce91129b4492e4dac0c9f2d0 (
.flogtanh_sel( I7ec1a328587b72a39c462083efea0ee0[flogtanh_SEL-1:0]),
.flogtanh( Ia884fcfa49cfe0b404bf49b99d7381aa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I46e9c76b19ed1ff21f102efe6ee5c732 = (I7ec1a328587b72a39c462083efea0ee0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia884fcfa49cfe0b404bf49b99d7381aa;


Ic3da32f100a43f826b89a492544e7812 I5f3fc4f2a681697a319cd30c57a8e154 (
.flogtanh_sel( Iaf028e7ab4dc77a7649f15d603834b5f[flogtanh_SEL-1:0]),
.flogtanh( Ie4ecd4c122ea5b478f3d7d2d632b8bf4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic75b8bbb1b80001ec188a0cd25623420 = (Iaf028e7ab4dc77a7649f15d603834b5f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie4ecd4c122ea5b478f3d7d2d632b8bf4;


Ic3da32f100a43f826b89a492544e7812 I7fbb9ac306c75381eb0cdc9c0ba91645 (
.flogtanh_sel( I58db79a8e9f0cd1ded379897ba2f27ae[flogtanh_SEL-1:0]),
.flogtanh( I82e534ecaabf5af6a9b6a567b862800a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idc7df6877bdb7e7d392307d78183d31c = (I58db79a8e9f0cd1ded379897ba2f27ae[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I82e534ecaabf5af6a9b6a567b862800a;


Ic3da32f100a43f826b89a492544e7812 I314e342874790132007847ff962fb257 (
.flogtanh_sel( I6d3cb4ccb4e51c7e6603d0abd1a082c4[flogtanh_SEL-1:0]),
.flogtanh( I1c9684b45467216a18a3a0d93b555b60),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib8b95ece5da3877b261a06e6d0571921 = (I6d3cb4ccb4e51c7e6603d0abd1a082c4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1c9684b45467216a18a3a0d93b555b60;


Ic3da32f100a43f826b89a492544e7812 I91e1da6d6dd70d4e7c23e3ddaa316ac3 (
.flogtanh_sel( I79f75f49ea8a29d684af396014b2f3ab[flogtanh_SEL-1:0]),
.flogtanh( Ice212c509101d6d41b52ea0cb85dacc0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic99654bf4833c9132912eeb4c0dc92fa = (I79f75f49ea8a29d684af396014b2f3ab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ice212c509101d6d41b52ea0cb85dacc0;


Ic3da32f100a43f826b89a492544e7812 I841b063bbd36b902525008afbdc7a566 (
.flogtanh_sel( I9c5ecd86bedb189fada40fae9d751a68[flogtanh_SEL-1:0]),
.flogtanh( I37ee7a2fab22cf8e6452fb408b849595),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2461055ef9b1aa2ffca0f5cac3300e71 = (I9c5ecd86bedb189fada40fae9d751a68[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I37ee7a2fab22cf8e6452fb408b849595;


Ic3da32f100a43f826b89a492544e7812 I9874b247fb1d910d5192723a4a190a10 (
.flogtanh_sel( Iad5f06e1989ead7d306c70a3b02cb8f4[flogtanh_SEL-1:0]),
.flogtanh( I0ec18ade132eede6849e0607af608726),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2bc3ffbe5b42b0833206437d3863278e = (Iad5f06e1989ead7d306c70a3b02cb8f4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0ec18ade132eede6849e0607af608726;


Ic3da32f100a43f826b89a492544e7812 I013eb27b843435071f412ec694d6f71a (
.flogtanh_sel( If6d1a410df5a4aea6a01337a6074fbd9[flogtanh_SEL-1:0]),
.flogtanh( I4651eab27cb766a1792f9564bcb2764a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id5e02d4c48fa6c3b0d45a9e66f09448f = (If6d1a410df5a4aea6a01337a6074fbd9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4651eab27cb766a1792f9564bcb2764a;


Ic3da32f100a43f826b89a492544e7812 Ia3f03ecfe9f03d4dd5b6ffbdec97758f (
.flogtanh_sel( I3bc40a4db14566b5099b14cee5f61135[flogtanh_SEL-1:0]),
.flogtanh( Ibbdbc4e4fc2ee018a0e7a4da29e85b56),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I40e99289d5762e77a3766eb8251eef00 = (I3bc40a4db14566b5099b14cee5f61135[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibbdbc4e4fc2ee018a0e7a4da29e85b56;


Ic3da32f100a43f826b89a492544e7812 I6cfbee6ca5c87cab6ceb26f12b4fae8f (
.flogtanh_sel( I7e683fd8235d7cfbf4ff407a286f07de[flogtanh_SEL-1:0]),
.flogtanh( Ic67b9e090d6815b2a745bdc4983f9c69),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I20beb3fdbe91936f74a200cd8ec9817b = (I7e683fd8235d7cfbf4ff407a286f07de[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic67b9e090d6815b2a745bdc4983f9c69;


Ic3da32f100a43f826b89a492544e7812 I53c7313ce802bcbc3bfa4e79d8bd4bd7 (
.flogtanh_sel( I97afcedf05e588b7976d6005191dc916[flogtanh_SEL-1:0]),
.flogtanh( I8327267045af5da02c066a5eab25f13a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id435b68afb53bef4afc7b70a9512e955 = (I97afcedf05e588b7976d6005191dc916[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8327267045af5da02c066a5eab25f13a;


Ic3da32f100a43f826b89a492544e7812 I2db62d36b303fde7bebba334792a3abb (
.flogtanh_sel( Ib8d8eec0aaa662adf2837c9b705fce7e[flogtanh_SEL-1:0]),
.flogtanh( Id91ef7e27c689cdf5ce50d705017e40e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0cf5cb4cd472502b84dbf6fe1af0be78 = (Ib8d8eec0aaa662adf2837c9b705fce7e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id91ef7e27c689cdf5ce50d705017e40e;


Ic3da32f100a43f826b89a492544e7812 I14c72fec82d0b879797d0784f2ad1d39 (
.flogtanh_sel( Icbd765be950123705955e2c5d7ace84b[flogtanh_SEL-1:0]),
.flogtanh( I60498760f3c03cf92ceeb99c5096fe54),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iacf6340a29a5592b61ea875304a2de48 = (Icbd765be950123705955e2c5d7ace84b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I60498760f3c03cf92ceeb99c5096fe54;


Ic3da32f100a43f826b89a492544e7812 I0b31fd06b941d51f51d979646cf3a922 (
.flogtanh_sel( I706e8f5617cfae1e6fc83db18c8b5fe3[flogtanh_SEL-1:0]),
.flogtanh( I63169dbc533400e0db5e37a8ebeca1aa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5dfc71255cba279420b7545df4d35c40 = (I706e8f5617cfae1e6fc83db18c8b5fe3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I63169dbc533400e0db5e37a8ebeca1aa;


Ic3da32f100a43f826b89a492544e7812 If49963db7c7b6760b0885240683dc3f6 (
.flogtanh_sel( I1dd8f8c7f1b673898096b1f3ae383197[flogtanh_SEL-1:0]),
.flogtanh( I150f11a565ad39c59d8f9e4c94d397e2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibadcb205c7e9a0f3345cac7eb41b5985 = (I1dd8f8c7f1b673898096b1f3ae383197[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I150f11a565ad39c59d8f9e4c94d397e2;


Ic3da32f100a43f826b89a492544e7812 Id68006b668cee94fab9322a825640bb1 (
.flogtanh_sel( I10ca8978cf4659265ed25a27d09acc1c[flogtanh_SEL-1:0]),
.flogtanh( Icadb816a238ba165425e5a30bd0bb8e6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I762b2abb876381eff6de97cef0798405 = (I10ca8978cf4659265ed25a27d09acc1c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icadb816a238ba165425e5a30bd0bb8e6;


Ic3da32f100a43f826b89a492544e7812 I7720484859df47c067b4e0b7b90ff9fd (
.flogtanh_sel( Iec4656b32460def4a608b6b0f6486af9[flogtanh_SEL-1:0]),
.flogtanh( I3b55785b9625ac53f6c00ba5a10a481b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib3e7633767b6e09e4ee54f6feaddd31e = (Iec4656b32460def4a608b6b0f6486af9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3b55785b9625ac53f6c00ba5a10a481b;


Ic3da32f100a43f826b89a492544e7812 I9efa5ea2a3e65d52878299cbae06c711 (
.flogtanh_sel( I5f4475897d1d58965da1b35fe0ef8c01[flogtanh_SEL-1:0]),
.flogtanh( If7317c81c9b6503386cab33fa812e80e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3f193e9c265c1dfaeada63d59db5b79f = (I5f4475897d1d58965da1b35fe0ef8c01[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If7317c81c9b6503386cab33fa812e80e;


Ic3da32f100a43f826b89a492544e7812 Ic878f2a16139e52738789e775aab03d7 (
.flogtanh_sel( Ife61469306df3cf220666b187f1496a9[flogtanh_SEL-1:0]),
.flogtanh( I095672e79ca3a6dd8589b7821f06cdb9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie72268e979cf069b88f6eadde789e5ab = (Ife61469306df3cf220666b187f1496a9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I095672e79ca3a6dd8589b7821f06cdb9;


Ic3da32f100a43f826b89a492544e7812 I5cfcd8767987de774d2e2e4fdf338a86 (
.flogtanh_sel( Ib49319b9dfa4914f92f423ceaf840014[flogtanh_SEL-1:0]),
.flogtanh( Ibf2f43980e835dd7ae7535957e3ec131),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5732fdb805258fc13c8ba4aaf56574ca = (Ib49319b9dfa4914f92f423ceaf840014[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibf2f43980e835dd7ae7535957e3ec131;


Ic3da32f100a43f826b89a492544e7812 I80d830be15d6fa8044e96b2126c89f46 (
.flogtanh_sel( I93ff2f879233cac9b9f0dd2f4c082c09[flogtanh_SEL-1:0]),
.flogtanh( Iaa980a50205025e3e1b09c6ce8ee53dd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3afe987d8f2c93cc19534a3221d1939c = (I93ff2f879233cac9b9f0dd2f4c082c09[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaa980a50205025e3e1b09c6ce8ee53dd;


Ic3da32f100a43f826b89a492544e7812 I672efd0ba9cf19654adaaf2fba3b49c1 (
.flogtanh_sel( I44597d694e9c5d29280e503d72a27c8d[flogtanh_SEL-1:0]),
.flogtanh( I829aa657f0dd13c3fb86baeda8a3b4c8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic66af6c3c0268cfb0e9f0776c4f4e961 = (I44597d694e9c5d29280e503d72a27c8d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I829aa657f0dd13c3fb86baeda8a3b4c8;


Ic3da32f100a43f826b89a492544e7812 Ic49f0cce261191fcfb823e6211dec290 (
.flogtanh_sel( I04a19448c5e75af8021ad02d1a708bb0[flogtanh_SEL-1:0]),
.flogtanh( I1ae4334c32094064c19df0dac77bd03d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia605d14205926b3edc6d1c2f69f70ac0 = (I04a19448c5e75af8021ad02d1a708bb0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1ae4334c32094064c19df0dac77bd03d;


Ic3da32f100a43f826b89a492544e7812 I0087701442769027b7b3a8c5103192e6 (
.flogtanh_sel( I71a3093121c2f19dcd1412b468652fa8[flogtanh_SEL-1:0]),
.flogtanh( I78788f7e0845e4353145012efa04a48c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0071f2168787bd42ab7f2370aed9d0f5 = (I71a3093121c2f19dcd1412b468652fa8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I78788f7e0845e4353145012efa04a48c;


Ic3da32f100a43f826b89a492544e7812 Ib492393f3c242238855217eaa83fdc4c (
.flogtanh_sel( I3ae09c82029c617034fe6aacbe9e94e6[flogtanh_SEL-1:0]),
.flogtanh( I359f3e3bb2a69349f8564466fa81a054),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4936f823841b0ffe32f801f5134c0211 = (I3ae09c82029c617034fe6aacbe9e94e6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I359f3e3bb2a69349f8564466fa81a054;


Ic3da32f100a43f826b89a492544e7812 I752debe043d8a9e578510fc89bd9998a (
.flogtanh_sel( Ie7af6b3b441f910b000a333afad6c76f[flogtanh_SEL-1:0]),
.flogtanh( I7b630e8ac26638fb858dd3b5d2d56385),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5975ef8f6cf53cf2132cdd9d707e7912 = (Ie7af6b3b441f910b000a333afad6c76f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7b630e8ac26638fb858dd3b5d2d56385;


Ic3da32f100a43f826b89a492544e7812 I19cd387db66c16866078925b41b27dea (
.flogtanh_sel( I4d71dfea8407aa5b5cbb991bc4fea963[flogtanh_SEL-1:0]),
.flogtanh( I859bef71501c2f2a994a0cdf8a94b2a7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I954ff0f9ee871a31774a3d786128fa13 = (I4d71dfea8407aa5b5cbb991bc4fea963[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I859bef71501c2f2a994a0cdf8a94b2a7;


Ic3da32f100a43f826b89a492544e7812 I873119ef3a274502f0b23de2c799ef67 (
.flogtanh_sel( I1a082caecc831a90e74674ba35da4183[flogtanh_SEL-1:0]),
.flogtanh( Ib51b9e41161f4273f6469e8965acd7dd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I31f6bbfbbbd4c20d0c5c71663da1d4c1 = (I1a082caecc831a90e74674ba35da4183[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib51b9e41161f4273f6469e8965acd7dd;


Ic3da32f100a43f826b89a492544e7812 I604529a12f6b8f7af57a74230a9acfe0 (
.flogtanh_sel( Iec1de44616a2354a56ab1f681059d4c5[flogtanh_SEL-1:0]),
.flogtanh( I78bb23c008613c0f07f6f85172482296),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1898bc3cc6a8b6f71d65c758d1f08366 = (Iec1de44616a2354a56ab1f681059d4c5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I78bb23c008613c0f07f6f85172482296;


Ic3da32f100a43f826b89a492544e7812 I4bdba4354d579b912c3d65c530e8384a (
.flogtanh_sel( Ie3c2318e64d0e218c3db557404c4aac8[flogtanh_SEL-1:0]),
.flogtanh( I8b883a5bc22b2cde03f4074357be7c88),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If86532f849bd392dbf599eeb2fae0545 = (Ie3c2318e64d0e218c3db557404c4aac8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8b883a5bc22b2cde03f4074357be7c88;


Ic3da32f100a43f826b89a492544e7812 I3f6b44c374283b77ac5d7d44561d61d9 (
.flogtanh_sel( I9a251d50f41e51b1a5cc2475f267e8a0[flogtanh_SEL-1:0]),
.flogtanh( Ic2727e097ffbce70f07fc9f3d9395b54),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia344734d285ac29b53cf401c08a0f987 = (I9a251d50f41e51b1a5cc2475f267e8a0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic2727e097ffbce70f07fc9f3d9395b54;


Ic3da32f100a43f826b89a492544e7812 Ifd307104e75317ef8514819a606451e2 (
.flogtanh_sel( I9b5767a49f7b9dcb8fdaea924835033c[flogtanh_SEL-1:0]),
.flogtanh( I096397439036b0056c979054528ce1fd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I502a8e382aa0881dc86f3c13e0566ca3 = (I9b5767a49f7b9dcb8fdaea924835033c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I096397439036b0056c979054528ce1fd;


Ic3da32f100a43f826b89a492544e7812 I191a16f6aea463947222fb9a48e1a3fa (
.flogtanh_sel( I6ca1e6700a19d03621a193c7240bff54[flogtanh_SEL-1:0]),
.flogtanh( Ifcc83d9007aafdf32acf04f062e008c8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic462cebbfc39190b22d20013259e39eb = (I6ca1e6700a19d03621a193c7240bff54[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifcc83d9007aafdf32acf04f062e008c8;


Ic3da32f100a43f826b89a492544e7812 I4988bbbf0393c477c27e18525478c364 (
.flogtanh_sel( I931c597ff12bffce581f653346202f83[flogtanh_SEL-1:0]),
.flogtanh( I53c01c60f4061d970e4491564ddf88ae),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I385d03def4cfb49f54867687ebd710ed = (I931c597ff12bffce581f653346202f83[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I53c01c60f4061d970e4491564ddf88ae;


Ic3da32f100a43f826b89a492544e7812 I60a6ca074cf6efff523e57ca4f867ff6 (
.flogtanh_sel( Ia3a2c5d59f6340917ca3933c05ba4678[flogtanh_SEL-1:0]),
.flogtanh( I0b4d34aa164c014f9315debd37fa534b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If8aa3ec1b5a4a3c122da82467be917da = (Ia3a2c5d59f6340917ca3933c05ba4678[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0b4d34aa164c014f9315debd37fa534b;


Ic3da32f100a43f826b89a492544e7812 Ic6f94dae8ab3ffffd030554ca80966e4 (
.flogtanh_sel( Ie83d0a8ee5ed214bc7577467748aaa04[flogtanh_SEL-1:0]),
.flogtanh( Iac97aad4ca2c93e387ff0c1340143029),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8daf79a0a2ee1bac7f055af441539fa4 = (Ie83d0a8ee5ed214bc7577467748aaa04[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iac97aad4ca2c93e387ff0c1340143029;


Ic3da32f100a43f826b89a492544e7812 Ia5b53bda226ff5622cd4c13acbc8b845 (
.flogtanh_sel( Iaac29552e5fc65aaf4f0116f917b707c[flogtanh_SEL-1:0]),
.flogtanh( I8b4c2d8a5f2b796029575ecf3b89e2b9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6261e0d339762cb2364421e6b87086cb = (Iaac29552e5fc65aaf4f0116f917b707c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8b4c2d8a5f2b796029575ecf3b89e2b9;


Ic3da32f100a43f826b89a492544e7812 Ib52108acb173b4adb948b41fcb3af6c2 (
.flogtanh_sel( Ie2c8eac7204b98139c03b6fbfff9af36[flogtanh_SEL-1:0]),
.flogtanh( I06dd747316fa36a8dbdbb4ddf011230b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0e2f746715b901feb69f6b3c94f3a828 = (Ie2c8eac7204b98139c03b6fbfff9af36[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I06dd747316fa36a8dbdbb4ddf011230b;


Ic3da32f100a43f826b89a492544e7812 I1ef56e8089070dcc71ce348b42e40479 (
.flogtanh_sel( Ied7fcdaec662cb3c2f89f131986fa102[flogtanh_SEL-1:0]),
.flogtanh( I1594e7dfaedd9e7f5818dc4d639bb663),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7b8da162c08f8aa2ae90522ee1526cf6 = (Ied7fcdaec662cb3c2f89f131986fa102[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1594e7dfaedd9e7f5818dc4d639bb663;


Ic3da32f100a43f826b89a492544e7812 I7af923c3db3b09f9a8e5e140ccb97715 (
.flogtanh_sel( Ib16a17d6430570b45a304d847ee2b11c[flogtanh_SEL-1:0]),
.flogtanh( Ic8111eb95e6b6ab35bcd8e2cafcd0c1e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5e8ecdbb018402b2fbc0049ee44bae8c = (Ib16a17d6430570b45a304d847ee2b11c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic8111eb95e6b6ab35bcd8e2cafcd0c1e;


Ic3da32f100a43f826b89a492544e7812 Ie86223e557b0c75a9379e6d7fa1a110a (
.flogtanh_sel( I42169e454756fe4d1c5f17f2eeb2e091[flogtanh_SEL-1:0]),
.flogtanh( I650b4641d233096a77ae15c8254a29b1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I06d859184884c07a14c83d2f06587ad5 = (I42169e454756fe4d1c5f17f2eeb2e091[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I650b4641d233096a77ae15c8254a29b1;


Ic3da32f100a43f826b89a492544e7812 If194a90e1c4c621b4d73ed6f1d4dc73a (
.flogtanh_sel( I6fde38a3a92e06fa77123e3279813c41[flogtanh_SEL-1:0]),
.flogtanh( Ia905d37c471bdf7258a547be95b85e4f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I79e3e49f57d47231c0fe6aaafdbc57f1 = (I6fde38a3a92e06fa77123e3279813c41[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia905d37c471bdf7258a547be95b85e4f;


Ic3da32f100a43f826b89a492544e7812 Id8ddef8242a2fd0c90aa17d1c4067c3f (
.flogtanh_sel( Id8ee16437e8d6d6da6d37440e04097b6[flogtanh_SEL-1:0]),
.flogtanh( Icfc2b5de1aa36d81de3f163880d48a68),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I12c07042202f66db926861c9ce7c2b25 = (Id8ee16437e8d6d6da6d37440e04097b6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icfc2b5de1aa36d81de3f163880d48a68;


Ic3da32f100a43f826b89a492544e7812 Ib0e06fdc8efc9aa8ceef18c92e84fd92 (
.flogtanh_sel( Ibf249d8e5acced9b064132575f40e001[flogtanh_SEL-1:0]),
.flogtanh( I3c6893d360627cd954db1c20f3c9d319),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9d0fdb45b9e86bd409740e538a690320 = (Ibf249d8e5acced9b064132575f40e001[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3c6893d360627cd954db1c20f3c9d319;


Ic3da32f100a43f826b89a492544e7812 Ie88762487a8c612f90ec8f2b79f85277 (
.flogtanh_sel( I580659084e3d17b48de6b1c66154fcf5[flogtanh_SEL-1:0]),
.flogtanh( Ibc971e0b7ade69365d2c23f30ba0c1ea),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id5fd6f25dc3df22a322434ae3c90dea6 = (I580659084e3d17b48de6b1c66154fcf5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibc971e0b7ade69365d2c23f30ba0c1ea;


Ic3da32f100a43f826b89a492544e7812 I954996c7ec1b22605b47730275c5c824 (
.flogtanh_sel( I7a14e45d43ab77b265501902152c8616[flogtanh_SEL-1:0]),
.flogtanh( I562d9a1676d27c7966d2920bb6be3b38),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id812a8ea2a3b4a912d151be582833fcf = (I7a14e45d43ab77b265501902152c8616[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I562d9a1676d27c7966d2920bb6be3b38;


Ic3da32f100a43f826b89a492544e7812 Id3c3281e8eff9dcdbbeea29df02af90e (
.flogtanh_sel( I81ba868784103e0eb05a44d981d4d666[flogtanh_SEL-1:0]),
.flogtanh( I8aa258f382bea1eb300b006c3083bec1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifd3638d44e1ba2285891fac152dee327 = (I81ba868784103e0eb05a44d981d4d666[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8aa258f382bea1eb300b006c3083bec1;


Ic3da32f100a43f826b89a492544e7812 I453035bf406c20d368ad06352205962b (
.flogtanh_sel( Ic6b88783957cbaf253648a30b22f6b1c[flogtanh_SEL-1:0]),
.flogtanh( Iec0e7232ec94c15d7d50866ad5eb85fb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idd1b6014de2f053554ed09c29bf3e640 = (Ic6b88783957cbaf253648a30b22f6b1c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iec0e7232ec94c15d7d50866ad5eb85fb;


Ic3da32f100a43f826b89a492544e7812 Ie187a264bd0fef2ef08b80bf5508a3a9 (
.flogtanh_sel( I4103c218a85a1d08db5c4f4b5686b2e5[flogtanh_SEL-1:0]),
.flogtanh( I0d252b23e06d25aee4afd84b4c5b4ba9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0d96336eb4d5071d7e1d350e86513b25 = (I4103c218a85a1d08db5c4f4b5686b2e5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0d252b23e06d25aee4afd84b4c5b4ba9;


Ic3da32f100a43f826b89a492544e7812 I0a99b359cf5fa031ceb4e1ff800a2c1d (
.flogtanh_sel( I0e6c0958af503e4a120a49d02a432863[flogtanh_SEL-1:0]),
.flogtanh( I430703cef7ec173f9099c8391132e5c4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I31e5b2cdc3dc571eafa37510076bcc64 = (I0e6c0958af503e4a120a49d02a432863[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I430703cef7ec173f9099c8391132e5c4;


Ic3da32f100a43f826b89a492544e7812 I7fb2497b689287cfbb3585cfba862cd9 (
.flogtanh_sel( I8f76b31e8f15c0e5fe24dcb723418111[flogtanh_SEL-1:0]),
.flogtanh( I5788d966ba8393f5d76dcfcb9294b52e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia8849f78971a45ed0daa2489e7d27dd7 = (I8f76b31e8f15c0e5fe24dcb723418111[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5788d966ba8393f5d76dcfcb9294b52e;


Ic3da32f100a43f826b89a492544e7812 I150a778c3a2a620c105a0af478dc121a (
.flogtanh_sel( Id1457221b58344b60070aa026436df2c[flogtanh_SEL-1:0]),
.flogtanh( Ied561890134d28b451f26da773ea5525),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie4749f8e9ad2b370f9f9814b5a463c43 = (Id1457221b58344b60070aa026436df2c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ied561890134d28b451f26da773ea5525;


Ic3da32f100a43f826b89a492544e7812 I3fc10e51814099b4ebd90fabcd8af525 (
.flogtanh_sel( Icc31966508e03d8869e81d8aeb243705[flogtanh_SEL-1:0]),
.flogtanh( I52e018ad790a1e406777510a0f4b6c29),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3096d11098113da669ee0a94686e600d = (Icc31966508e03d8869e81d8aeb243705[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I52e018ad790a1e406777510a0f4b6c29;


Ic3da32f100a43f826b89a492544e7812 I64daef8db512ef764c759740d316e0a7 (
.flogtanh_sel( I9dcccf542ba434b6e0fde6f012f98f92[flogtanh_SEL-1:0]),
.flogtanh( I25eb66d8589cbb35b32cd25539a24f7f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I09a1d04c307fcb8a0e30925d86df3fe9 = (I9dcccf542ba434b6e0fde6f012f98f92[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I25eb66d8589cbb35b32cd25539a24f7f;


Ic3da32f100a43f826b89a492544e7812 I7e8896a311fdca4590b4b896ae2fab0b (
.flogtanh_sel( I51ccbb824a5e1e340eefd173c4491728[flogtanh_SEL-1:0]),
.flogtanh( Icd4716d0d66d95a532544461c4872d11),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idb0a98cea3ee6cd4308bfc2414a003e1 = (I51ccbb824a5e1e340eefd173c4491728[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icd4716d0d66d95a532544461c4872d11;


Ic3da32f100a43f826b89a492544e7812 I6d846f729b3bd7d15edd7edd18a962c2 (
.flogtanh_sel( Ib7ae1730dcd8bc708bbfcc6a9f97ac66[flogtanh_SEL-1:0]),
.flogtanh( I266ba4229056534d310d982253b5f9b9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id4788855f9a503e8b506d012aaeea445 = (Ib7ae1730dcd8bc708bbfcc6a9f97ac66[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I266ba4229056534d310d982253b5f9b9;


Ic3da32f100a43f826b89a492544e7812 Ice68b02b2aa9080e68fb6a46b61439a7 (
.flogtanh_sel( I4714f5c91203fcfa552f0fcf71b87442[flogtanh_SEL-1:0]),
.flogtanh( I86498c8c820d276ac12764b5df267252),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5b937934e7aae1f916c2848889f12685 = (I4714f5c91203fcfa552f0fcf71b87442[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I86498c8c820d276ac12764b5df267252;


Ic3da32f100a43f826b89a492544e7812 I3c0a3121ae11d7a9ec428add5b080f3c (
.flogtanh_sel( I3b6d1e84fdd1019249886fa5fe65895b[flogtanh_SEL-1:0]),
.flogtanh( I7bb9ad1a2cd32966746b05b7604a09b6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9275bb36e58e0f17964e13ee7f027ab7 = (I3b6d1e84fdd1019249886fa5fe65895b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7bb9ad1a2cd32966746b05b7604a09b6;


Ic3da32f100a43f826b89a492544e7812 I889e113801b481e602307b82f01cbe24 (
.flogtanh_sel( Ia8a7d4207dbabc7970bf36f3fe74f72d[flogtanh_SEL-1:0]),
.flogtanh( Id0998cc2848a6a72ed2701a8e720946e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I02330ade2eed926076cc071e45eed82c = (Ia8a7d4207dbabc7970bf36f3fe74f72d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id0998cc2848a6a72ed2701a8e720946e;


Ic3da32f100a43f826b89a492544e7812 I5edf8bd34ffbb793f1a072b4e21e20ff (
.flogtanh_sel( I84047457b43ef33874f4550c3b773460[flogtanh_SEL-1:0]),
.flogtanh( If1ed051cd94d42e7836f82c10538b302),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I296bc392d4223cbdd6f77be6523df819 = (I84047457b43ef33874f4550c3b773460[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If1ed051cd94d42e7836f82c10538b302;


Ic3da32f100a43f826b89a492544e7812 Ide77db16d85c807676405e55cb72c583 (
.flogtanh_sel( I5e51563c3e69beca0b463742e6e5f9ee[flogtanh_SEL-1:0]),
.flogtanh( I780afd116929565d1ff9b3833ba242d5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I31b0f2fe98cfddbc05dbd14be8be394b = (I5e51563c3e69beca0b463742e6e5f9ee[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I780afd116929565d1ff9b3833ba242d5;


Ic3da32f100a43f826b89a492544e7812 I2fef22b0a3f67a751197c43d12a230d2 (
.flogtanh_sel( I6c8d14e31c80811ccab1b6ab09d28089[flogtanh_SEL-1:0]),
.flogtanh( I89ee99e699676bcec20031b6cad0e2ac),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia71663e8f563041c27cd21a0c9c27a28 = (I6c8d14e31c80811ccab1b6ab09d28089[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I89ee99e699676bcec20031b6cad0e2ac;


Ic3da32f100a43f826b89a492544e7812 I3abd34d32f67155bbb9e76c18a990b48 (
.flogtanh_sel( I50b3b7490c9b65b6e662cc86b163a2df[flogtanh_SEL-1:0]),
.flogtanh( I862b467403c045e4694fb57d59e10064),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib46b13498ec14ceaa56719f26f18febb = (I50b3b7490c9b65b6e662cc86b163a2df[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I862b467403c045e4694fb57d59e10064;


Ic3da32f100a43f826b89a492544e7812 I544cddffa373016b01f6c54c9b89d589 (
.flogtanh_sel( I8351a2110a3d73ad8803cf17e3317017[flogtanh_SEL-1:0]),
.flogtanh( Ic3b554c66f652f027159dbc0fccc5ba3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9bc2d5692474b8368c570d92835191b3 = (I8351a2110a3d73ad8803cf17e3317017[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic3b554c66f652f027159dbc0fccc5ba3;


Ic3da32f100a43f826b89a492544e7812 I868923006897c0c59b3934ee560ee267 (
.flogtanh_sel( I1e6c696951688d581f21ab2302593335[flogtanh_SEL-1:0]),
.flogtanh( I04635713f6d70142b7ab3ecb5ffe6ac9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If8b0b96a659183e3651c691a2848b86b = (I1e6c696951688d581f21ab2302593335[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I04635713f6d70142b7ab3ecb5ffe6ac9;


Ic3da32f100a43f826b89a492544e7812 If8e88f32c9cb4c1f89d416f472c6cb42 (
.flogtanh_sel( Ie9840e28133eebdca0be313552195c7b[flogtanh_SEL-1:0]),
.flogtanh( I1917eae0dbcc0a941718c3248c7d4b11),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I87d958c00fc6209d901147831b0c951c = (Ie9840e28133eebdca0be313552195c7b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1917eae0dbcc0a941718c3248c7d4b11;


Ic3da32f100a43f826b89a492544e7812 I5f9659087b55397213a8e7438f6e31f7 (
.flogtanh_sel( I82812258a8032e273cab7139266be1b6[flogtanh_SEL-1:0]),
.flogtanh( Ifa60c3079164485f31442d9cf12bd2ad),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie4e4eaf3e5d2f581210af8054df71c6c = (I82812258a8032e273cab7139266be1b6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifa60c3079164485f31442d9cf12bd2ad;


Ic3da32f100a43f826b89a492544e7812 I361852ce4f21de3ebde870e8026b17de (
.flogtanh_sel( I27ab6fd9927518e29ed36d7a7a241498[flogtanh_SEL-1:0]),
.flogtanh( I5616405acf49c3e8608ae4d2b544b0d6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0b557cf102da41afd26936cbdb64b6e8 = (I27ab6fd9927518e29ed36d7a7a241498[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5616405acf49c3e8608ae4d2b544b0d6;


Ic3da32f100a43f826b89a492544e7812 Ib27e57de9c87f97e250ec5892c54338a (
.flogtanh_sel( I05b0f33a3808ac53b29d8d8309447650[flogtanh_SEL-1:0]),
.flogtanh( Ie6f9ae463fa1add4de23463435a23d25),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I49eb064043f91112c854e31e4eb9b885 = (I05b0f33a3808ac53b29d8d8309447650[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie6f9ae463fa1add4de23463435a23d25;


Ic3da32f100a43f826b89a492544e7812 I637b750e4ae79f2d0d91b45b3e57277d (
.flogtanh_sel( If150ebf242231f0d22c996a71552f6eb[flogtanh_SEL-1:0]),
.flogtanh( Ib16a67d67a4650e53547312e3af60363),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1039bc43e88eee527d2ed6adb8c7d1ba = (If150ebf242231f0d22c996a71552f6eb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib16a67d67a4650e53547312e3af60363;


Ic3da32f100a43f826b89a492544e7812 I099572371eef8a853a3618de5c6c0b15 (
.flogtanh_sel( If2d0a2b58510715e74787cb60719cb5b[flogtanh_SEL-1:0]),
.flogtanh( I8fa4ad645ca2ef21dea8669d2e2afbe2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9aab16e89f1b64117caece8ca8af5940 = (If2d0a2b58510715e74787cb60719cb5b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8fa4ad645ca2ef21dea8669d2e2afbe2;


Ic3da32f100a43f826b89a492544e7812 I5103ae3e1695e713b5a3439a2def56c1 (
.flogtanh_sel( Ib6745a6d17034a29501e022bd846bf2f[flogtanh_SEL-1:0]),
.flogtanh( I41ea2e3d798ff8e0a95f04e4773c59b4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I343df614f97cf732e57cf2ad3f95dc9e = (Ib6745a6d17034a29501e022bd846bf2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41ea2e3d798ff8e0a95f04e4773c59b4;


Ic3da32f100a43f826b89a492544e7812 I7df444d3b5785dfef2490545e87403c6 (
.flogtanh_sel( Iae09c127dfe86c9f7bdbeff447c777f5[flogtanh_SEL-1:0]),
.flogtanh( Id7f4c6208197cdbf48fecdb2a18b81fc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie02de90d8eb06b16314946d21299500c = (Iae09c127dfe86c9f7bdbeff447c777f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id7f4c6208197cdbf48fecdb2a18b81fc;


Ic3da32f100a43f826b89a492544e7812 I412ac07316c9f52e5f9d927c7feccc6e (
.flogtanh_sel( I742128de6b237ed48e3a7ccd3788f0d7[flogtanh_SEL-1:0]),
.flogtanh( I0adb66417482782dd71da1678c1f7412),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3353a7916b569f2c0ca122180608dccc = (I742128de6b237ed48e3a7ccd3788f0d7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0adb66417482782dd71da1678c1f7412;


Ic3da32f100a43f826b89a492544e7812 If36873ecaf128f8033f9c22c3af060f0 (
.flogtanh_sel( Id5e8fda13ba8f6d95d694d0f30da75bb[flogtanh_SEL-1:0]),
.flogtanh( I2abe89a1366a1ad862266ad88101baa2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibfe760474fcac99f1e5ffa2e008fef99 = (Id5e8fda13ba8f6d95d694d0f30da75bb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2abe89a1366a1ad862266ad88101baa2;


Ic3da32f100a43f826b89a492544e7812 Idc49f18e909ac800f57bd8437a7988ec (
.flogtanh_sel( I1aa5a04e40f9b1685c77e4d101c3ccf4[flogtanh_SEL-1:0]),
.flogtanh( I8d10f0c6dc026005f7882ca013283099),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3caf1211dcbcdc746a3e4c7fbbdae4a8 = (I1aa5a04e40f9b1685c77e4d101c3ccf4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8d10f0c6dc026005f7882ca013283099;


Ic3da32f100a43f826b89a492544e7812 I18714ed2a5ad9652f7d42e3a4733251d (
.flogtanh_sel( Ife1adea26d13bc299bb2de241ad4a6ea[flogtanh_SEL-1:0]),
.flogtanh( I4ef16908ce9b89771f94068eec1a983e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2dcc0d17b9fcac35693bf32b5c5540fd = (Ife1adea26d13bc299bb2de241ad4a6ea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4ef16908ce9b89771f94068eec1a983e;


Ic3da32f100a43f826b89a492544e7812 I1b95a03881d2f23ad2a5efcbf2569cdd (
.flogtanh_sel( Ifcf6c761f0f253921710af87ab1d2247[flogtanh_SEL-1:0]),
.flogtanh( I4f6bcd6e0bcd77730248b69d2b93c904),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie6764a631310e312ba5c2c1e601d828f = (Ifcf6c761f0f253921710af87ab1d2247[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4f6bcd6e0bcd77730248b69d2b93c904;


Ic3da32f100a43f826b89a492544e7812 I6fa8917dae215a86c17655573a6e3cb1 (
.flogtanh_sel( I1478e6a9113c124bdc4361908af6643f[flogtanh_SEL-1:0]),
.flogtanh( Iea1ae39e18f083fb8f855fd9ad3d4f8e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I220f8e45e5fe6e69f02cded87f12e1e5 = (I1478e6a9113c124bdc4361908af6643f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iea1ae39e18f083fb8f855fd9ad3d4f8e;


Ic3da32f100a43f826b89a492544e7812 I3af6f5b66a9a99ecb9b89b2d60ac120f (
.flogtanh_sel( I0afd42151925883835844cf5deef6156[flogtanh_SEL-1:0]),
.flogtanh( I795ae30dec63ef2952917eb3355148a2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I896cd566a3d078b0f697a788efd223f2 = (I0afd42151925883835844cf5deef6156[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I795ae30dec63ef2952917eb3355148a2;


Ic3da32f100a43f826b89a492544e7812 I72979f9f549b7229d29c723980bba7f5 (
.flogtanh_sel( I2b4ab0aadffb3a1bb86f45ebc8acf085[flogtanh_SEL-1:0]),
.flogtanh( I188813c5474bf304b59dbe07c78bef6f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7caa41076a293edf18c7c4309fdcfc91 = (I2b4ab0aadffb3a1bb86f45ebc8acf085[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I188813c5474bf304b59dbe07c78bef6f;


Ic3da32f100a43f826b89a492544e7812 I13a343511d5bf4755a879af1c34fc8ed (
.flogtanh_sel( Iffa867719ba9c31a8756cc5e6bf81147[flogtanh_SEL-1:0]),
.flogtanh( I1760a42d85513ea751e94a8b829b5f1a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I928a0e4951208aab170656596f456209 = (Iffa867719ba9c31a8756cc5e6bf81147[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1760a42d85513ea751e94a8b829b5f1a;


Ic3da32f100a43f826b89a492544e7812 I8edadee2eb2ce40fa390fb24710b75d4 (
.flogtanh_sel( Ibb62b6cb003f0d5549c864075f23d19b[flogtanh_SEL-1:0]),
.flogtanh( I8c652055cfcd230426887e171eaf2511),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia3d129fd297905bee180293c0c39d9ef = (Ibb62b6cb003f0d5549c864075f23d19b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8c652055cfcd230426887e171eaf2511;


Ic3da32f100a43f826b89a492544e7812 I2de6d68b88909d4f19b775e47917b75b (
.flogtanh_sel( I3690d101ae99f258cc58b4482cc378c8[flogtanh_SEL-1:0]),
.flogtanh( I9a88a91b0fcc6dd1a7b4ed24e676d9e1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id555c88cf7f0904db74d45cc75c8f5d6 = (I3690d101ae99f258cc58b4482cc378c8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9a88a91b0fcc6dd1a7b4ed24e676d9e1;


Ic3da32f100a43f826b89a492544e7812 I45a273cb3fc7275abc7a565cbc649855 (
.flogtanh_sel( Id597e95ce8a168ab67890085a26870d0[flogtanh_SEL-1:0]),
.flogtanh( I89f6566e2295d58668e63b9529d94df8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1ddfd31bbf062aa5c3c71d61e492e3a2 = (Id597e95ce8a168ab67890085a26870d0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I89f6566e2295d58668e63b9529d94df8;


Ic3da32f100a43f826b89a492544e7812 Id6b2ce96e394f9990d90980b600460c8 (
.flogtanh_sel( I98df60eb8f65641f9cccce4023be905c[flogtanh_SEL-1:0]),
.flogtanh( I08295c218fd06a8900974edc9c2924f2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iae9e023628eb6686708b2656f15616cc = (I98df60eb8f65641f9cccce4023be905c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I08295c218fd06a8900974edc9c2924f2;


Ic3da32f100a43f826b89a492544e7812 Id7b8820c207d8d3942751014cf3e396b (
.flogtanh_sel( Ibcb4fbdee372353b79c460cdeafdfe4e[flogtanh_SEL-1:0]),
.flogtanh( I0a39fdea8b5bfac1862f199152e26ffe),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If4b100d26126e460c41b8c1bc8fbbb96 = (Ibcb4fbdee372353b79c460cdeafdfe4e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0a39fdea8b5bfac1862f199152e26ffe;


Ic3da32f100a43f826b89a492544e7812 Iceefc682a14ccad2db03fca7c8e642fe (
.flogtanh_sel( I74dbf75966d047a4a9e91c1bc793666f[flogtanh_SEL-1:0]),
.flogtanh( Ib36a71ff310882325be0a2745e48f708),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I85a7fede715578be0634d71e9c7951cd = (I74dbf75966d047a4a9e91c1bc793666f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib36a71ff310882325be0a2745e48f708;


Ic3da32f100a43f826b89a492544e7812 Iccfc8c17cb1e9b04bbd05d30c68ce8b0 (
.flogtanh_sel( I79b8d9f9447c4c1b551ec6c1e8903040[flogtanh_SEL-1:0]),
.flogtanh( I75e4d037cc2ed0b0f75fc1fe9cb21da3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2d7715a3af03d9664729fa6df85034a2 = (I79b8d9f9447c4c1b551ec6c1e8903040[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I75e4d037cc2ed0b0f75fc1fe9cb21da3;


Ic3da32f100a43f826b89a492544e7812 I70b1e8cb0062241b4b53fb479349c4ae (
.flogtanh_sel( Ib34b66548621fabe0753223712b1369f[flogtanh_SEL-1:0]),
.flogtanh( Iee9e9849924642a9579a10655624fa17),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I571ddcb0a10938e4c0816c965214b4a8 = (Ib34b66548621fabe0753223712b1369f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iee9e9849924642a9579a10655624fa17;


Ic3da32f100a43f826b89a492544e7812 I9894896829f7e6b6454cc4937e975b99 (
.flogtanh_sel( Ie5b3eb4c00bedfaecc3215d43ff28362[flogtanh_SEL-1:0]),
.flogtanh( I0a267feb8313c9fa5c663a3fe68284dd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8bf8b0cf27a2654a0e7fdf3255945b67 = (Ie5b3eb4c00bedfaecc3215d43ff28362[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0a267feb8313c9fa5c663a3fe68284dd;


Ic3da32f100a43f826b89a492544e7812 Ia6c85fc15efe23d7c59d2dd588ddff07 (
.flogtanh_sel( Icf3a1b0b6dbcf959b44379024f3c4169[flogtanh_SEL-1:0]),
.flogtanh( I0e0ff3511e65a1dda10ec944c89d09d7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I63f82f075d53205b5b556c0054f1a0b8 = (Icf3a1b0b6dbcf959b44379024f3c4169[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0e0ff3511e65a1dda10ec944c89d09d7;


Ic3da32f100a43f826b89a492544e7812 Id4d710fa03d3e930baf2ae4d7cd0388a (
.flogtanh_sel( I918c2bbe7c71f8c6a07b0bad8811f4e7[flogtanh_SEL-1:0]),
.flogtanh( I4504a0a17633d26163a0afae21ad0f43),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3c6fb0df5846a19228a4e6cf9f9106ac = (I918c2bbe7c71f8c6a07b0bad8811f4e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4504a0a17633d26163a0afae21ad0f43;


Ic3da32f100a43f826b89a492544e7812 I788854048c9db748bb88305142d5de3c (
.flogtanh_sel( Iedd960a21b1c08b4a5293cff200218b3[flogtanh_SEL-1:0]),
.flogtanh( Ibd7b7f4ba86b6c61a0dd38f71c67ae05),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7168b0efdd2fae57292379c9d15c62eb = (Iedd960a21b1c08b4a5293cff200218b3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibd7b7f4ba86b6c61a0dd38f71c67ae05;


Ic3da32f100a43f826b89a492544e7812 Ic7bc684be7299f38971cbd8c2dfb495c (
.flogtanh_sel( If9722c28747df3a59b0ecf8200907e98[flogtanh_SEL-1:0]),
.flogtanh( Icddd184270ffda26b803956883400ad0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibe502ebbb366f54a8f8fda4e361308e3 = (If9722c28747df3a59b0ecf8200907e98[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icddd184270ffda26b803956883400ad0;


Ic3da32f100a43f826b89a492544e7812 Ic487f2b1d45a998959bf6d278969aa9b (
.flogtanh_sel( Ib83df72c8b73a333d0699a8bbbec16be[flogtanh_SEL-1:0]),
.flogtanh( Id3da7061c05091ffc520d4480058e8e9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifce70fefde8f5ea4d2c1857236f66d65 = (Ib83df72c8b73a333d0699a8bbbec16be[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id3da7061c05091ffc520d4480058e8e9;


Ic3da32f100a43f826b89a492544e7812 Ie9af7acffee6de1eb96634b24d9f13a2 (
.flogtanh_sel( Ide3798a77f709a9f694523338b081f70[flogtanh_SEL-1:0]),
.flogtanh( Ie63d649228270b34d8ed25e7c4b09883),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice2c390d296e09b117d60905343e9098 = (Ide3798a77f709a9f694523338b081f70[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie63d649228270b34d8ed25e7c4b09883;


Ic3da32f100a43f826b89a492544e7812 Iacab793a98e6b438a0b250dfa775296b (
.flogtanh_sel( I0a9722a805604433562f85c62b168b96[flogtanh_SEL-1:0]),
.flogtanh( I8eed3f7b36c046fff1e41dd52a300d29),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4b94402a53d981e953c21ef316c709b7 = (I0a9722a805604433562f85c62b168b96[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8eed3f7b36c046fff1e41dd52a300d29;


Ic3da32f100a43f826b89a492544e7812 I2deed88b7f179b7dc0a41ddc90019c22 (
.flogtanh_sel( If9480ec13cd538ed03a43e56bd6264a6[flogtanh_SEL-1:0]),
.flogtanh( Iefcebe38e0c2d6d570017e165d70d3b1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I450c0d6ad5d3b1f18bb28e3a432b5442 = (If9480ec13cd538ed03a43e56bd6264a6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iefcebe38e0c2d6d570017e165d70d3b1;


Ic3da32f100a43f826b89a492544e7812 I68dd079497d998561260a755b82dc3fa (
.flogtanh_sel( I433ecf86b7704c5552e5fb5cafe0d529[flogtanh_SEL-1:0]),
.flogtanh( Ia153222350357443978d7426663c3eaa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2587a5800a5a9ffeabc4dca503e3d964 = (I433ecf86b7704c5552e5fb5cafe0d529[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia153222350357443978d7426663c3eaa;


Ic3da32f100a43f826b89a492544e7812 Ib3967ce8b1f89fdd3114782355b14377 (
.flogtanh_sel( I8326f0b2d25139609e2c5e466724f224[flogtanh_SEL-1:0]),
.flogtanh( I06f0fd2d9d46a2fdb4221217ee2496d1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1182655739d7ab5bbe4a6546a5ca36fd = (I8326f0b2d25139609e2c5e466724f224[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I06f0fd2d9d46a2fdb4221217ee2496d1;


Ic3da32f100a43f826b89a492544e7812 Ife592791cd5e41d80eb7d9eb77270cb1 (
.flogtanh_sel( Ibbe211d9955cdf2810c9003d1fb78074[flogtanh_SEL-1:0]),
.flogtanh( I9533ff0882ed01409795d7269329fd76),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8110a5a62607093b21b7cd088b1d9ee0 = (Ibbe211d9955cdf2810c9003d1fb78074[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9533ff0882ed01409795d7269329fd76;


Ic3da32f100a43f826b89a492544e7812 I5e7adcb3ed1429927a76a244d2527d69 (
.flogtanh_sel( If15e950b569a92b590127d0ca6f20a16[flogtanh_SEL-1:0]),
.flogtanh( Ia9eb9821e7dc31c23d7e60839949c1ff),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8b611f7c12ddd81de403ba74e212857f = (If15e950b569a92b590127d0ca6f20a16[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia9eb9821e7dc31c23d7e60839949c1ff;


Ic3da32f100a43f826b89a492544e7812 I1edc59047920506549ace5959da95ce5 (
.flogtanh_sel( I03e0532841ba39eb1d4ae823c4de2f7d[flogtanh_SEL-1:0]),
.flogtanh( I3663fc86620d6244a850819bd3ebe72c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I84a62a133dbceb5a32a7c907f371663d = (I03e0532841ba39eb1d4ae823c4de2f7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3663fc86620d6244a850819bd3ebe72c;


Ic3da32f100a43f826b89a492544e7812 Iac037e6522d597b13d321532915df713 (
.flogtanh_sel( I1be81a7b73987ee023e396cec87312d1[flogtanh_SEL-1:0]),
.flogtanh( I11293e7cdeddf352011d46abd6c3bb72),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia2fc8a1bbc3cb0dd7d89a7f05b04909c = (I1be81a7b73987ee023e396cec87312d1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I11293e7cdeddf352011d46abd6c3bb72;


Ic3da32f100a43f826b89a492544e7812 I5768df3b7be6734f8d1caf13d5240321 (
.flogtanh_sel( I4ce1a767a78673590c4074f3f03bad8d[flogtanh_SEL-1:0]),
.flogtanh( Ic9339e415d0f756e34bcd930de63ad87),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2a3eb42a4402e873d081f94a14a99c20 = (I4ce1a767a78673590c4074f3f03bad8d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic9339e415d0f756e34bcd930de63ad87;


Ic3da32f100a43f826b89a492544e7812 I6d771fb02e713cfc4bf7929f466cea18 (
.flogtanh_sel( I57806bb7da625881e68ae315543f70d6[flogtanh_SEL-1:0]),
.flogtanh( Icf109f65e24d3a23ecad9e7d4cc54dc1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I58447d6ae49a6be2d043477a06f83df0 = (I57806bb7da625881e68ae315543f70d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icf109f65e24d3a23ecad9e7d4cc54dc1;


Ic3da32f100a43f826b89a492544e7812 Ic9d658321948865c46728be562b7f6e5 (
.flogtanh_sel( I8b0ab476b4790150575abb06bcdce2b3[flogtanh_SEL-1:0]),
.flogtanh( Idf7dd0ff83b2d56693e729a1a375fabb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I83292bcda4645233d8e8a1dfe8e5f60b = (I8b0ab476b4790150575abb06bcdce2b3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idf7dd0ff83b2d56693e729a1a375fabb;


Ic3da32f100a43f826b89a492544e7812 Ie2f5f74057b157c17dfa7ac49c834399 (
.flogtanh_sel( I8846a8961b7d557df4fc62dada679c33[flogtanh_SEL-1:0]),
.flogtanh( I312a248019372261c0959cdc9378ec93),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic5e0a84cf1a2ef907b2456559ea26c75 = (I8846a8961b7d557df4fc62dada679c33[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I312a248019372261c0959cdc9378ec93;


Ic3da32f100a43f826b89a492544e7812 I0589c76d81ca182d7be41b4803590154 (
.flogtanh_sel( I7909a0f96a92e93f95023cddc742a5eb[flogtanh_SEL-1:0]),
.flogtanh( I8e311b9891dda272762da2c640019e8c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2cefbf897bb7f6f67ca500727e85c683 = (I7909a0f96a92e93f95023cddc742a5eb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8e311b9891dda272762da2c640019e8c;


Ic3da32f100a43f826b89a492544e7812 Id0ec5ecfff5e14158a26024268ceb744 (
.flogtanh_sel( I43ac4857544c0fb79d04e850435ef673[flogtanh_SEL-1:0]),
.flogtanh( I1874dd9f7c0a93310873173561402912),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If47be2ca4617a426258c51f8d977ba3f = (I43ac4857544c0fb79d04e850435ef673[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1874dd9f7c0a93310873173561402912;


Ic3da32f100a43f826b89a492544e7812 If6ebd2295760a0536ad245a16f8430be (
.flogtanh_sel( Ia6dfa47c465325c1d9fb9b9c5ce08f01[flogtanh_SEL-1:0]),
.flogtanh( I04adb3964e739a106098a6c4d2f49e94),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7c68e0ae30efc4ca4d68b6047119c6c3 = (Ia6dfa47c465325c1d9fb9b9c5ce08f01[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I04adb3964e739a106098a6c4d2f49e94;


Ic3da32f100a43f826b89a492544e7812 I398652d5ace1fbbcae9c343935f133a2 (
.flogtanh_sel( I2e9eda5bea0cc3d88359ce8a7a82f21f[flogtanh_SEL-1:0]),
.flogtanh( I9135b709c3c802a42c7186087b5664cc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iccca1936f4c1c9496205e77b588e9985 = (I2e9eda5bea0cc3d88359ce8a7a82f21f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9135b709c3c802a42c7186087b5664cc;


Ic3da32f100a43f826b89a492544e7812 I5580ab45adaac9d7872faec2063c6301 (
.flogtanh_sel( I53ec2486418e41b2ccfa8fd82777eaf0[flogtanh_SEL-1:0]),
.flogtanh( Ia236dfe34ff4938456d76f787d2db945),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I59d4567d3355fdae5660a1364d1b8d00 = (I53ec2486418e41b2ccfa8fd82777eaf0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia236dfe34ff4938456d76f787d2db945;


Ic3da32f100a43f826b89a492544e7812 Icd58ab459e5144889f6b44c545b17dea (
.flogtanh_sel( I18387c05cef21970ecbc39c20a87aafb[flogtanh_SEL-1:0]),
.flogtanh( I41c98bae5fbdb31bac0913930573e80c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4600963866dcb9bbea2515c805f885cb = (I18387c05cef21970ecbc39c20a87aafb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41c98bae5fbdb31bac0913930573e80c;


Ic3da32f100a43f826b89a492544e7812 I71ee711d784840d722a1c99c9756ebb7 (
.flogtanh_sel( I2b23eae78cb925008ad59f45e80e165b[flogtanh_SEL-1:0]),
.flogtanh( I226befd72285893998aca87fe34d9aaf),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If26d90629e70c5a871e6f5b14471b8cf = (I2b23eae78cb925008ad59f45e80e165b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I226befd72285893998aca87fe34d9aaf;


Ic3da32f100a43f826b89a492544e7812 I53ac521d87e8564003f755f0f40d2a34 (
.flogtanh_sel( Ic69eb7677638a90b7a54389d47be46de[flogtanh_SEL-1:0]),
.flogtanh( I20ab7c6174af39aee99492f704b2748c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iedb9bb14951bf67bc8865b0983490c14 = (Ic69eb7677638a90b7a54389d47be46de[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I20ab7c6174af39aee99492f704b2748c;


Ic3da32f100a43f826b89a492544e7812 Ife82bce13890ef71870777fcaabd7328 (
.flogtanh_sel( I8cb9a216f4da7c27f678386cb214c59d[flogtanh_SEL-1:0]),
.flogtanh( I0a1c5724ffa14df653142a1f8bcf44a4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6a3854ed571e8c262aa3ec377c247778 = (I8cb9a216f4da7c27f678386cb214c59d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0a1c5724ffa14df653142a1f8bcf44a4;


Ic3da32f100a43f826b89a492544e7812 I902a7c06c049f3a0bf00e617b039782e (
.flogtanh_sel( I48cb720a6323697084ac3bbd8fcadfcb[flogtanh_SEL-1:0]),
.flogtanh( I481973954b81accf069dd80830fba3bc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I05028975b49ec0c089bd981696f85a8b = (I48cb720a6323697084ac3bbd8fcadfcb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I481973954b81accf069dd80830fba3bc;


Ic3da32f100a43f826b89a492544e7812 I771f015e478d35df6c17e7aba6c0c2be (
.flogtanh_sel( Ib8dc3c1885c92cdcce7fcb58d65d03e7[flogtanh_SEL-1:0]),
.flogtanh( Ia6825c3edc9d2a6832db7a7d684faf98),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ife732309efcc740cfff5c747aab2e3d6 = (Ib8dc3c1885c92cdcce7fcb58d65d03e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia6825c3edc9d2a6832db7a7d684faf98;


Ic3da32f100a43f826b89a492544e7812 I7dc3d63e6dd55aff3cb0682ea4c4262c (
.flogtanh_sel( Ic3aa51a5c758405fa6e2dbed707555b2[flogtanh_SEL-1:0]),
.flogtanh( I5c964036207f47629302e282d56fef7b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idcef10a0465614cf38e0d6f503b5174a = (Ic3aa51a5c758405fa6e2dbed707555b2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5c964036207f47629302e282d56fef7b;


Ic3da32f100a43f826b89a492544e7812 I26eab18d515ed85631102b8d6118f52c (
.flogtanh_sel( I4d418179c859feb8bc7d750416bb1004[flogtanh_SEL-1:0]),
.flogtanh( I00b74ed4d6730b37c6fbfd42dee42584),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibd4aaf02982068ffbfd1b8b3795d9217 = (I4d418179c859feb8bc7d750416bb1004[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I00b74ed4d6730b37c6fbfd42dee42584;


Ic3da32f100a43f826b89a492544e7812 I2805a2c28f51eb01e4a3ac38f589649b (
.flogtanh_sel( If207b2adc6f668f85cb76bf54673fe18[flogtanh_SEL-1:0]),
.flogtanh( I0345fc4a507f9e3be3e1d46b71693de1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I788c64785b992c675fe348a1fa181525 = (If207b2adc6f668f85cb76bf54673fe18[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0345fc4a507f9e3be3e1d46b71693de1;


Ic3da32f100a43f826b89a492544e7812 I4d3994b2adacfc7dfb4dab2832c79006 (
.flogtanh_sel( Ib08b8067ea75e210e83526ca4a37217e[flogtanh_SEL-1:0]),
.flogtanh( I9f0735c1cf5d1af7c82a251ef4886f9c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib235af5b28d56f24372d3f0af816f2c2 = (Ib08b8067ea75e210e83526ca4a37217e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9f0735c1cf5d1af7c82a251ef4886f9c;


Ic3da32f100a43f826b89a492544e7812 I51d662becc68b93ec29d4a5653e112b2 (
.flogtanh_sel( I95b30f641cbf7bec1886643c4468017d[flogtanh_SEL-1:0]),
.flogtanh( I861cf5dffb18c84953013dc4026bd08a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4c03a6569d1b954d088053e38827e811 = (I95b30f641cbf7bec1886643c4468017d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I861cf5dffb18c84953013dc4026bd08a;


Ic3da32f100a43f826b89a492544e7812 I25d2a0e341a013a5ceed9a901a1abc32 (
.flogtanh_sel( I1978531a6f8d1d25ee6d404025ec4753[flogtanh_SEL-1:0]),
.flogtanh( I19722ceada71cc9cc06edde39142ff17),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idda26504e422367082caeafbb29871f9 = (I1978531a6f8d1d25ee6d404025ec4753[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I19722ceada71cc9cc06edde39142ff17;


Ic3da32f100a43f826b89a492544e7812 I07ac8362dbacc6edced4066157a81b30 (
.flogtanh_sel( I6c9698ba88db16b8d22ccebd58cc541d[flogtanh_SEL-1:0]),
.flogtanh( Id8349128e2c391df008828494da928c6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I195c3a82123142d509886ee37dc6fc98 = (I6c9698ba88db16b8d22ccebd58cc541d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id8349128e2c391df008828494da928c6;


Ic3da32f100a43f826b89a492544e7812 Id20751b5b475f62b5b63511b4619263e (
.flogtanh_sel( I0d8ac5e09b200a55bf5ba6f834cc9174[flogtanh_SEL-1:0]),
.flogtanh( I27209805df490a07f1726875a7b69922),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1abb512ca0383c9e7104418e07281841 = (I0d8ac5e09b200a55bf5ba6f834cc9174[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I27209805df490a07f1726875a7b69922;


Ic3da32f100a43f826b89a492544e7812 I89ee2b86dd74bf6052337b196a6998ec (
.flogtanh_sel( Ib58b7d3d77a54ff1a180c6fa5f1400e6[flogtanh_SEL-1:0]),
.flogtanh( I7532c1f0624a2d5a94321c89c73e38df),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I00ff1331b1900bb031ee81d2a58c1bd5 = (Ib58b7d3d77a54ff1a180c6fa5f1400e6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7532c1f0624a2d5a94321c89c73e38df;


Ic3da32f100a43f826b89a492544e7812 I554c8e771ba4596299971e3b434cfaae (
.flogtanh_sel( Icf6b990098b7ab91800bfcf1e643153c[flogtanh_SEL-1:0]),
.flogtanh( Ife892846e66e2522c06b170811a11ada),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If65eb5e743a7b1878fb232ef2fe13cb0 = (Icf6b990098b7ab91800bfcf1e643153c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ife892846e66e2522c06b170811a11ada;


Ic3da32f100a43f826b89a492544e7812 I5689239e01c4c9ff9ec7faefd9b47e0e (
.flogtanh_sel( Ie4308b9ac6fb6de9329ba02b1eeb0e8a[flogtanh_SEL-1:0]),
.flogtanh( Ib905ede2830f7e3c8cf993075f07345c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I24ae7de3549a84f4f88f561b6017b7a8 = (Ie4308b9ac6fb6de9329ba02b1eeb0e8a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib905ede2830f7e3c8cf993075f07345c;


Ic3da32f100a43f826b89a492544e7812 Ia62426cb98358c486613704e158e9a10 (
.flogtanh_sel( I01d4f02a356c51d7e4e1993de0d8eebd[flogtanh_SEL-1:0]),
.flogtanh( Ibf169f844d9e00eca8f3821ddc952ef0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I449c77140475475b138d839a74078337 = (I01d4f02a356c51d7e4e1993de0d8eebd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibf169f844d9e00eca8f3821ddc952ef0;


Ic3da32f100a43f826b89a492544e7812 Iadb3a9c38fb173e837e0eba8272858fa (
.flogtanh_sel( I36c351e3641b01cc43e1dd5de0a649e5[flogtanh_SEL-1:0]),
.flogtanh( I3137f75629e72f78abdac088e18608d5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia9e102d8679943c079f16c0228f0f0d1 = (I36c351e3641b01cc43e1dd5de0a649e5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3137f75629e72f78abdac088e18608d5;


Ic3da32f100a43f826b89a492544e7812 I3e3abeb5aa8eabbe133c5aa74b96cc41 (
.flogtanh_sel( I4fc983e94c5b8f7bafca61fb0d351c08[flogtanh_SEL-1:0]),
.flogtanh( I8fbcabc2f5c30fcf1c5b46de5dfe887d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibf1c9d86665f696d91c554db748ff42b = (I4fc983e94c5b8f7bafca61fb0d351c08[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8fbcabc2f5c30fcf1c5b46de5dfe887d;


Ic3da32f100a43f826b89a492544e7812 Ied1a943823b3662e58652c459fb5f589 (
.flogtanh_sel( I1fcb82fdf96cda14a55fa6358cb62c1e[flogtanh_SEL-1:0]),
.flogtanh( Ie7acfb624aa6242b558481350c85fda3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieb0336a1974a2aec0966f4f59f460802 = (I1fcb82fdf96cda14a55fa6358cb62c1e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie7acfb624aa6242b558481350c85fda3;


Ic3da32f100a43f826b89a492544e7812 Id9c9cec648944074216cbcc0fad50c84 (
.flogtanh_sel( I665e54ea6bdca483149d3b7f3ee42a2b[flogtanh_SEL-1:0]),
.flogtanh( I11e0b915338d5d649c800455b9a7695f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic0819ccefe784a6379716b3633ae0196 = (I665e54ea6bdca483149d3b7f3ee42a2b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I11e0b915338d5d649c800455b9a7695f;


Ic3da32f100a43f826b89a492544e7812 Iba327dc6674a5c45a4f569679a095ab3 (
.flogtanh_sel( I925df2307b5af6d1b166e5435641d3bd[flogtanh_SEL-1:0]),
.flogtanh( Ia9e4e68dcd3d0281decde939eed0c3bd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0c4bbd1827b1859caabb067e864ce4b3 = (I925df2307b5af6d1b166e5435641d3bd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia9e4e68dcd3d0281decde939eed0c3bd;


Ic3da32f100a43f826b89a492544e7812 I6469111b19d850549b05e8ddf2687a24 (
.flogtanh_sel( I9b14f48aa357d09e460a445da86cdf89[flogtanh_SEL-1:0]),
.flogtanh( Id508f63a381fc565a28fe4e662b33efb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I004c98da87996b77b5761d366210f782 = (I9b14f48aa357d09e460a445da86cdf89[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id508f63a381fc565a28fe4e662b33efb;


Ic3da32f100a43f826b89a492544e7812 I7f338f3b782de1a3986a9ee0a724aa22 (
.flogtanh_sel( I78e94ecb6c92fa8ee24edaff33b6f82d[flogtanh_SEL-1:0]),
.flogtanh( I33582dc83370e68b0ae7b22b553276b4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia457938da4efe847cb06f645f2a54a52 = (I78e94ecb6c92fa8ee24edaff33b6f82d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I33582dc83370e68b0ae7b22b553276b4;


Ic3da32f100a43f826b89a492544e7812 I15cfeea64b61228a248d1de64c0141ff (
.flogtanh_sel( I5ebeb9ce5adee72a7c9527ea6d3a3028[flogtanh_SEL-1:0]),
.flogtanh( I8aeca996ad6820edcc6fcbaa8a0f15ce),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7e0474089ebc1c34747be1bc17a81d72 = (I5ebeb9ce5adee72a7c9527ea6d3a3028[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8aeca996ad6820edcc6fcbaa8a0f15ce;


Ic3da32f100a43f826b89a492544e7812 I09a1588018f0d894d61c7c14003b89a6 (
.flogtanh_sel( I90d7b28ec09142ca8086836fc0c5ea0d[flogtanh_SEL-1:0]),
.flogtanh( Ica86e8037319b868c8cb89f3cb02b136),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib0b46b99e61d724ae664d9d1fec1e29f = (I90d7b28ec09142ca8086836fc0c5ea0d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ica86e8037319b868c8cb89f3cb02b136;


Ic3da32f100a43f826b89a492544e7812 Iccf9e114b4d5025a5b8afb458103ff19 (
.flogtanh_sel( I27d9985415e6d0b117e5a4c2863aa7f8[flogtanh_SEL-1:0]),
.flogtanh( Ia95013b19d9fc12d19ff9924007113d4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I56d1025271f1f7704a40dd7f0df02b0b = (I27d9985415e6d0b117e5a4c2863aa7f8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia95013b19d9fc12d19ff9924007113d4;


Ic3da32f100a43f826b89a492544e7812 Idb28cb6a9327327e5f957e388fd05a71 (
.flogtanh_sel( Idf9b563e5d10c2bdbcc07e81d74467eb[flogtanh_SEL-1:0]),
.flogtanh( Ifcf979b713b014f22c1c8ce1d42132c2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I72c2256ba47cf03f95143df8f741fd83 = (Idf9b563e5d10c2bdbcc07e81d74467eb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifcf979b713b014f22c1c8ce1d42132c2;


Ic3da32f100a43f826b89a492544e7812 I7324e5bb447f4337582fa0086dd5ca7b (
.flogtanh_sel( Ie351922194483938302ff6cafc477e4a[flogtanh_SEL-1:0]),
.flogtanh( I973b3306021532f286cf248084398c26),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I733c3fa4d84e5680792b16a70bb1a51d = (Ie351922194483938302ff6cafc477e4a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I973b3306021532f286cf248084398c26;


Ic3da32f100a43f826b89a492544e7812 I32a42430f75f148cd3dd2b5bb8997498 (
.flogtanh_sel( Ifb2da5faf236ca8636677bc1dc35c4db[flogtanh_SEL-1:0]),
.flogtanh( Iea7940bb396d1a436f56806fc533edee),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If367d63311c96726517240de13bd2a4b = (Ifb2da5faf236ca8636677bc1dc35c4db[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iea7940bb396d1a436f56806fc533edee;


Ic3da32f100a43f826b89a492544e7812 I766c2db7e949837f12d18c93aa6648b2 (
.flogtanh_sel( Ie15825d216685ae241b528fa9c158ff3[flogtanh_SEL-1:0]),
.flogtanh( Ied55045b003302c294591a8d2a6a39fd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icc6d895d943e14f2801c22e79ce190e8 = (Ie15825d216685ae241b528fa9c158ff3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ied55045b003302c294591a8d2a6a39fd;


Ic3da32f100a43f826b89a492544e7812 Id2386ff2b294a3f4e9803d984171349c (
.flogtanh_sel( Id92c2d8bc61245c0c8e40bec2424c3c8[flogtanh_SEL-1:0]),
.flogtanh( Ib64e948413d5dce1d9309fe95c0919ab),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieb664ac9be65fba2e25960141f7fb4b6 = (Id92c2d8bc61245c0c8e40bec2424c3c8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib64e948413d5dce1d9309fe95c0919ab;


Ic3da32f100a43f826b89a492544e7812 I7964fa1ce64fd652015522deb8728091 (
.flogtanh_sel( Icd9fd8d7114b6e894dbee493b6797df6[flogtanh_SEL-1:0]),
.flogtanh( I682fe6c6c621db5dd867574e8573d8ed),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I66071f20991b414140869a2e3b750471 = (Icd9fd8d7114b6e894dbee493b6797df6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I682fe6c6c621db5dd867574e8573d8ed;


Ic3da32f100a43f826b89a492544e7812 I65bcf5f3157a35f102555eccbd26a341 (
.flogtanh_sel( I29ff688c085f2b18e7a3af969f18af76[flogtanh_SEL-1:0]),
.flogtanh( I508b57f6ebc45eb70aa7b114096a7d12),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iffeefa89a2ba7d032db5db64cbf05e20 = (I29ff688c085f2b18e7a3af969f18af76[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I508b57f6ebc45eb70aa7b114096a7d12;


Ic3da32f100a43f826b89a492544e7812 I9119e7640366214578b9fd7c79af8561 (
.flogtanh_sel( I6d56db9fcfe69dfcd747521a1ff62297[flogtanh_SEL-1:0]),
.flogtanh( I8e82b8914260669ed1d88a690467a7b4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9ab3cea6ee8d8473221da21bae06066b = (I6d56db9fcfe69dfcd747521a1ff62297[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8e82b8914260669ed1d88a690467a7b4;


Ic3da32f100a43f826b89a492544e7812 Iad61cc3f07670a7faa2718fe03c6ea73 (
.flogtanh_sel( I2f17f7c79a0118b39a63894917c6affa[flogtanh_SEL-1:0]),
.flogtanh( I525feb94b558fb4bb8db8eead9f05afa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3403ce6e697b523a9f441d8fd5e2d420 = (I2f17f7c79a0118b39a63894917c6affa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I525feb94b558fb4bb8db8eead9f05afa;


Ic3da32f100a43f826b89a492544e7812 Ief318368d992d8c255649de3ba14d9e4 (
.flogtanh_sel( I7350af5d5ee09ad28c459e3674a829ab[flogtanh_SEL-1:0]),
.flogtanh( Ie5e4cf2b42054822a9091f5ef67cd968),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia98a70144e466b356d2998948dc4b602 = (I7350af5d5ee09ad28c459e3674a829ab[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie5e4cf2b42054822a9091f5ef67cd968;


Ic3da32f100a43f826b89a492544e7812 I81eacd051031fdc622878857cdc7a4d5 (
.flogtanh_sel( I67b6415c5135e3d6a41d56d98d3f8315[flogtanh_SEL-1:0]),
.flogtanh( I0d08d26e31c8b69ed8c089cdcd055a50),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie4ca0836695d951ee09622892ee35928 = (I67b6415c5135e3d6a41d56d98d3f8315[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0d08d26e31c8b69ed8c089cdcd055a50;


Ic3da32f100a43f826b89a492544e7812 I588de0617014fb8432bf5bf26901c7b3 (
.flogtanh_sel( I4a6fffd8bb7244599383f2aa3a1c8916[flogtanh_SEL-1:0]),
.flogtanh( I877f44c880a781381bfa8a8f8471d697),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I485a48b4ff4da08f977425fd10e6d392 = (I4a6fffd8bb7244599383f2aa3a1c8916[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I877f44c880a781381bfa8a8f8471d697;


Ic3da32f100a43f826b89a492544e7812 Ic051a5f98debf78822778d3c7510c4c8 (
.flogtanh_sel( I7dbcd21016231546b76aab175cac9f74[flogtanh_SEL-1:0]),
.flogtanh( I7fc78273dc765cf1c03b3c1a043b35f8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie8c79e6a5378808c0ead5a4b24319ce9 = (I7dbcd21016231546b76aab175cac9f74[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7fc78273dc765cf1c03b3c1a043b35f8;


Ic3da32f100a43f826b89a492544e7812 I4bd2826194e6ec3b098dae91b88c4e97 (
.flogtanh_sel( I9aeff3dc44ed0d0f32518590a900dcc9[flogtanh_SEL-1:0]),
.flogtanh( Ie67275a4b3fdc050f0f6e7ac7d1eebfc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9ca81c841a75a9ac242835956509e0fe = (I9aeff3dc44ed0d0f32518590a900dcc9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie67275a4b3fdc050f0f6e7ac7d1eebfc;


Ic3da32f100a43f826b89a492544e7812 I93de51261c003913fd304c99bd84a8c1 (
.flogtanh_sel( I988b7d5d56d22d2c77c5c8c125129a50[flogtanh_SEL-1:0]),
.flogtanh( I41f9acc96650353174155a5f378d5cc5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id50f18f642f3b00ffa34986f78a0eae6 = (I988b7d5d56d22d2c77c5c8c125129a50[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41f9acc96650353174155a5f378d5cc5;


Ic3da32f100a43f826b89a492544e7812 I25d4b99b5a3cd798a33034ff312f1fa8 (
.flogtanh_sel( Iff35cd97f2a6d37a7861b9cc1a655ef5[flogtanh_SEL-1:0]),
.flogtanh( I0d73c905b2ed777acd71d560928dcf0b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I75838ca09e301b8e1301cbf603a1f8c2 = (Iff35cd97f2a6d37a7861b9cc1a655ef5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0d73c905b2ed777acd71d560928dcf0b;


Ic3da32f100a43f826b89a492544e7812 I42533b9a42dd5381e666ff145dd05c40 (
.flogtanh_sel( Ifb3f2a1bedfe41c73d198046a2a3f177[flogtanh_SEL-1:0]),
.flogtanh( I2b6b1c25caf8b00d19ccc98156a8ca2b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id968b34075e351ab01d65abcb4ed8cca = (Ifb3f2a1bedfe41c73d198046a2a3f177[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2b6b1c25caf8b00d19ccc98156a8ca2b;


Ic3da32f100a43f826b89a492544e7812 I7b4b0ba0f46c4232b9b092443921a095 (
.flogtanh_sel( I37ddc6ccbc188a3eb8c33a501de820be[flogtanh_SEL-1:0]),
.flogtanh( I28ea2b207bcd3518a85ff150466a6a08),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I84da4ce7441e132e775167c1cd81dbe5 = (I37ddc6ccbc188a3eb8c33a501de820be[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I28ea2b207bcd3518a85ff150466a6a08;


Ic3da32f100a43f826b89a492544e7812 I35a3bb68a517dc6bb869bd634c361967 (
.flogtanh_sel( Ica608f1136da397e2ab61bd4a5d83201[flogtanh_SEL-1:0]),
.flogtanh( I7d0a1c64b2e85e1bf0bf99423321466b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If19dc22d45cc4664c85a043ec4c00617 = (Ica608f1136da397e2ab61bd4a5d83201[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7d0a1c64b2e85e1bf0bf99423321466b;


Ic3da32f100a43f826b89a492544e7812 I3d20646f5683308fffafd4f21ca6b946 (
.flogtanh_sel( I80636a3df4541bf29780bcb4d0ee48f9[flogtanh_SEL-1:0]),
.flogtanh( I3b9b9b41b54ff194314b572a15daf606),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibf482db0f5058be72061267c42ebc292 = (I80636a3df4541bf29780bcb4d0ee48f9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3b9b9b41b54ff194314b572a15daf606;


Ic3da32f100a43f826b89a492544e7812 Id532485b1bd48873a9696f01318a6e47 (
.flogtanh_sel( I9ad99d544187db3cc7090b92c9933a31[flogtanh_SEL-1:0]),
.flogtanh( Ic914f847e623d9c52e2d9ae5076c21c3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6d2dbb953a58b91dafa7f0d34d41bdc3 = (I9ad99d544187db3cc7090b92c9933a31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic914f847e623d9c52e2d9ae5076c21c3;


Ic3da32f100a43f826b89a492544e7812 I066535c63c22185e258cc43ecf60574b (
.flogtanh_sel( Iaa8a2b6fcd469869efcf0b75ca38e68f[flogtanh_SEL-1:0]),
.flogtanh( I46fc20938dd554b23b5af5f7c3e39480),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib393146d81d3cf031466543311cee2ad = (Iaa8a2b6fcd469869efcf0b75ca38e68f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I46fc20938dd554b23b5af5f7c3e39480;


Ic3da32f100a43f826b89a492544e7812 I4c85b76161932951c3e304c6c3e1c8cd (
.flogtanh_sel( I9a171d2d8eee362a0073ab7b139d3037[flogtanh_SEL-1:0]),
.flogtanh( I1fa8b37b4697ae60cf399285d9524b8d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I42564ec6a794ea803795f0b5b3523a93 = (I9a171d2d8eee362a0073ab7b139d3037[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1fa8b37b4697ae60cf399285d9524b8d;


Ic3da32f100a43f826b89a492544e7812 I998b8a7b4239c02de65776c266aa158b (
.flogtanh_sel( I84cdcba86bc5991feb391003cd7be40b[flogtanh_SEL-1:0]),
.flogtanh( I66c8261df769288836e188ecb32b6dc6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4a0033a180d7edce81fcfef603532e28 = (I84cdcba86bc5991feb391003cd7be40b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I66c8261df769288836e188ecb32b6dc6;


Ic3da32f100a43f826b89a492544e7812 I120ff224dcc3a4ed4e9c87f87b4f60a7 (
.flogtanh_sel( If9e5c3a848acce5daf570458f78f6aad[flogtanh_SEL-1:0]),
.flogtanh( I267714c8a5aa14bae9c74da272a60aa5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic7a21921e2716fba55aad2e351f4498a = (If9e5c3a848acce5daf570458f78f6aad[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I267714c8a5aa14bae9c74da272a60aa5;


Ic3da32f100a43f826b89a492544e7812 I1bf5df75ac3e874444f05c422cd46219 (
.flogtanh_sel( I73247d4348333f67a491fc607b15af0e[flogtanh_SEL-1:0]),
.flogtanh( I47a34c8d2174c12f96041e82ad835db2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9a3f0b4867087790c78f674b719dbf7b = (I73247d4348333f67a491fc607b15af0e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I47a34c8d2174c12f96041e82ad835db2;


Ic3da32f100a43f826b89a492544e7812 I742ea019a0dd217b84ee013b3c166ab3 (
.flogtanh_sel( I021c745eee4b85a2cd91d9d8d2b18b2c[flogtanh_SEL-1:0]),
.flogtanh( If99ca487495a015063fd8dc54ae596aa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I138f008a6206a1067bb0e22ce3d90990 = (I021c745eee4b85a2cd91d9d8d2b18b2c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If99ca487495a015063fd8dc54ae596aa;


Ic3da32f100a43f826b89a492544e7812 I987c7e10b6a42e17b9a7c50bef1ccc61 (
.flogtanh_sel( I1381c0a0bd28b1c5542992084635b355[flogtanh_SEL-1:0]),
.flogtanh( I1043f1b92b49a8c304a23c0b5c615def),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I48ad9b737892d7c49340ed679f46e034 = (I1381c0a0bd28b1c5542992084635b355[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1043f1b92b49a8c304a23c0b5c615def;


Ic3da32f100a43f826b89a492544e7812 Ifb2bf39243945ac599d6994b1a6e8055 (
.flogtanh_sel( Ie74eeddc21428254a8fc4c3e293b5eb7[flogtanh_SEL-1:0]),
.flogtanh( Icafa102383ef33455236ba268b1b7460),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I04a9c9765fd468a7e841577f09fc287b = (Ie74eeddc21428254a8fc4c3e293b5eb7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icafa102383ef33455236ba268b1b7460;


Ic3da32f100a43f826b89a492544e7812 I34e160be46791b4d21848c5f2090cd10 (
.flogtanh_sel( Ib1d0f94258b45de4bfe610086d8990c5[flogtanh_SEL-1:0]),
.flogtanh( I677fca8017154fed3e6cd54362e829db),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7b929c228c865112f00bc6b4dcc95b52 = (Ib1d0f94258b45de4bfe610086d8990c5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I677fca8017154fed3e6cd54362e829db;


Ic3da32f100a43f826b89a492544e7812 I0c878da4bc007d57a9f77fe262ca5ffc (
.flogtanh_sel( I138d6d5d60df37870cdbb1d9c51a94af[flogtanh_SEL-1:0]),
.flogtanh( I826fe051a6b09d5cacf712431ce89b7c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2b54a135e59945901e9c11580a29ee3d = (I138d6d5d60df37870cdbb1d9c51a94af[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I826fe051a6b09d5cacf712431ce89b7c;


Ic3da32f100a43f826b89a492544e7812 Id9d543bc9a9601676f98cb4d50127304 (
.flogtanh_sel( I706378735e63e15c8d5395446ea41db8[flogtanh_SEL-1:0]),
.flogtanh( I23f781ebfa449cec7975b94179d72259),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I566221060f06e724676ec9bec861d7de = (I706378735e63e15c8d5395446ea41db8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I23f781ebfa449cec7975b94179d72259;


Ic3da32f100a43f826b89a492544e7812 Iffe64346beb2561305131e02f57eeae3 (
.flogtanh_sel( If8680a7fc4f5532a660006bf4ca6a66e[flogtanh_SEL-1:0]),
.flogtanh( Ia383b5dc3b7ce1bc7987926535639668),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icd9a876a0feb16ea62bcad5be2004dac = (If8680a7fc4f5532a660006bf4ca6a66e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia383b5dc3b7ce1bc7987926535639668;


Ic3da32f100a43f826b89a492544e7812 I497cdc03af4fb0d3546ad3f57b1b07f9 (
.flogtanh_sel( Ic59d1ff3051a95166c3c2d5a2881221b[flogtanh_SEL-1:0]),
.flogtanh( I40ae857caffae41564c2ecb0c7e9777b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8f8273c4cb2a9ace8a09847efd4bdec7 = (Ic59d1ff3051a95166c3c2d5a2881221b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I40ae857caffae41564c2ecb0c7e9777b;


Ic3da32f100a43f826b89a492544e7812 I93eb1eb39d8011cd1dad9ccfa1796dba (
.flogtanh_sel( I54a551af28c505601cdfaf8faaa94afb[flogtanh_SEL-1:0]),
.flogtanh( I569d56a2673a104f3050d851d767af8a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I96ef4b631a7f63e19f67f3920685f0e6 = (I54a551af28c505601cdfaf8faaa94afb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I569d56a2673a104f3050d851d767af8a;


Ic3da32f100a43f826b89a492544e7812 I92d07fa26c11e6f1421c67de23603976 (
.flogtanh_sel( I6a3124c03eb83d41c16704133bd1cfde[flogtanh_SEL-1:0]),
.flogtanh( I2022005072d2979dae84b6e4491a3ce2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9e2de71442b8f504358e582087a6d19f = (I6a3124c03eb83d41c16704133bd1cfde[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2022005072d2979dae84b6e4491a3ce2;


Ic3da32f100a43f826b89a492544e7812 I6343f2f05c746c228383c3fe533b1439 (
.flogtanh_sel( Ie9ee27b9761af611ab96f0010abd47a3[flogtanh_SEL-1:0]),
.flogtanh( I98524ad028e4d832ebbcd92956dac08c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1fb13d7500f5ac3821c424bd3688cf4e = (Ie9ee27b9761af611ab96f0010abd47a3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I98524ad028e4d832ebbcd92956dac08c;


Ic3da32f100a43f826b89a492544e7812 I602773c88e41bb06fe19399941e842c4 (
.flogtanh_sel( I305436919f84066a22ab1417ebabd737[flogtanh_SEL-1:0]),
.flogtanh( I4d24e2ba47093eee6669f537374ecce7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2aabda12ff89e708d04b4399472b5203 = (I305436919f84066a22ab1417ebabd737[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4d24e2ba47093eee6669f537374ecce7;


Ic3da32f100a43f826b89a492544e7812 Ia1dc8afcceac6a6e161adee409e6214b (
.flogtanh_sel( I78e63717f436493b756efa32d66cdefd[flogtanh_SEL-1:0]),
.flogtanh( I227232e7189020459c16b3413e881b80),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8c733a5d394e6b8d045eede5cc7451f6 = (I78e63717f436493b756efa32d66cdefd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I227232e7189020459c16b3413e881b80;


Ic3da32f100a43f826b89a492544e7812 I5ddfcb36c35d03af44f019f352a1b420 (
.flogtanh_sel( Ic965ba971642db19ca773eb68dc0b9bf[flogtanh_SEL-1:0]),
.flogtanh( If4359aebd4cc66c75cf2a44f681ccc72),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4f45dd50d2825ab338b8a2a8264096c0 = (Ic965ba971642db19ca773eb68dc0b9bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If4359aebd4cc66c75cf2a44f681ccc72;


Ic3da32f100a43f826b89a492544e7812 I4f33dfb8a61f65531a495883eb135fe6 (
.flogtanh_sel( I579480a66a5f6331fb46de13090ce888[flogtanh_SEL-1:0]),
.flogtanh( I8d2e10b8c474f1a915825ec78072ad56),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib45caf6b563d22144be3e9225a99a1cd = (I579480a66a5f6331fb46de13090ce888[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8d2e10b8c474f1a915825ec78072ad56;


Ic3da32f100a43f826b89a492544e7812 I68e15e60a73f03a40c416ade83f75c05 (
.flogtanh_sel( I38d78b447217271a63f30f78b424e2ae[flogtanh_SEL-1:0]),
.flogtanh( Ie5b3748f3c81d9eeec767d546b29cbd8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9d6730140c690037b5ca58aa30103f5b = (I38d78b447217271a63f30f78b424e2ae[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie5b3748f3c81d9eeec767d546b29cbd8;


Ic3da32f100a43f826b89a492544e7812 Ide128e81c2e631105ca0b5651a08f58d (
.flogtanh_sel( I4c8d7e5474b19a7c63444d0cb6143728[flogtanh_SEL-1:0]),
.flogtanh( Ib764a6d1978dc61cb4499b15c45cb1b4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9df5b63f66c162d517daa69f5d0e6095 = (I4c8d7e5474b19a7c63444d0cb6143728[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib764a6d1978dc61cb4499b15c45cb1b4;


Ic3da32f100a43f826b89a492544e7812 Iab10286ef2d840325576e235813295a9 (
.flogtanh_sel( Ia4bc4b7414bf31305ec8f63e7eda61e7[flogtanh_SEL-1:0]),
.flogtanh( I4fbe7db2d4288676183dc69ed56c9c68),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1b40adfd6fa6c943dfa8d230d9e65514 = (Ia4bc4b7414bf31305ec8f63e7eda61e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4fbe7db2d4288676183dc69ed56c9c68;


Ic3da32f100a43f826b89a492544e7812 I2b08883ac8edaf243d1c789c7077a16b (
.flogtanh_sel( Ibbebe287d56c7d627f3ffcf706575e77[flogtanh_SEL-1:0]),
.flogtanh( I99f0cc5986099cb57fbebf9e5e262c56),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0eb3df4d4094e09e6c4b3c788baed61f = (Ibbebe287d56c7d627f3ffcf706575e77[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I99f0cc5986099cb57fbebf9e5e262c56;


Ic3da32f100a43f826b89a492544e7812 I36de683cc30dd15bd0e7bee30ceeece7 (
.flogtanh_sel( I83867e6ee369fff7e39ef5c8d5398fef[flogtanh_SEL-1:0]),
.flogtanh( I4f5bb7e206563a334d7e2dd100b37c35),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id6f7923a16cc5adc96a730083153ca6d = (I83867e6ee369fff7e39ef5c8d5398fef[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4f5bb7e206563a334d7e2dd100b37c35;


Ic3da32f100a43f826b89a492544e7812 I1c88ba6df8a727790c8e0b00c2b738a6 (
.flogtanh_sel( I1d40df7dbf99674f987bd06db714a702[flogtanh_SEL-1:0]),
.flogtanh( I59ecb14b5f34ebab3da4784709de66a4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idf8ebc0d747ae143aa61866e33d458c0 = (I1d40df7dbf99674f987bd06db714a702[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I59ecb14b5f34ebab3da4784709de66a4;


Ic3da32f100a43f826b89a492544e7812 I87bb8679b6fb1fe2d6bf9252edf3dbea (
.flogtanh_sel( I92f42789cb81760ff2973e3a5fe915c3[flogtanh_SEL-1:0]),
.flogtanh( I54f5a8caf0e1c2df9477b37157d94995),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id682e531735437bc24abbf3d3d51e18b = (I92f42789cb81760ff2973e3a5fe915c3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I54f5a8caf0e1c2df9477b37157d94995;


Ic3da32f100a43f826b89a492544e7812 I325e2fdd785ee73b7b21b81231c7e0d3 (
.flogtanh_sel( Idbd5f2a25ab05808721cf9c403017565[flogtanh_SEL-1:0]),
.flogtanh( I77e1bed2da0ccf1475dcfe908d64f82c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I05ecce409cca00ea5b0df25de5a50cf2 = (Idbd5f2a25ab05808721cf9c403017565[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I77e1bed2da0ccf1475dcfe908d64f82c;


Ic3da32f100a43f826b89a492544e7812 I2c51c458a95acd7982eba2ae9f785493 (
.flogtanh_sel( I7ca5f07d6d3c2a045dfd55ae5214dd65[flogtanh_SEL-1:0]),
.flogtanh( I1a450ec193ccde2946f6ca20c0fa894c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I831d214dcb4f8d534b5ddaaeaeeb81ce = (I7ca5f07d6d3c2a045dfd55ae5214dd65[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1a450ec193ccde2946f6ca20c0fa894c;


Ic3da32f100a43f826b89a492544e7812 Ib02168d6dba7e0fca55580b2958516b8 (
.flogtanh_sel( I7f4e1445c68abbadce23944b99d206f9[flogtanh_SEL-1:0]),
.flogtanh( I01fbfc3b5c14733738f93a3487e54f35),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia540866403683bc30504bace19bdda7b = (I7f4e1445c68abbadce23944b99d206f9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I01fbfc3b5c14733738f93a3487e54f35;


Ic3da32f100a43f826b89a492544e7812 I15ad3388c6707f20b81099dc66348dc9 (
.flogtanh_sel( Id9f28016678e5e2127d9f0aa93e0b534[flogtanh_SEL-1:0]),
.flogtanh( Icff5d12020f78478c77210d9c692dfbe),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I05fb1982415bd3fa78dd9a00af7a3d4a = (Id9f28016678e5e2127d9f0aa93e0b534[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icff5d12020f78478c77210d9c692dfbe;


Ic3da32f100a43f826b89a492544e7812 I1c9006b4914bfe480d90983e7a7a55f4 (
.flogtanh_sel( I6b939c57a8b7c7c51ab43e1b1df12f6a[flogtanh_SEL-1:0]),
.flogtanh( I6eb28698ab4105a74c6510dbcfefbc3c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I977864efb0d94149cce7dc4d165f11de = (I6b939c57a8b7c7c51ab43e1b1df12f6a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6eb28698ab4105a74c6510dbcfefbc3c;


Ic3da32f100a43f826b89a492544e7812 I5cd46b41fb2b8cac2f693e5d3934d624 (
.flogtanh_sel( Ic5d0df586d56bf4cb322d4c3ad677385[flogtanh_SEL-1:0]),
.flogtanh( I7cc0f835ad7a18683e1fdb5bcbfb7f2f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9362b615a612599239e3b752a9334e8c = (Ic5d0df586d56bf4cb322d4c3ad677385[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7cc0f835ad7a18683e1fdb5bcbfb7f2f;


Ic3da32f100a43f826b89a492544e7812 If93135a28738e973e39e4d9ba9bfe549 (
.flogtanh_sel( I2e287724873cf6761799eaf464ed6302[flogtanh_SEL-1:0]),
.flogtanh( I9389a0dfe5a82a903c89e1a468f0ad57),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5d4fb4b5a5ad3dc48beebfa0e0cebbed = (I2e287724873cf6761799eaf464ed6302[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9389a0dfe5a82a903c89e1a468f0ad57;


Ic3da32f100a43f826b89a492544e7812 I0cea1aa59bacb04d36583b0f52a0bb2c (
.flogtanh_sel( Ia7a10cffe31a53aafa1104b97543280b[flogtanh_SEL-1:0]),
.flogtanh( Idc4ce4afd846e212526d21a5e0cd1c14),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifb9b29c43f435452cc761218c509f5df = (Ia7a10cffe31a53aafa1104b97543280b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idc4ce4afd846e212526d21a5e0cd1c14;


Ic3da32f100a43f826b89a492544e7812 I8f084479560c53da76219cc04b326d8b (
.flogtanh_sel( Ieeb089c6a18791a2227c8571913d689a[flogtanh_SEL-1:0]),
.flogtanh( I38a0ba1e69b467d4aed306e76ec3bfdb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If2143db72bf9a02b64eb45b3a4faa39d = (Ieeb089c6a18791a2227c8571913d689a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I38a0ba1e69b467d4aed306e76ec3bfdb;


Ic3da32f100a43f826b89a492544e7812 I9c6f1545dddecedcce8b8bf0e63ed432 (
.flogtanh_sel( Ib29b00328971c3cd67209a5ea5b63b0a[flogtanh_SEL-1:0]),
.flogtanh( I66279b0fa707a272f43ee929cb297945),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice780b1695a8e80607a03dee3c426ffe = (Ib29b00328971c3cd67209a5ea5b63b0a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I66279b0fa707a272f43ee929cb297945;


Ic3da32f100a43f826b89a492544e7812 I48d1d5fc3d471b54863f783d505a611b (
.flogtanh_sel( I517e0868f2bb9a22c287a1f3eeaad2f3[flogtanh_SEL-1:0]),
.flogtanh( Ib091954846c14743e01fd4e7bafda1b5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I90b0296f5ef87dfaa6110fc2e9d6ed9d = (I517e0868f2bb9a22c287a1f3eeaad2f3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib091954846c14743e01fd4e7bafda1b5;


Ic3da32f100a43f826b89a492544e7812 Ifc5e96f6d55cd4077e745f594632ac03 (
.flogtanh_sel( I2bc9f76469e2a3f9846560ad1975cf54[flogtanh_SEL-1:0]),
.flogtanh( I3b8663f2adecb8da2c84dbb37341e25f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icd37da8ea84a606529e32b2db4eb7f5f = (I2bc9f76469e2a3f9846560ad1975cf54[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3b8663f2adecb8da2c84dbb37341e25f;


Ic3da32f100a43f826b89a492544e7812 Iad978a09c0cf77c2833cca261956e66b (
.flogtanh_sel( I9f089315e435cd69d2929fdd936a8a77[flogtanh_SEL-1:0]),
.flogtanh( I19bc03089c6c288e1778bd1f197a3ce3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie626a24e3680f7d3995dd0c2ce60cbcc = (I9f089315e435cd69d2929fdd936a8a77[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I19bc03089c6c288e1778bd1f197a3ce3;


Ic3da32f100a43f826b89a492544e7812 I9012b9f20a606e72d00a3b7e8d63ab29 (
.flogtanh_sel( I9b54c9fb4179423c731217286e329930[flogtanh_SEL-1:0]),
.flogtanh( I0988382a446b21da209d49d0d00bd6df),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iebee55168fb47664095b11c9f6641124 = (I9b54c9fb4179423c731217286e329930[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0988382a446b21da209d49d0d00bd6df;


Ic3da32f100a43f826b89a492544e7812 Ic40dae9287348c46281920f4da0f01e8 (
.flogtanh_sel( I82fb41ab743146badfd2e82258afb310[flogtanh_SEL-1:0]),
.flogtanh( I19f5cb50b27b6c5e40012df9397aa288),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic0954671eb1dc893c3932e456800fadf = (I82fb41ab743146badfd2e82258afb310[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I19f5cb50b27b6c5e40012df9397aa288;


Ic3da32f100a43f826b89a492544e7812 Ic18d2f208631a4085f42a264080f3ffb (
.flogtanh_sel( I5619b91de99eead78befdcba1c62411e[flogtanh_SEL-1:0]),
.flogtanh( I706ca74386e5778b30eca35432429bc3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia4131464996aabab8aae1db85f6a50e4 = (I5619b91de99eead78befdcba1c62411e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I706ca74386e5778b30eca35432429bc3;


Ic3da32f100a43f826b89a492544e7812 Id9815b8b85433860f62acef909eae612 (
.flogtanh_sel( I83dd2047dece99cd841b2e7955819d57[flogtanh_SEL-1:0]),
.flogtanh( If6af0cc7a120b2897c3a69d54a554e86),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2de1ca2c390bdd3011fff4a359bb5332 = (I83dd2047dece99cd841b2e7955819d57[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If6af0cc7a120b2897c3a69d54a554e86;


Ic3da32f100a43f826b89a492544e7812 I6940ba6624872e10fea51a9e6cd53c84 (
.flogtanh_sel( I8c927e66ccbf4d19f07af5ef9fbfe3fb[flogtanh_SEL-1:0]),
.flogtanh( I88ebe846173f486b07d2051a80bd055f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6fb55222b69475b7168874423226ec9c = (I8c927e66ccbf4d19f07af5ef9fbfe3fb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I88ebe846173f486b07d2051a80bd055f;


Ic3da32f100a43f826b89a492544e7812 I72be6a96d5bde170dea9299599eaf0d2 (
.flogtanh_sel( I0793fa8938acdf65486e5582d01b9e5a[flogtanh_SEL-1:0]),
.flogtanh( I2c577b130db6f4673704c858d454f3ea),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9b09b800a9dcd8ac36f25cb0324e748d = (I0793fa8938acdf65486e5582d01b9e5a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2c577b130db6f4673704c858d454f3ea;


Ic3da32f100a43f826b89a492544e7812 I4001e2462b038b65b179127689b9af00 (
.flogtanh_sel( Ied68d7ba0ee9974eb33767e737760b4d[flogtanh_SEL-1:0]),
.flogtanh( I383f23d4e769bbdc1c8acd9c660a0b3e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I74ac0327175f50f508a5013df298df02 = (Ied68d7ba0ee9974eb33767e737760b4d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I383f23d4e769bbdc1c8acd9c660a0b3e;


Ic3da32f100a43f826b89a492544e7812 I54ef2322948ea1e0a279176aa8ad9bb4 (
.flogtanh_sel( I95ba37056659b29fd4318a68d85445e8[flogtanh_SEL-1:0]),
.flogtanh( Iea20a6ecf4bbf907d1a102bde797284f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ica26f542586d50c56ce0f3c00f36b388 = (I95ba37056659b29fd4318a68d85445e8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iea20a6ecf4bbf907d1a102bde797284f;


Ic3da32f100a43f826b89a492544e7812 I50b15718c2d4920e806970e65b88e56e (
.flogtanh_sel( I08d7051a18f358d08728f1c401c15c47[flogtanh_SEL-1:0]),
.flogtanh( I77d655383c0c22b1af75d9308fab2e4f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7c6862830daffc98cb2c1fc121d82c38 = (I08d7051a18f358d08728f1c401c15c47[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I77d655383c0c22b1af75d9308fab2e4f;


Ic3da32f100a43f826b89a492544e7812 I765de144c4e405d975e573fb33e38fad (
.flogtanh_sel( I768b6f55827ac49eb6ac2655e9397be1[flogtanh_SEL-1:0]),
.flogtanh( I4a4ebb2f3389d67c4b7671e12fc5cd92),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icf19dd665616a8c96146b3ab9f46c741 = (I768b6f55827ac49eb6ac2655e9397be1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4a4ebb2f3389d67c4b7671e12fc5cd92;


Ic3da32f100a43f826b89a492544e7812 I121fe3dea1c412926e20e406ed9e35ad (
.flogtanh_sel( Ic66f737fe60c55d4c10e5d72b307a061[flogtanh_SEL-1:0]),
.flogtanh( Ibc927d678e218397e23147b5c0654fd9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I97f2813ec39bbf1513faf66b3e38838a = (Ic66f737fe60c55d4c10e5d72b307a061[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibc927d678e218397e23147b5c0654fd9;


Ic3da32f100a43f826b89a492544e7812 I82b2e7546a321545f51e1aa934de55a2 (
.flogtanh_sel( I5653779f15c6c9b0f3b26927c48d6234[flogtanh_SEL-1:0]),
.flogtanh( Ib0358b6f47edcd54971935de215203f8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I716ee53e79883f69aa045380a357e913 = (I5653779f15c6c9b0f3b26927c48d6234[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib0358b6f47edcd54971935de215203f8;


Ic3da32f100a43f826b89a492544e7812 I7c34f9c887442ebc58a33045e284a8c9 (
.flogtanh_sel( Iac550729fc437fd67151fab57134ec88[flogtanh_SEL-1:0]),
.flogtanh( Iaa6f2bbd8a343ebf878da57badb4572b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I25c324feaca84e80f58075597e8c448f = (Iac550729fc437fd67151fab57134ec88[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaa6f2bbd8a343ebf878da57badb4572b;


Ic3da32f100a43f826b89a492544e7812 I95e98963cb4dfba642e84a8e416bb722 (
.flogtanh_sel( I853b03c5826eedc3c67a2fae7a640212[flogtanh_SEL-1:0]),
.flogtanh( I823f1a0d2d757d5ca83dc7b5ca08e0f8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7fc190647082a3d71614f46f670167bc = (I853b03c5826eedc3c67a2fae7a640212[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I823f1a0d2d757d5ca83dc7b5ca08e0f8;


Ic3da32f100a43f826b89a492544e7812 Ie1735ed691e4c4bdab20970aa3c9e487 (
.flogtanh_sel( If46a6b47c1c52243cc0bc92d1edb594f[flogtanh_SEL-1:0]),
.flogtanh( I1a650234a61a3ff90ea079e29d322069),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iebdf938a28594624f4d4a337356485cb = (If46a6b47c1c52243cc0bc92d1edb594f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1a650234a61a3ff90ea079e29d322069;


Ic3da32f100a43f826b89a492544e7812 If928be4a9c6f2e8b73a7da5a7bf34f49 (
.flogtanh_sel( I75b36a9b429cd657afc8151b9613aca6[flogtanh_SEL-1:0]),
.flogtanh( I70a7b1083c9593840759854430ee9d62),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3fd068d55154441ffd005999ea823fd0 = (I75b36a9b429cd657afc8151b9613aca6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I70a7b1083c9593840759854430ee9d62;


Ic3da32f100a43f826b89a492544e7812 I01ec4c83564dc147544f89f98ad95196 (
.flogtanh_sel( Ife682dd9f677da4d27294fb61b141948[flogtanh_SEL-1:0]),
.flogtanh( I99aa55a3e285e62e9a8b50174e84b68c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic5ca74b66763c6e5591c7c2bfeeb0663 = (Ife682dd9f677da4d27294fb61b141948[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I99aa55a3e285e62e9a8b50174e84b68c;


Ic3da32f100a43f826b89a492544e7812 Ia792bc5779ef305ad9c4a0c6d1ea01d1 (
.flogtanh_sel( Ic2b6177a9c586b274b68b25584e6df2c[flogtanh_SEL-1:0]),
.flogtanh( Ief099d2084b84e0e23599d98102a13b7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5ab556386d2973354a5551ba9823e4ba = (Ic2b6177a9c586b274b68b25584e6df2c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ief099d2084b84e0e23599d98102a13b7;


Ic3da32f100a43f826b89a492544e7812 I552c5629b3d0039e678cd25449a22551 (
.flogtanh_sel( I0d23011c4381496a19cced7bf7960546[flogtanh_SEL-1:0]),
.flogtanh( I84aa89bab681c2fc7a8c7c6b47200dec),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I64f65df774d29696425ba460dda09b68 = (I0d23011c4381496a19cced7bf7960546[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I84aa89bab681c2fc7a8c7c6b47200dec;


Ic3da32f100a43f826b89a492544e7812 Ia85d999d97c6100b4044cf7bf69e549e (
.flogtanh_sel( Ic5992d5eaeafd5dded641a7d9801e763[flogtanh_SEL-1:0]),
.flogtanh( I101b9397639b59fd53a88d17425e0c96),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9e09c25be9f877c1e1aaf79bf12c7943 = (Ic5992d5eaeafd5dded641a7d9801e763[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I101b9397639b59fd53a88d17425e0c96;


Ic3da32f100a43f826b89a492544e7812 I67134d40050d977d9d0a419d080a963a (
.flogtanh_sel( Ic9e7fe68b9045c6c9eb86185b5f5872e[flogtanh_SEL-1:0]),
.flogtanh( Ic302f050dba883d8f4bd20b1030ba14d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I42c1d469ff97913cbf15e3ebee6fdfa8 = (Ic9e7fe68b9045c6c9eb86185b5f5872e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic302f050dba883d8f4bd20b1030ba14d;


Ic3da32f100a43f826b89a492544e7812 I6b2093ed3fcd637becbdf92f71b0d255 (
.flogtanh_sel( I51ad746720b5e6e09ab50f0283552f1a[flogtanh_SEL-1:0]),
.flogtanh( I848425f041888d7433b68900f259732a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If9f2a53dbf6e9b9a335a7657b7a2b468 = (I51ad746720b5e6e09ab50f0283552f1a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I848425f041888d7433b68900f259732a;


Ic3da32f100a43f826b89a492544e7812 I7b55d36fb01e3fa4e01f7b734fe73b80 (
.flogtanh_sel( I0c8964888a1315507f5d71959dd24cf0[flogtanh_SEL-1:0]),
.flogtanh( I2b4671193178503f5329954e74a399b3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I495f8be463b15db906474c518e0741e2 = (I0c8964888a1315507f5d71959dd24cf0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2b4671193178503f5329954e74a399b3;


Ic3da32f100a43f826b89a492544e7812 Ic9f654621fe49ace3022d80a05650ff5 (
.flogtanh_sel( Id4d4f814a0bb3418cbf70c306acf048f[flogtanh_SEL-1:0]),
.flogtanh( I97b93c6d963d51a819b1dc9ab3bf28ea),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3e265a7dcf29687248b9275df49771fb = (Id4d4f814a0bb3418cbf70c306acf048f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I97b93c6d963d51a819b1dc9ab3bf28ea;


Ic3da32f100a43f826b89a492544e7812 I6be204c36c2ea0b1ac868a142e06b3ef (
.flogtanh_sel( Ic91bd7b4bd148e526ca21d4a5ba87be9[flogtanh_SEL-1:0]),
.flogtanh( I2593b1b30f4c97845a1f77c3f558b263),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iffd94cf3a8a4681ff3327c90bf89bd8b = (Ic91bd7b4bd148e526ca21d4a5ba87be9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2593b1b30f4c97845a1f77c3f558b263;


Ic3da32f100a43f826b89a492544e7812 I1ce3a48699f634292542bfa5146bd075 (
.flogtanh_sel( I7959dddc32f0f181b3ba39149afe1016[flogtanh_SEL-1:0]),
.flogtanh( I3a4695c79b62f6baa47cdc939c4e2974),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iea71417e738c6ca54c50aa014cc38627 = (I7959dddc32f0f181b3ba39149afe1016[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3a4695c79b62f6baa47cdc939c4e2974;


Ic3da32f100a43f826b89a492544e7812 I5f7d70dcbdbb154ce7d84cdc8a4716fd (
.flogtanh_sel( I087263600b5f38be072a4f1db787aea7[flogtanh_SEL-1:0]),
.flogtanh( Ibc577b2948aec87c0696c860d7efa1d7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic8df04756f67e6dd29f3374c5f86d451 = (I087263600b5f38be072a4f1db787aea7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibc577b2948aec87c0696c860d7efa1d7;


Ic3da32f100a43f826b89a492544e7812 Icdd9b114d49efbbe685ad9d6123ead43 (
.flogtanh_sel( I78d17a56de5cbe08191ef23b9731c485[flogtanh_SEL-1:0]),
.flogtanh( I08401e4e9a1766a0034f45933b5bb29a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I546122346a22ad64a6ab2b4978cde095 = (I78d17a56de5cbe08191ef23b9731c485[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I08401e4e9a1766a0034f45933b5bb29a;


Ic3da32f100a43f826b89a492544e7812 Id275849e3670b109fed780738dde5063 (
.flogtanh_sel( I82f713a43596df3b935d6da6f8041dc2[flogtanh_SEL-1:0]),
.flogtanh( I5e5bb0de4fe6682a6beaa86f6cd1ca32),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icaae0fb0f460f68d690ab00697355a49 = (I82f713a43596df3b935d6da6f8041dc2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5e5bb0de4fe6682a6beaa86f6cd1ca32;


Ic3da32f100a43f826b89a492544e7812 Iaeffb06cb0480028cc417d05e4075aaa (
.flogtanh_sel( I422987396853a6a39dabb6e7ddbf91fb[flogtanh_SEL-1:0]),
.flogtanh( Ia487e80f0010e7cb34aa12471e62a62f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I42455e7e4d0c63f97702d204d18a446e = (I422987396853a6a39dabb6e7ddbf91fb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia487e80f0010e7cb34aa12471e62a62f;


Ic3da32f100a43f826b89a492544e7812 I3eb86409ea46b9e06d4d5b451e75fa8f (
.flogtanh_sel( Ibb6556671e104141dd33188ea5fc024d[flogtanh_SEL-1:0]),
.flogtanh( I3bee9305e2f4456aae800bbb174b7843),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaec2f15665e83416bc140890f3cdde9a = (Ibb6556671e104141dd33188ea5fc024d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3bee9305e2f4456aae800bbb174b7843;


Ic3da32f100a43f826b89a492544e7812 If924bd06ddd4705e62497d0e279abe2b (
.flogtanh_sel( Ie42ce76076a2a5e887e0112086012da6[flogtanh_SEL-1:0]),
.flogtanh( I14f1aa0dbf6f1f0fbf6b5f996e229a04),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I487391402b6aa27bf212724a37ea9c33 = (Ie42ce76076a2a5e887e0112086012da6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I14f1aa0dbf6f1f0fbf6b5f996e229a04;


Ic3da32f100a43f826b89a492544e7812 I990d855e86abded668d588f68fa51e03 (
.flogtanh_sel( I4aea430599b9c0702b3bebd5960b5c91[flogtanh_SEL-1:0]),
.flogtanh( If87afc1cf342dca9986f798c38a69dab),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia9f375709014a9d553d46cff2799b59f = (I4aea430599b9c0702b3bebd5960b5c91[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If87afc1cf342dca9986f798c38a69dab;


Ic3da32f100a43f826b89a492544e7812 I9016b3cc58ad66529907803e873f64a3 (
.flogtanh_sel( Icbe11a3970136e485eee1bc5053e7273[flogtanh_SEL-1:0]),
.flogtanh( Ibb1c020ea255a966e54c00fc7cc745b5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I34d428a56bd0142a9be9f627f1c3c87f = (Icbe11a3970136e485eee1bc5053e7273[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibb1c020ea255a966e54c00fc7cc745b5;


Ic3da32f100a43f826b89a492544e7812 I0fe7f64845563025b0777948ab4d3f58 (
.flogtanh_sel( I0a7f1ea1719c1f5ff104445a4130a5a8[flogtanh_SEL-1:0]),
.flogtanh( Icae8a2980dd7403caf72820ae508885b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I57db98eb439d59a895dabe029c6a3a8b = (I0a7f1ea1719c1f5ff104445a4130a5a8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icae8a2980dd7403caf72820ae508885b;


Ic3da32f100a43f826b89a492544e7812 I55b424cc9358d653f64c09db0c0b84e9 (
.flogtanh_sel( I1802d759f26dd919bc315bfd4156238d[flogtanh_SEL-1:0]),
.flogtanh( Ic8f858d7f7a16b771933741d31679dc1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9937af6fcf9d834f308bc3683d524981 = (I1802d759f26dd919bc315bfd4156238d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic8f858d7f7a16b771933741d31679dc1;


Ic3da32f100a43f826b89a492544e7812 I54d7cab766278c006349b1c7c0589cca (
.flogtanh_sel( I2148493e253783fad70f4f2807b83008[flogtanh_SEL-1:0]),
.flogtanh( I9dcf19da38f352fe7fa27c22bff08c19),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I463f4f370e1ecad71de44780eff10df4 = (I2148493e253783fad70f4f2807b83008[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9dcf19da38f352fe7fa27c22bff08c19;


Ic3da32f100a43f826b89a492544e7812 Ic43b6c3cfe97e2292dcbbae85ead8d36 (
.flogtanh_sel( I39e7f78d33aa7f50264908d2efe23634[flogtanh_SEL-1:0]),
.flogtanh( I2bc787aa749db4a5f48bd917715a11d5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I53309409a6059c3bd39f037c23ec3458 = (I39e7f78d33aa7f50264908d2efe23634[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2bc787aa749db4a5f48bd917715a11d5;


Ic3da32f100a43f826b89a492544e7812 I3412014bad8f40f5c8596a53ce51203f (
.flogtanh_sel( I844be5874def16af98de935019f35fe8[flogtanh_SEL-1:0]),
.flogtanh( I3d072e173fd12ac9d802a29a0ff4378c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2603e0b8b93f6680e44c9c8883f6512c = (I844be5874def16af98de935019f35fe8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3d072e173fd12ac9d802a29a0ff4378c;


Ic3da32f100a43f826b89a492544e7812 I660129cd827148d7960a4cb2a6ca39b6 (
.flogtanh_sel( Iee5172ba70a6e368b4903f9ff1d93471[flogtanh_SEL-1:0]),
.flogtanh( I2115d62275a57ec7273e3631c0a32872),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iab354cc9ac1173335c0efeef694f3567 = (Iee5172ba70a6e368b4903f9ff1d93471[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2115d62275a57ec7273e3631c0a32872;


Ic3da32f100a43f826b89a492544e7812 Ib27702f34d6d9a9064cf8edb1ea72f39 (
.flogtanh_sel( I1f34b473283291e0970879465c005e2f[flogtanh_SEL-1:0]),
.flogtanh( I91bc663fcd7f86a066b8b3f93b1dcfc2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6c19936ca2edeb0e261e880a1055e964 = (I1f34b473283291e0970879465c005e2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I91bc663fcd7f86a066b8b3f93b1dcfc2;


Ic3da32f100a43f826b89a492544e7812 Ib7f3c5f1b3d627e0ab306fff3d461ba9 (
.flogtanh_sel( Ie1e0b5120737a7f4bf845618ccd22239[flogtanh_SEL-1:0]),
.flogtanh( I988c0d94f97329dd1cff7d913cb449e7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifebfa58419ecd22a334ed4b67f5c3581 = (Ie1e0b5120737a7f4bf845618ccd22239[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I988c0d94f97329dd1cff7d913cb449e7;


Ic3da32f100a43f826b89a492544e7812 Ie12f94674838a51e9139f0387d7159fa (
.flogtanh_sel( I8abec3020ee5358f8768e5595e9992b4[flogtanh_SEL-1:0]),
.flogtanh( If444a37a85774dcc2769ffd74b785e46),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I71a28e8525f07dabeabe4b4f45f353d0 = (I8abec3020ee5358f8768e5595e9992b4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If444a37a85774dcc2769ffd74b785e46;


Ic3da32f100a43f826b89a492544e7812 I84061f1530957bc7a3926a63a68fa11d (
.flogtanh_sel( I6fe683073211a484cb6e3c416b365d9f[flogtanh_SEL-1:0]),
.flogtanh( Idbb89639b8399b57b190efd898643328),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I514830acdad20c4ff3d078477e939b4b = (I6fe683073211a484cb6e3c416b365d9f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idbb89639b8399b57b190efd898643328;


Ic3da32f100a43f826b89a492544e7812 Ic57710877cacb8a03c27a9068b6e8443 (
.flogtanh_sel( Id7d764da58ade36853e8a45b5ee19dc3[flogtanh_SEL-1:0]),
.flogtanh( Ib1d70f302858eb7c78fb834071616a9b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I036342f6be0f2e2f1f4927099a5c4a78 = (Id7d764da58ade36853e8a45b5ee19dc3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib1d70f302858eb7c78fb834071616a9b;


Ic3da32f100a43f826b89a492544e7812 I514442e48b89cb349a8b86f680826b34 (
.flogtanh_sel( I3cee2fdf353643deac7d6bca20c8fb52[flogtanh_SEL-1:0]),
.flogtanh( I82bd4ea32da7ae3a0d5938fc8a1424c5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iedb655aa25e5f0e35137ec6c3acdc527 = (I3cee2fdf353643deac7d6bca20c8fb52[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I82bd4ea32da7ae3a0d5938fc8a1424c5;


Ic3da32f100a43f826b89a492544e7812 Ib0c7895cbf1ae166ff4e477c025602de (
.flogtanh_sel( Ie9b8f8f0434fe3783c3d8f68fef30e50[flogtanh_SEL-1:0]),
.flogtanh( I6964f2e681e9cdf63fbc0358cb6edcca),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0c59e8c82a31aacbf5977ff778a7ff49 = (Ie9b8f8f0434fe3783c3d8f68fef30e50[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6964f2e681e9cdf63fbc0358cb6edcca;


Ic3da32f100a43f826b89a492544e7812 Ib4909091697a330fd2b3003ef429399a (
.flogtanh_sel( I68cba8ad7742cbb34d0b1fb16be4a58a[flogtanh_SEL-1:0]),
.flogtanh( I41aeb75239ce0d636288e8ceb0665b34),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1b6d20c64b9f23fb6c30f723546aa285 = (I68cba8ad7742cbb34d0b1fb16be4a58a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I41aeb75239ce0d636288e8ceb0665b34;


Ic3da32f100a43f826b89a492544e7812 I5a29ed353f3c5dc5fb2bebd1dfca9933 (
.flogtanh_sel( Idcea56657d40e0fdf9a1c2d920938fd6[flogtanh_SEL-1:0]),
.flogtanh( Ie0d3fd5e7c38c10fdcae3f1b217c28f4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0d66aa55747362354aa81d96057bc4c2 = (Idcea56657d40e0fdf9a1c2d920938fd6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie0d3fd5e7c38c10fdcae3f1b217c28f4;


Ic3da32f100a43f826b89a492544e7812 Ifc92d1d97bc372be37f4b240b5605245 (
.flogtanh_sel( Ic549ffab8f0ce161a177faa2ffd1326d[flogtanh_SEL-1:0]),
.flogtanh( Ia8b7d74eaf227e697c3eb58b31eb355f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1ea33707e40a2e41513fdb3118371437 = (Ic549ffab8f0ce161a177faa2ffd1326d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia8b7d74eaf227e697c3eb58b31eb355f;


Ic3da32f100a43f826b89a492544e7812 I12e444dc3a5a422f1c9ec6fbf2705734 (
.flogtanh_sel( I4d463d500f93f74b2724972ec1d62439[flogtanh_SEL-1:0]),
.flogtanh( I79034cd4180d03348de2c101927048a7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I68c85727adecde0aa8aa66ed08c4b502 = (I4d463d500f93f74b2724972ec1d62439[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I79034cd4180d03348de2c101927048a7;


Ic3da32f100a43f826b89a492544e7812 I6186334ae58166879980196a4192c684 (
.flogtanh_sel( Iba2f362e263953331649c726afa9c481[flogtanh_SEL-1:0]),
.flogtanh( Id23895e0696cdd27e3087294fb52a65b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iebd050e29044153d5881ef80b2db8c28 = (Iba2f362e263953331649c726afa9c481[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id23895e0696cdd27e3087294fb52a65b;


Ic3da32f100a43f826b89a492544e7812 I47687e56550b7c072b3b8a8f65242b40 (
.flogtanh_sel( I6a053d931fb030e03d4882856d3bda75[flogtanh_SEL-1:0]),
.flogtanh( I43939a168f9f5e476262ace39c6ae483),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3c057d64cf4fca0238a874f0ced99c76 = (I6a053d931fb030e03d4882856d3bda75[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I43939a168f9f5e476262ace39c6ae483;


Ic3da32f100a43f826b89a492544e7812 I8c88f2622f0bf7ad4ae5a77a84ba153a (
.flogtanh_sel( I27ede93004e0c240efaa56cc8c570910[flogtanh_SEL-1:0]),
.flogtanh( Ie5167faac3e6510d4b208a1bdc0cd44c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I066cd52173ec5dbce9a3f470d73325af = (I27ede93004e0c240efaa56cc8c570910[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie5167faac3e6510d4b208a1bdc0cd44c;


Ic3da32f100a43f826b89a492544e7812 I0c76ad072804d93cdba16c88d72a5196 (
.flogtanh_sel( I61a11c1711ca10eefea3438722b40bff[flogtanh_SEL-1:0]),
.flogtanh( I1cad8b885a541dd049093ce60c3f8a06),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic7ad59f6a232a997706d17b4098e0324 = (I61a11c1711ca10eefea3438722b40bff[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1cad8b885a541dd049093ce60c3f8a06;


Ic3da32f100a43f826b89a492544e7812 I4e4b3d72471351d05bd62699a33b479e (
.flogtanh_sel( Ia7924c88692cfddf24fb1eff66eacb7e[flogtanh_SEL-1:0]),
.flogtanh( Icd2d69f12d4744ce7b09fce7f27ab830),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icf8cfc800f0a2aa5140a7f83f035b0cc = (Ia7924c88692cfddf24fb1eff66eacb7e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icd2d69f12d4744ce7b09fce7f27ab830;


Ic3da32f100a43f826b89a492544e7812 I7ba543d3d81e23b35b1850246b68e03e (
.flogtanh_sel( Ibcfd01e622f7f5a5156dd9b335b4e5e0[flogtanh_SEL-1:0]),
.flogtanh( Ic9ee0243e36f66f462eb3d4ce93fdde9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6bfbf7ff79ff0a6facc9ba5031239644 = (Ibcfd01e622f7f5a5156dd9b335b4e5e0[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic9ee0243e36f66f462eb3d4ce93fdde9;


Ic3da32f100a43f826b89a492544e7812 I2f486d368f2270674b8782d9d23e4e1a (
.flogtanh_sel( I7f6f418ea51b4298da8758bda3f6a21b[flogtanh_SEL-1:0]),
.flogtanh( I5353c3239ddb4d7fa7094e413b5303b1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I78ade92efd265027807c861be44a10af = (I7f6f418ea51b4298da8758bda3f6a21b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5353c3239ddb4d7fa7094e413b5303b1;


Ic3da32f100a43f826b89a492544e7812 I03616136956550eed69c0d53c917f9de (
.flogtanh_sel( I7185da8937449e23abdd0f39a4b3ed7d[flogtanh_SEL-1:0]),
.flogtanh( Idfca1b1d8041e5808799499e8c8dcf5e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2bc5a10c587d89d10021aa5eaafb490a = (I7185da8937449e23abdd0f39a4b3ed7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idfca1b1d8041e5808799499e8c8dcf5e;


Ic3da32f100a43f826b89a492544e7812 Iebf1eceacf4cb012fda57927c36af5d8 (
.flogtanh_sel( Idc3e3ffa31d9b76c7cf9358a5b2e65d7[flogtanh_SEL-1:0]),
.flogtanh( I4710d61c763098027934286c6a9f3714),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I30080cc6c03bbe933165d266558a822c = (Idc3e3ffa31d9b76c7cf9358a5b2e65d7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4710d61c763098027934286c6a9f3714;


Ic3da32f100a43f826b89a492544e7812 Iaa16f7af8d66dd832af1d9c4783e0cbd (
.flogtanh_sel( I31fe8c887c4aff7c69336676cd31aaa1[flogtanh_SEL-1:0]),
.flogtanh( If6a04c29b7205c5db5f2ff3cf302c45f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7e28234bdf66ab5489d36d15678db797 = (I31fe8c887c4aff7c69336676cd31aaa1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If6a04c29b7205c5db5f2ff3cf302c45f;


Ic3da32f100a43f826b89a492544e7812 Ia4a8d659699ee0d16dfb16f75dc2e08e (
.flogtanh_sel( I59684d5fe6bbb4b54ac097bd25fceef5[flogtanh_SEL-1:0]),
.flogtanh( Ib5d9348a114627a8b1f56aca968d20b1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I74b3c9dd3a8168aacd4369b9ff68fdfd = (I59684d5fe6bbb4b54ac097bd25fceef5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib5d9348a114627a8b1f56aca968d20b1;


Ic3da32f100a43f826b89a492544e7812 Ie18b13c4d332608ae361b7247d45e0fa (
.flogtanh_sel( I86a7cd69148f9590ce91d0aa270d6c54[flogtanh_SEL-1:0]),
.flogtanh( I4e2b59a03731959106d469ffee7b7d33),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia7046faae1ab05978e4b32bd44049fb9 = (I86a7cd69148f9590ce91d0aa270d6c54[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4e2b59a03731959106d469ffee7b7d33;


Ic3da32f100a43f826b89a492544e7812 I5ea8416b1af042ec2d6c033db039a497 (
.flogtanh_sel( Iabce1ccdd968980f622f0e137b159d11[flogtanh_SEL-1:0]),
.flogtanh( Ic6d519691c7543b1bd0707a8c9899088),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0c5250aaca86185fed5978438c8861b6 = (Iabce1ccdd968980f622f0e137b159d11[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic6d519691c7543b1bd0707a8c9899088;


Ic3da32f100a43f826b89a492544e7812 Ibe9d815daef6b021f6cf82c79b07d5ce (
.flogtanh_sel( Iff02977d7b4c733cca1794246f630931[flogtanh_SEL-1:0]),
.flogtanh( Icc6bde490bd8df2ce5efe8cfb24cf5f5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic78949e07e643f571f23df7e8f15d9fb = (Iff02977d7b4c733cca1794246f630931[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icc6bde490bd8df2ce5efe8cfb24cf5f5;


Ic3da32f100a43f826b89a492544e7812 I6099baa4a0bdbae94ecdd8560211e3b8 (
.flogtanh_sel( I9026c904e5ead7ff2994c4f781d61466[flogtanh_SEL-1:0]),
.flogtanh( I861bd8df5caf968dc6edd7a05d690033),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ifb8b3586a5b69b20cf03eabf51344ab6 = (I9026c904e5ead7ff2994c4f781d61466[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I861bd8df5caf968dc6edd7a05d690033;


Ic3da32f100a43f826b89a492544e7812 I13417159878003c4357c5e5bf3a76af3 (
.flogtanh_sel( I99d7489ba87c629c6dd9702a9bbfd3c8[flogtanh_SEL-1:0]),
.flogtanh( I6f44882493f9eadbdbe1ac46a3d2a43b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9ea09f27ce4484f2e7fc3a6b6d6ecb7c = (I99d7489ba87c629c6dd9702a9bbfd3c8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6f44882493f9eadbdbe1ac46a3d2a43b;


Ic3da32f100a43f826b89a492544e7812 I8a045948391b57c3c79d915997bb4705 (
.flogtanh_sel( Ifaf191e0d00ba6da7019c2efcf08e1d9[flogtanh_SEL-1:0]),
.flogtanh( I5a3ec39885fba8d015009d671a1cb544),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If0b9225e759438be175c4128c78605ea = (Ifaf191e0d00ba6da7019c2efcf08e1d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5a3ec39885fba8d015009d671a1cb544;


Ic3da32f100a43f826b89a492544e7812 I0ae1fadba76ede609941439e0988ce47 (
.flogtanh_sel( I4c295991fb08c90862a2f3ba6489000a[flogtanh_SEL-1:0]),
.flogtanh( Ic4e6d76148a8170d1af0c95f370367a5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I33d941ad9d4858fcfb77f0f6cf99d2ec = (I4c295991fb08c90862a2f3ba6489000a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic4e6d76148a8170d1af0c95f370367a5;


Ic3da32f100a43f826b89a492544e7812 I23d8c5e870f2475f3518698121078d1b (
.flogtanh_sel( Iee61d179da125934298400256788cbb8[flogtanh_SEL-1:0]),
.flogtanh( I244bd772f9d750b4e1800e0b0ca67d63),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia0868eee7e7e0640ce1a4d3ca9c001cb = (Iee61d179da125934298400256788cbb8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I244bd772f9d750b4e1800e0b0ca67d63;


Ic3da32f100a43f826b89a492544e7812 Ice9a7abb642f414e712c1b940931cbc8 (
.flogtanh_sel( If87c84440426fb24070372dc1d4bf315[flogtanh_SEL-1:0]),
.flogtanh( I00c203d60e09f1cccdadb8ebff2de650),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icb3ab2c67a87b2ee158e0021b72fc186 = (If87c84440426fb24070372dc1d4bf315[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I00c203d60e09f1cccdadb8ebff2de650;


Ic3da32f100a43f826b89a492544e7812 Ib04bd2633b44e70b4d2d7fca6d9418cd (
.flogtanh_sel( Ib9259a807b31c1b7a528d336bfc403ee[flogtanh_SEL-1:0]),
.flogtanh( I20c7780e77b49d31808e59cae58968a9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5b64997d083769666741c794dd92fb7f = (Ib9259a807b31c1b7a528d336bfc403ee[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I20c7780e77b49d31808e59cae58968a9;


Ic3da32f100a43f826b89a492544e7812 I8c4e156747d4539b4a0677dda038fec9 (
.flogtanh_sel( I411c4d909b2a571e685cd703245516d7[flogtanh_SEL-1:0]),
.flogtanh( Ia332fad029505e5975156f8e13910358),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0a3323aac825506435068f6746aee974 = (I411c4d909b2a571e685cd703245516d7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia332fad029505e5975156f8e13910358;


Ic3da32f100a43f826b89a492544e7812 I67c2529ac0f7cba02e73270ba3244711 (
.flogtanh_sel( If8425453cca8fc8623cb85375c4b8a1d[flogtanh_SEL-1:0]),
.flogtanh( I9cc95185621ad5718a905092c03315f8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibec442c099da091afcf75a7c970bf8ea = (If8425453cca8fc8623cb85375c4b8a1d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9cc95185621ad5718a905092c03315f8;


Ic3da32f100a43f826b89a492544e7812 I625cfb70b6fa2987709bea65abbf07cb (
.flogtanh_sel( I654b497f62df75fa283127b5de29b1ad[flogtanh_SEL-1:0]),
.flogtanh( Iba2a341076f0506aeac3769e71b91f43),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If3a79ede332c39a8d2a276de833242f6 = (I654b497f62df75fa283127b5de29b1ad[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iba2a341076f0506aeac3769e71b91f43;


Ic3da32f100a43f826b89a492544e7812 I523ed12282a559d0154ae052f98619ac (
.flogtanh_sel( I2768519342f7b8a1ee40c1d5ac502b66[flogtanh_SEL-1:0]),
.flogtanh( Ic9e82f153d0e690d5ea47ee159523b72),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I49ccb3e14fe61618806e791ecb4f4eae = (I2768519342f7b8a1ee40c1d5ac502b66[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic9e82f153d0e690d5ea47ee159523b72;


Ic3da32f100a43f826b89a492544e7812 Ib54c9e40b094ddcb3a7792461dfe2439 (
.flogtanh_sel( I8e354c1c5ba44fe5430887248ce0c43b[flogtanh_SEL-1:0]),
.flogtanh( Ia265b95249953a7867c611d475d01169),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I461ebbf3a02ae63e2eb27531b1370f24 = (I8e354c1c5ba44fe5430887248ce0c43b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia265b95249953a7867c611d475d01169;


Ic3da32f100a43f826b89a492544e7812 I9c7df7de90e074eb759943cae32b9265 (
.flogtanh_sel( I8970d8a8aea29913e8696c14c153d16e[flogtanh_SEL-1:0]),
.flogtanh( I5ef2899606d7f08aa6d0028f9f113e38),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice66c108aa66981051df71e226cb0e4d = (I8970d8a8aea29913e8696c14c153d16e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5ef2899606d7f08aa6d0028f9f113e38;


Ic3da32f100a43f826b89a492544e7812 Ia75a2cfd79745c670ef9b0b7e65be876 (
.flogtanh_sel( I3555c6e2fd480a6be11549bf95a9b0b1[flogtanh_SEL-1:0]),
.flogtanh( Idf3a6723fec1ef62c1e37a419590122c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I645ff0d8c0a87ba7f792fc83f342b958 = (I3555c6e2fd480a6be11549bf95a9b0b1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idf3a6723fec1ef62c1e37a419590122c;


Ic3da32f100a43f826b89a492544e7812 I16ac4d1f7e879b2d4b65b9d8db0e140c (
.flogtanh_sel( I8d5600a352e8ba4756f917f912fda6dd[flogtanh_SEL-1:0]),
.flogtanh( I0bde2fc197586c74374ffb402956baf5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ica94017f26e96fb22a47add326ee126e = (I8d5600a352e8ba4756f917f912fda6dd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0bde2fc197586c74374ffb402956baf5;


Ic3da32f100a43f826b89a492544e7812 Ie39ff2f40e0c97a452013d08f13112f4 (
.flogtanh_sel( I7e99d73c95e7ae5c3fe07a3c60ef52eb[flogtanh_SEL-1:0]),
.flogtanh( I9182b3349816b6ddaffde1cbec78339e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id32e7ad5b1aa825732d9b26d0fa02ca1 = (I7e99d73c95e7ae5c3fe07a3c60ef52eb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9182b3349816b6ddaffde1cbec78339e;


Ic3da32f100a43f826b89a492544e7812 I6b1712ed71f6796852f4cff92fbf2dc1 (
.flogtanh_sel( I831633aebe5c6a52b98d630205376f3a[flogtanh_SEL-1:0]),
.flogtanh( I5bf9702e2afd6c791b28c76c84aeb886),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I51b5e641856239367cf43f9b5679b268 = (I831633aebe5c6a52b98d630205376f3a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5bf9702e2afd6c791b28c76c84aeb886;


Ic3da32f100a43f826b89a492544e7812 I51c4b24bdcc943dcfb48540619125594 (
.flogtanh_sel( I82e35482de74223be0d2558334ac2dfb[flogtanh_SEL-1:0]),
.flogtanh( Ifbd7b868d9cb7e04bf2189922bcb9c92),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2d1a5645b126761fc7fb70d24e37189a = (I82e35482de74223be0d2558334ac2dfb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifbd7b868d9cb7e04bf2189922bcb9c92;


Ic3da32f100a43f826b89a492544e7812 I6295920fefd94563a91961e7ed5b1221 (
.flogtanh_sel( Iae2a6f9649ef1bb193e4f0ab5ecbc3e3[flogtanh_SEL-1:0]),
.flogtanh( Ib78e7602e521bc064d5cd9efe10ec6b1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I49f5f87662fbb540d72c94bfd1acd060 = (Iae2a6f9649ef1bb193e4f0ab5ecbc3e3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib78e7602e521bc064d5cd9efe10ec6b1;


Ic3da32f100a43f826b89a492544e7812 I13ee33df653e6e8f19278058de5c2836 (
.flogtanh_sel( Ie8eca65d791ad2f6e8f4ed244f22ae3d[flogtanh_SEL-1:0]),
.flogtanh( I0497115b3dd67c6538039969368e03ae),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I30253dc91301ca27b5732312c01145e0 = (Ie8eca65d791ad2f6e8f4ed244f22ae3d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0497115b3dd67c6538039969368e03ae;


Ic3da32f100a43f826b89a492544e7812 Ic444b4592f1da1512f7c023f26160ea5 (
.flogtanh_sel( Ic24146b01094df9b9ccd455a791f239d[flogtanh_SEL-1:0]),
.flogtanh( Ieba8e28ee660b8e2d78909d61ced3233),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I143f5e324716a94d24ada126886bf895 = (Ic24146b01094df9b9ccd455a791f239d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieba8e28ee660b8e2d78909d61ced3233;


Ic3da32f100a43f826b89a492544e7812 I6f64f03cce94f52d615f8555aa287e78 (
.flogtanh_sel( I1c9031fd54ff9417d44c9fb17dc1fc63[flogtanh_SEL-1:0]),
.flogtanh( I12e6fe32f6159ce6bb8be6411af2b7bb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If64aa8c220b9ab6652e081da7e404e80 = (I1c9031fd54ff9417d44c9fb17dc1fc63[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I12e6fe32f6159ce6bb8be6411af2b7bb;


Ic3da32f100a43f826b89a492544e7812 I26f354f24a092797e87d73bb913d6b51 (
.flogtanh_sel( Idefa20487bc5ba6daff03e6b327d76c6[flogtanh_SEL-1:0]),
.flogtanh( I03392e42f99b06cb65b38122c1e4dc81),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1092325b801600fa7ec85fa640167da9 = (Idefa20487bc5ba6daff03e6b327d76c6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I03392e42f99b06cb65b38122c1e4dc81;


Ic3da32f100a43f826b89a492544e7812 I502b51b80c531fc4ebf2da31063dafb1 (
.flogtanh_sel( I6f984fd9ea27b40ab3afeac8afd29ade[flogtanh_SEL-1:0]),
.flogtanh( I32270eb6cf0594020ee19abb2edfe93d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib028686da9c849e827cf249a744b7db3 = (I6f984fd9ea27b40ab3afeac8afd29ade[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I32270eb6cf0594020ee19abb2edfe93d;


Ic3da32f100a43f826b89a492544e7812 Id528fdf6ce0594d7fcb939bc03e1ef41 (
.flogtanh_sel( I0be92debced4961df5f461fe81e80bf1[flogtanh_SEL-1:0]),
.flogtanh( Ib135d3d7d338f5ff3a1f504aec754bbd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5f3ff7fa8686f7a380302d71b88cfb4b = (I0be92debced4961df5f461fe81e80bf1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib135d3d7d338f5ff3a1f504aec754bbd;


Ic3da32f100a43f826b89a492544e7812 Iacc24303e39b4216b23c2a68d79c3760 (
.flogtanh_sel( Ia7bdaba4c6601b7146498aea6c9a3e07[flogtanh_SEL-1:0]),
.flogtanh( Id9cbc2e4b0f437840f028c7273d49416),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic01904f7c518990eff2dc1de127676c4 = (Ia7bdaba4c6601b7146498aea6c9a3e07[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id9cbc2e4b0f437840f028c7273d49416;


Ic3da32f100a43f826b89a492544e7812 I41193efbb1eef8488f97ddf7a70ab0ab (
.flogtanh_sel( Id450c0a1cabe087be051fbf4158e6016[flogtanh_SEL-1:0]),
.flogtanh( I98b5a84c247422b51abf63a705fbb5f7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I43f2ddd9780f86af489f8deae51168ec = (Id450c0a1cabe087be051fbf4158e6016[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I98b5a84c247422b51abf63a705fbb5f7;


Ic3da32f100a43f826b89a492544e7812 I533d3c82e5232b2ca3ce76b9b3485729 (
.flogtanh_sel( I656d0d69f6e243746b87ad67764dbc3d[flogtanh_SEL-1:0]),
.flogtanh( I0ae39e89061b4f8c5c0e56eba2f48889),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0a013fff6c792363bd7feb03d9691db8 = (I656d0d69f6e243746b87ad67764dbc3d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0ae39e89061b4f8c5c0e56eba2f48889;


Ic3da32f100a43f826b89a492544e7812 I4e2edb90a128904b516b98a1aa48e191 (
.flogtanh_sel( Iab9d870dc1ad159bbaecb20a9b72f005[flogtanh_SEL-1:0]),
.flogtanh( If612cf94a3cefcfb844d6e975ba4aada),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7cf8401bf6893eab0b9f33a0f91ddd05 = (Iab9d870dc1ad159bbaecb20a9b72f005[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If612cf94a3cefcfb844d6e975ba4aada;


Ic3da32f100a43f826b89a492544e7812 I73501caaa0c66c23a09bf28721b9433a (
.flogtanh_sel( Id53b60854f19e095c38f2c255dc57f29[flogtanh_SEL-1:0]),
.flogtanh( I3dab04eb1045e1b3b6bb47e0f4c390ad),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic7ccbeaf4ab94d0660eb7a0533723e24 = (Id53b60854f19e095c38f2c255dc57f29[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3dab04eb1045e1b3b6bb47e0f4c390ad;


Ic3da32f100a43f826b89a492544e7812 I9c98628051943d48097d419973055f06 (
.flogtanh_sel( If9ba44a2e4a8f0b61692fc69ebeb82bd[flogtanh_SEL-1:0]),
.flogtanh( I447db5cb14c9588418037bbb793a6274),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I08043393cb7f2558c145a698ea6652c9 = (If9ba44a2e4a8f0b61692fc69ebeb82bd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I447db5cb14c9588418037bbb793a6274;


Ic3da32f100a43f826b89a492544e7812 I0d62647bebb49e474712d473753800d0 (
.flogtanh_sel( Ief95e8620a1c8ddfd6df673a3a223bd8[flogtanh_SEL-1:0]),
.flogtanh( Ic1227b130f19411495bed64035ea317b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I84865c4f872c0845124b78fabf695c2c = (Ief95e8620a1c8ddfd6df673a3a223bd8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic1227b130f19411495bed64035ea317b;


Ic3da32f100a43f826b89a492544e7812 I450dbbafef894421f919453e0545523c (
.flogtanh_sel( I61519bc0aa02ed461dbb91851d0ae19e[flogtanh_SEL-1:0]),
.flogtanh( I6861b48d33277dd057c6f09ba630d700),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I57b9dd7a7deea6695dcd03439c9723cf = (I61519bc0aa02ed461dbb91851d0ae19e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6861b48d33277dd057c6f09ba630d700;


Ic3da32f100a43f826b89a492544e7812 I174d247b5d5c52b3a5cc288bbcf82245 (
.flogtanh_sel( Ie0c11d584811174a66ca221baf87c36b[flogtanh_SEL-1:0]),
.flogtanh( I022bebca44e2f0b8f9877dd0e709b29f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1cd6b35bcdfd461db69a4c1bdb1d387f = (Ie0c11d584811174a66ca221baf87c36b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I022bebca44e2f0b8f9877dd0e709b29f;


Ic3da32f100a43f826b89a492544e7812 I2989b1a7e719287806cc126c32b445ab (
.flogtanh_sel( If10f4f45ff0fd17541735934ad20f187[flogtanh_SEL-1:0]),
.flogtanh( I8e3d5a48955fe19e24975579d55f4e14),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I40a1ecabded8add5bffe316f2d8beda9 = (If10f4f45ff0fd17541735934ad20f187[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8e3d5a48955fe19e24975579d55f4e14;


Ic3da32f100a43f826b89a492544e7812 I6db3aa1b08b872905f0f90dbea6ebc03 (
.flogtanh_sel( I445919f07a6fa8654211301a9a6126bd[flogtanh_SEL-1:0]),
.flogtanh( I7ee915ffb1c7b8985788c5e6af532ce3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7c52ae4af926267b5e27a530202fcce0 = (I445919f07a6fa8654211301a9a6126bd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7ee915ffb1c7b8985788c5e6af532ce3;


Ic3da32f100a43f826b89a492544e7812 Ic30142e2018ff9879932bdd9f0b212aa (
.flogtanh_sel( I64102b82893352549abd2e2132b19476[flogtanh_SEL-1:0]),
.flogtanh( Ia897087d82c2deac4697755c31766241),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1a5c6c50817db8bde279d5f0b5095d76 = (I64102b82893352549abd2e2132b19476[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia897087d82c2deac4697755c31766241;


Ic3da32f100a43f826b89a492544e7812 Idc80987b1241ef6f1b89c9b27b9aecff (
.flogtanh_sel( I1fc1933fe891ac26f35a42a1b242d919[flogtanh_SEL-1:0]),
.flogtanh( I4c23326dc80b54231289f9f18c4db711),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idf0c1b85712fcbbbcc12915158ebff62 = (I1fc1933fe891ac26f35a42a1b242d919[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4c23326dc80b54231289f9f18c4db711;


Ic3da32f100a43f826b89a492544e7812 I54b19e7dd9da31eea302f3218ad96bd9 (
.flogtanh_sel( I84dfba8bcf8ad3b85f9472fd60d607b5[flogtanh_SEL-1:0]),
.flogtanh( I8326b063a9b9688fb3014667c49ada1b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6b32298e8c61e75d0a38bca3084c0528 = (I84dfba8bcf8ad3b85f9472fd60d607b5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I8326b063a9b9688fb3014667c49ada1b;


Ic3da32f100a43f826b89a492544e7812 I63ce05969f49477fe74e1700d82dd397 (
.flogtanh_sel( I4302fccefe5ee13161f9ad49f9ddf43c[flogtanh_SEL-1:0]),
.flogtanh( Ic41133a438fcea4a1cad9f5e5ee05a03),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5b0d72cedc120406402076148e2d30b0 = (I4302fccefe5ee13161f9ad49f9ddf43c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic41133a438fcea4a1cad9f5e5ee05a03;


Ic3da32f100a43f826b89a492544e7812 Ia48c992069620368c8884a807adc17d5 (
.flogtanh_sel( I59d7153724d3b3805af799692fbe245a[flogtanh_SEL-1:0]),
.flogtanh( I1ac5e426032b874b250cb8adad5b345a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaf624549f73b0d13c1a73c850b99f810 = (I59d7153724d3b3805af799692fbe245a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1ac5e426032b874b250cb8adad5b345a;


Ic3da32f100a43f826b89a492544e7812 I860b806ae381ee99bddb5d9b62140e04 (
.flogtanh_sel( Id1650d0e39be078027493f58e9bbcbdd[flogtanh_SEL-1:0]),
.flogtanh( If9aca7e28f987bf6c7f2fb9b6f11962f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaaf7efeae9f6dc9e8222dc2b10122000 = (Id1650d0e39be078027493f58e9bbcbdd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If9aca7e28f987bf6c7f2fb9b6f11962f;


Ic3da32f100a43f826b89a492544e7812 I278dbdbf1d03d3581a92aeb13ff6ed2e (
.flogtanh_sel( If40ad4aca8dbb3bf7dde8c2ff2e5b8f2[flogtanh_SEL-1:0]),
.flogtanh( Id98a58cd8017fd149ea4f5b295f7ec80),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iea1cd2321d2ac9b891b344e2ba2363d3 = (If40ad4aca8dbb3bf7dde8c2ff2e5b8f2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id98a58cd8017fd149ea4f5b295f7ec80;


Ic3da32f100a43f826b89a492544e7812 If635c8bd23fc7234d8fe2e59d50551e4 (
.flogtanh_sel( Ie49f173549396caeab1d13da36e37c65[flogtanh_SEL-1:0]),
.flogtanh( Ib9e45e75ce8cdd3b548eaf3e41a091ce),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia544fa24b953fe91800978895e3e610e = (Ie49f173549396caeab1d13da36e37c65[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib9e45e75ce8cdd3b548eaf3e41a091ce;


Ic3da32f100a43f826b89a492544e7812 If87a69ebcdba279ba22cd1f970111d0a (
.flogtanh_sel( I3002a0e0cdf8e79bc7186a876410d106[flogtanh_SEL-1:0]),
.flogtanh( I9fcedcbd532cefe1e66ec94b22457cf4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7fa710c37f5f96c3cdc35612a702a71c = (I3002a0e0cdf8e79bc7186a876410d106[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9fcedcbd532cefe1e66ec94b22457cf4;


Ic3da32f100a43f826b89a492544e7812 Ic41ef18644785c9dea69e3d3d76ad18e (
.flogtanh_sel( I2b50fa03f584d10e9af3be085a02a12c[flogtanh_SEL-1:0]),
.flogtanh( Ic627802cf228a709638c14adf83091f8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I98fd105696fca11c1075f9bd30013747 = (I2b50fa03f584d10e9af3be085a02a12c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic627802cf228a709638c14adf83091f8;


Ic3da32f100a43f826b89a492544e7812 I9fb32194e6b2ff18148a61be4e66a9cd (
.flogtanh_sel( If473d172a7bff5aeae99245bbb72978d[flogtanh_SEL-1:0]),
.flogtanh( Ib6bd27a683e11d238fcb775bb44dd913),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I61345963ceabdaa0f25f8a463fc9fe5d = (If473d172a7bff5aeae99245bbb72978d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib6bd27a683e11d238fcb775bb44dd913;


Ic3da32f100a43f826b89a492544e7812 Iac6763d8190a7f31544def1a562589a9 (
.flogtanh_sel( Ib89f7b5625995290a64bcfb143d978ca[flogtanh_SEL-1:0]),
.flogtanh( I3affcbe66b25dc7f11f98b4e444937a2),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9e8375af6af10f4bac3e87e416d430ee = (Ib89f7b5625995290a64bcfb143d978ca[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3affcbe66b25dc7f11f98b4e444937a2;


Ic3da32f100a43f826b89a492544e7812 I25da31087ebccd2bf633db240822dcc5 (
.flogtanh_sel( Iebe0c9b4a87d58a1c55e2ee6b01603c4[flogtanh_SEL-1:0]),
.flogtanh( Ib537657951962c85ad92d43777458588),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ida1cd844022bbf1b8431225e66b2b78f = (Iebe0c9b4a87d58a1c55e2ee6b01603c4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib537657951962c85ad92d43777458588;


Ic3da32f100a43f826b89a492544e7812 Idb8d5cccf82dc4bfa68dae9eee873f88 (
.flogtanh_sel( I104411bb641d2445c7e1385a809bb682[flogtanh_SEL-1:0]),
.flogtanh( Id0af2b1d8b0aa3ba9764ea6a22fafc8c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I30e9ab592e97dbc5fb6ab58d2ffbf8d4 = (I104411bb641d2445c7e1385a809bb682[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id0af2b1d8b0aa3ba9764ea6a22fafc8c;


Ic3da32f100a43f826b89a492544e7812 I4201c4d0b1e09078d310e5fcb2980406 (
.flogtanh_sel( I47dd28b4ae4f7151aff5bb271e35b716[flogtanh_SEL-1:0]),
.flogtanh( I3f934c17beeba9f2d2ca58b3677fe1f3),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2ec2a6de2be39b1bc259b0be72e35a0f = (I47dd28b4ae4f7151aff5bb271e35b716[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3f934c17beeba9f2d2ca58b3677fe1f3;


Ic3da32f100a43f826b89a492544e7812 I2576686eadabda47ae0e79d911ae4e0c (
.flogtanh_sel( I3a27d5573b748df459b90a5a347f9d09[flogtanh_SEL-1:0]),
.flogtanh( Ie3e094ae62dc2a694777f4792c78c886),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic32e349efae2ca419e095ee5e15a501d = (I3a27d5573b748df459b90a5a347f9d09[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie3e094ae62dc2a694777f4792c78c886;


Ic3da32f100a43f826b89a492544e7812 Ibd59cafd11b6731c1e6e40e159c5a3ff (
.flogtanh_sel( I2dbef85d2b2b95af39c3a98c4e143253[flogtanh_SEL-1:0]),
.flogtanh( Idea1d2f5e910ebadc99d356dee8646bd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1befb935ee9cb871c9a7476c1fc0da3f = (I2dbef85d2b2b95af39c3a98c4e143253[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idea1d2f5e910ebadc99d356dee8646bd;


Ic3da32f100a43f826b89a492544e7812 I7307d95396f67a5000c4d6dde4b7da2e (
.flogtanh_sel( I510d39830ae7b0a857ac11baa7c144d3[flogtanh_SEL-1:0]),
.flogtanh( I7cf160bea55d67417a4ee9ce9b252871),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I01c57f697f2af7d2c6ae904319f10725 = (I510d39830ae7b0a857ac11baa7c144d3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7cf160bea55d67417a4ee9ce9b252871;


Ic3da32f100a43f826b89a492544e7812 I333ffd8175ff0f92bdde2890dbd231f3 (
.flogtanh_sel( I2751a94a66ea4cb44c512df4c509937f[flogtanh_SEL-1:0]),
.flogtanh( I196915263bfb62cc21659f81572438b4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id580f8a2748efff9b6b747c497c16e9c = (I2751a94a66ea4cb44c512df4c509937f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I196915263bfb62cc21659f81572438b4;


Ic3da32f100a43f826b89a492544e7812 Ia0b93a9927b1e11ac38ac1270046eeef (
.flogtanh_sel( Ic9a003bfb70ac2da6c229fcad09246d4[flogtanh_SEL-1:0]),
.flogtanh( I548af5c4ccd2816978de565c0c02f176),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I77b54488bd26318f14b4364035cd1836 = (Ic9a003bfb70ac2da6c229fcad09246d4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I548af5c4ccd2816978de565c0c02f176;


Ic3da32f100a43f826b89a492544e7812 I3db014e8dc73657b5011e941c43ac7f3 (
.flogtanh_sel( I34ed986182a3311a8cb005b3dccc224b[flogtanh_SEL-1:0]),
.flogtanh( Ifb7004286169cd9b229b083aea58a408),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I786338397f55073dce91e1c8c5f8e298 = (I34ed986182a3311a8cb005b3dccc224b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifb7004286169cd9b229b083aea58a408;


Ic3da32f100a43f826b89a492544e7812 I7dc26b94819bbe821ea8e0764f9aa819 (
.flogtanh_sel( Ic79281755397f6099ff30c5d07d7e6de[flogtanh_SEL-1:0]),
.flogtanh( Ib04408fcc6f4d26fcdb5599b03b1b534),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0e5931219d94c8e8e1f4af081404dcab = (Ic79281755397f6099ff30c5d07d7e6de[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib04408fcc6f4d26fcdb5599b03b1b534;


Ic3da32f100a43f826b89a492544e7812 If3103d9724829b00ec29c261c1a8907c (
.flogtanh_sel( I8d6559ccc33cbc663584923a55b928b5[flogtanh_SEL-1:0]),
.flogtanh( Ifda1a58a6f54318a30faa98dc1982e8e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8d96b419b010f8076311420d7b9c8a18 = (I8d6559ccc33cbc663584923a55b928b5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifda1a58a6f54318a30faa98dc1982e8e;


Ic3da32f100a43f826b89a492544e7812 If4cf503e643c409e3dc4ec28cea73d5e (
.flogtanh_sel( I4f0a4c241844e390318f11899a0f2c5a[flogtanh_SEL-1:0]),
.flogtanh( I799ce64e6df49e2b62dc6beda4500146),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ife13f962c7a8df3845cde104a959f678 = (I4f0a4c241844e390318f11899a0f2c5a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I799ce64e6df49e2b62dc6beda4500146;


Ic3da32f100a43f826b89a492544e7812 I24dd2cdeba135350b76fae4278c21711 (
.flogtanh_sel( I45fffa266ce3838f82d755b59216a4d6[flogtanh_SEL-1:0]),
.flogtanh( Ia592b65aa89be2fcd981cf144683a298),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7f701ff37ad3fc34d2f4efafe5ff5351 = (I45fffa266ce3838f82d755b59216a4d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia592b65aa89be2fcd981cf144683a298;


Ic3da32f100a43f826b89a492544e7812 I845de6351f6beca36d80512dc360bb00 (
.flogtanh_sel( I8f0e65f5db47d5460d4ec2172807a3e1[flogtanh_SEL-1:0]),
.flogtanh( Ib52365bf14aedf524bb23a4a6fe10551),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I43c815a8ce0b2df9744a525328969691 = (I8f0e65f5db47d5460d4ec2172807a3e1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib52365bf14aedf524bb23a4a6fe10551;


Ic3da32f100a43f826b89a492544e7812 I9a5b2dec4e4606e1f1558dfb14502b22 (
.flogtanh_sel( I34127c0d1af2438e13b6f4709ece80ba[flogtanh_SEL-1:0]),
.flogtanh( Ieba74e8bf3d692612c544af3ce6046fd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6c4a1ded9bf39091cf302ebe0103e2f0 = (I34127c0d1af2438e13b6f4709ece80ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieba74e8bf3d692612c544af3ce6046fd;


Ic3da32f100a43f826b89a492544e7812 I78103c1f21068a9c0bba813ff6893733 (
.flogtanh_sel( I3a67de0e76bbf29d8c77c21865abda2f[flogtanh_SEL-1:0]),
.flogtanh( I6cc1587e659f3f97d636485b708b1eeb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icd4ff8d14af2699db2b5168027894ebb = (I3a67de0e76bbf29d8c77c21865abda2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6cc1587e659f3f97d636485b708b1eeb;


Ic3da32f100a43f826b89a492544e7812 Ib5064cb3cf001b8a99212aaadee06b9d (
.flogtanh_sel( Ic64e64aeb754249b868e14311ea19759[flogtanh_SEL-1:0]),
.flogtanh( I84b09aba55d2335f19faa5762aeedb89),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia79d52fe2130426c07890fcaa50137db = (Ic64e64aeb754249b868e14311ea19759[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I84b09aba55d2335f19faa5762aeedb89;


Ic3da32f100a43f826b89a492544e7812 I07987b16b313b685813c635fdc7adea7 (
.flogtanh_sel( Ic4aa0dc9014c8445f8d9a7723d7263f5[flogtanh_SEL-1:0]),
.flogtanh( I3c4b9082ba72cade4d52924eff135135),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I308aaa8ac500b5589aa4af533a9062bf = (Ic4aa0dc9014c8445f8d9a7723d7263f5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3c4b9082ba72cade4d52924eff135135;


Ic3da32f100a43f826b89a492544e7812 I31ac6d0c4276c60aabee4e0551dded9a (
.flogtanh_sel( I47b988d017580bdfe8f443904b1f3aac[flogtanh_SEL-1:0]),
.flogtanh( I65f6c14ae4e7139fd858d7637ec3fd46),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iac91f4037e542d9fda30fadafe7e79ac = (I47b988d017580bdfe8f443904b1f3aac[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I65f6c14ae4e7139fd858d7637ec3fd46;


Ic3da32f100a43f826b89a492544e7812 I49a309080c74c55e248856f2d1bfb69c (
.flogtanh_sel( Ica9ff13e8c3850be6c70b0b06c1d9fbf[flogtanh_SEL-1:0]),
.flogtanh( I02425810db970e5ef0b791dc4be103a9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8cd5970682bc84881489c12ff073212c = (Ica9ff13e8c3850be6c70b0b06c1d9fbf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I02425810db970e5ef0b791dc4be103a9;


Ic3da32f100a43f826b89a492544e7812 I122cf9e037c0943593493c409ca7db6b (
.flogtanh_sel( If2efeb489911f295dd7722cb22ea521d[flogtanh_SEL-1:0]),
.flogtanh( Id0bc7b00dec58136a8016979d8a9faad),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1ee27be7e1a38aff0039b21c45f406d1 = (If2efeb489911f295dd7722cb22ea521d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id0bc7b00dec58136a8016979d8a9faad;


Ic3da32f100a43f826b89a492544e7812 I55c0e94fb8f677783b44556b31566df0 (
.flogtanh_sel( Iaa16dffcc01e41e6ff17e92bdefe3df5[flogtanh_SEL-1:0]),
.flogtanh( I7c61892052c3c32343ed172d4ae354cc),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idf90f01353ad1057e11fd060442f4e53 = (Iaa16dffcc01e41e6ff17e92bdefe3df5[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7c61892052c3c32343ed172d4ae354cc;


Ic3da32f100a43f826b89a492544e7812 I7e367ba994f0ce92f0fcdc2efa3e7c02 (
.flogtanh_sel( Ie8857b9841fbd795a4192976ef7ecc25[flogtanh_SEL-1:0]),
.flogtanh( I7cd312338aa5a86e1b05cc28ab7a2b23),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id45f4e0f142b6c3925f24a37dcf7c0ae = (Ie8857b9841fbd795a4192976ef7ecc25[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7cd312338aa5a86e1b05cc28ab7a2b23;


Ic3da32f100a43f826b89a492544e7812 I41547a01e1721217848fefc522f14954 (
.flogtanh_sel( If12aef69eea28052aa3bdb6ac31af205[flogtanh_SEL-1:0]),
.flogtanh( I88d4372b4f7bfddd2af726c2df391287),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I52a9bcfbd2d3a763671f19cfeaf7bb8b = (If12aef69eea28052aa3bdb6ac31af205[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I88d4372b4f7bfddd2af726c2df391287;


Ic3da32f100a43f826b89a492544e7812 I29b72fef263a81166d14a1138932d9c6 (
.flogtanh_sel( I0b3c6162ae2b9221738a18a29489887f[flogtanh_SEL-1:0]),
.flogtanh( Ic8978ad86275ac6f4a0cf80ebefc5b27),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia3cc6acf2cae41e560e09993007ffd2b = (I0b3c6162ae2b9221738a18a29489887f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic8978ad86275ac6f4a0cf80ebefc5b27;


Ic3da32f100a43f826b89a492544e7812 I453a66ca7a6ddf07f50693094e15bdfd (
.flogtanh_sel( I08211bba29e87faf4079152bcc973e7d[flogtanh_SEL-1:0]),
.flogtanh( I99745124c45f37d3882064590394a0aa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iba0d2f08788f2208a648ae7b5414195d = (I08211bba29e87faf4079152bcc973e7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I99745124c45f37d3882064590394a0aa;


Ic3da32f100a43f826b89a492544e7812 Ia4195932342cae834eeb7578df124b7d (
.flogtanh_sel( Ibff3da265f1c3f21548f5b019e1a9dc1[flogtanh_SEL-1:0]),
.flogtanh( I33fe34f9be3c51b4b93f89c3f862e332),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9f7df6ad60284c812aeb522974578e0b = (Ibff3da265f1c3f21548f5b019e1a9dc1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I33fe34f9be3c51b4b93f89c3f862e332;


Ic3da32f100a43f826b89a492544e7812 I0459a8ee45e2acfc69c15ffa657a96d2 (
.flogtanh_sel( Ie9fa1762d7844b0d781afdfb0771cea9[flogtanh_SEL-1:0]),
.flogtanh( Iecda9a183e74f78b9fd5ce34e80d712e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iab1fb7006598181bd8749ed90c519b13 = (Ie9fa1762d7844b0d781afdfb0771cea9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iecda9a183e74f78b9fd5ce34e80d712e;


Ic3da32f100a43f826b89a492544e7812 I41a6c7b1fd7f1cd6bee3d02e9337c147 (
.flogtanh_sel( Ia677d504b9f7fc2698c0345f236428ba[flogtanh_SEL-1:0]),
.flogtanh( I5293b996bbf152abf110df1205ad4856),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieef3b299ec35075c71ef9fb10525bfc4 = (Ia677d504b9f7fc2698c0345f236428ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5293b996bbf152abf110df1205ad4856;


Ic3da32f100a43f826b89a492544e7812 I9a3861c2b2068be74e2b5da53789c4b4 (
.flogtanh_sel( Idebce29121c0481df83d755b60ff632c[flogtanh_SEL-1:0]),
.flogtanh( Ia99c08ee345bdc1489ce82a62481ef3b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I58a7c08adf48d0737c5803e2a818c045 = (Idebce29121c0481df83d755b60ff632c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia99c08ee345bdc1489ce82a62481ef3b;


Ic3da32f100a43f826b89a492544e7812 I507b2febb42b9c336c4ca442801d15ef (
.flogtanh_sel( Iad2c780a6386674d50cca54d8c4ebd86[flogtanh_SEL-1:0]),
.flogtanh( Iaa314530e04145eb73672ebb150858af),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I30a1c8fcd9a510a6ed559f07dd809b90 = (Iad2c780a6386674d50cca54d8c4ebd86[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iaa314530e04145eb73672ebb150858af;


Ic3da32f100a43f826b89a492544e7812 Iee55e7f1b448c7684b887f970ea182d6 (
.flogtanh_sel( If1d7944e7c4828ddb91ffea28609cbc7[flogtanh_SEL-1:0]),
.flogtanh( I05f7363bfcc34691280079e82f6f5449),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic4f5e9d49419e1c57cfa387761ab643d = (If1d7944e7c4828ddb91ffea28609cbc7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I05f7363bfcc34691280079e82f6f5449;


Ic3da32f100a43f826b89a492544e7812 I47c162f63f223552f690bb29493b8be6 (
.flogtanh_sel( I843a68ceb0adab829091f31d0de56eb6[flogtanh_SEL-1:0]),
.flogtanh( Ica5ce135e77ed1d7cbc8277344ffeaeb),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id3dd71ea0bf0f2996fbe42b8c3318762 = (I843a68ceb0adab829091f31d0de56eb6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ica5ce135e77ed1d7cbc8277344ffeaeb;


Ic3da32f100a43f826b89a492544e7812 I46ef8dd6d06dc52635d66f393a3f0bac (
.flogtanh_sel( I59701b9eb54dda2744a79cebe7d73f3b[flogtanh_SEL-1:0]),
.flogtanh( Iac98c702c4d9d78460fc7c212bce7841),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib834b91bf81067e8efa9d470023e8b9d = (I59701b9eb54dda2744a79cebe7d73f3b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iac98c702c4d9d78460fc7c212bce7841;


Ic3da32f100a43f826b89a492544e7812 I1705314f8e142466610b5adb5af0d5a0 (
.flogtanh_sel( If63cf5e8f47e4e51176401f0d954ea23[flogtanh_SEL-1:0]),
.flogtanh( I1fe269380ba03e78a8e41c17aa4bd757),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic6ead78ed741442f17a15a157cd6ef9c = (If63cf5e8f47e4e51176401f0d954ea23[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1fe269380ba03e78a8e41c17aa4bd757;


Ic3da32f100a43f826b89a492544e7812 I8e55722b79fe2ea3d9afc8c546629738 (
.flogtanh_sel( Id09454844b525697de3e3727d89551e4[flogtanh_SEL-1:0]),
.flogtanh( Ib19549130ee3307413b69c50042f7302),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4e257dbd6f196a02dc0f5a2e5f6047d7 = (Id09454844b525697de3e3727d89551e4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib19549130ee3307413b69c50042f7302;


Ic3da32f100a43f826b89a492544e7812 I12dbfce9f98fb8ef277b4408a4c06bf4 (
.flogtanh_sel( I6d1b2ce4368945b56eee7814638471cc[flogtanh_SEL-1:0]),
.flogtanh( Iad6acaf97d307fdbe0f20bf010acb468),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3dbfbd34d1fdfd4f422d900154123b6b = (I6d1b2ce4368945b56eee7814638471cc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iad6acaf97d307fdbe0f20bf010acb468;


Ic3da32f100a43f826b89a492544e7812 Ibab8cb9bc13be76eaeb076f79edc4283 (
.flogtanh_sel( I6079945faa57335b1c902ccf7f960a70[flogtanh_SEL-1:0]),
.flogtanh( I67c9882f9e19df5a7b9bd0d900bb2f75),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I529b763dace1924613d184c6c70c2708 = (I6079945faa57335b1c902ccf7f960a70[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I67c9882f9e19df5a7b9bd0d900bb2f75;


Ic3da32f100a43f826b89a492544e7812 I94ab36ac1f8f613ae3c0dd3c539454dc (
.flogtanh_sel( Ie7752906ac55cf51f3e96e8c0046f1aa[flogtanh_SEL-1:0]),
.flogtanh( I3099768bc986a11350656e472fc21ac1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7a600aeb6cf8c3311c10afa4d82767a1 = (Ie7752906ac55cf51f3e96e8c0046f1aa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3099768bc986a11350656e472fc21ac1;


Ic3da32f100a43f826b89a492544e7812 I5137c20d83b2058d562a4bcbb47f3bb0 (
.flogtanh_sel( I2d7d4135a94f5df949283c043228791f[flogtanh_SEL-1:0]),
.flogtanh( Ifba5972f9d38199dbc675432a29934e4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8c7aab31f8cb705ea13a41a5bd349303 = (I2d7d4135a94f5df949283c043228791f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifba5972f9d38199dbc675432a29934e4;


Ic3da32f100a43f826b89a492544e7812 I7e377ea010a57e6d6b2af33313847851 (
.flogtanh_sel( I99c75e3d26c5d01f6ae9abcd05407d8c[flogtanh_SEL-1:0]),
.flogtanh( I0934fb292b19451a050fb3374a7bd1a7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I171149dcaab2c0f0e2a10547ad95084d = (I99c75e3d26c5d01f6ae9abcd05407d8c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0934fb292b19451a050fb3374a7bd1a7;


Ic3da32f100a43f826b89a492544e7812 Ib5536c4d92da5817957f8fa20780019e (
.flogtanh_sel( I81e6f97621dbfb2fed6fc236005a2b19[flogtanh_SEL-1:0]),
.flogtanh( I9a3d1741c77fb1bbc1a54383874de82a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I23b60ca4da2df0ec40c1df62d058deef = (I81e6f97621dbfb2fed6fc236005a2b19[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9a3d1741c77fb1bbc1a54383874de82a;


Ic3da32f100a43f826b89a492544e7812 I3c3ff8b5625fc01b6fe4c10ed3851b44 (
.flogtanh_sel( Ieac60532dcfc916a65054e35cf31d6d2[flogtanh_SEL-1:0]),
.flogtanh( If89f2ce813bab91af88f73ddc570d5a1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7978d2d800b4438d0644ae3df6bcac9c = (Ieac60532dcfc916a65054e35cf31d6d2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If89f2ce813bab91af88f73ddc570d5a1;


Ic3da32f100a43f826b89a492544e7812 I0d138477b99cb1a594f9e019da8fb474 (
.flogtanh_sel( Ib7eb83ba73e0dc17f69c357b6ca555bf[flogtanh_SEL-1:0]),
.flogtanh( Ibc0dfcffac26f4898d42808534f6588f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibc4eddc0f1768e9ec7e38e951a28ec42 = (Ib7eb83ba73e0dc17f69c357b6ca555bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibc0dfcffac26f4898d42808534f6588f;


Ic3da32f100a43f826b89a492544e7812 I2a52739a417d5f48d370614b3ce6e4e7 (
.flogtanh_sel( I5139d8a7a099e3c619c60647c15b7420[flogtanh_SEL-1:0]),
.flogtanh( I3a0a6f3d0141e8ad04d89c4bf306a96f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1c97fd1d21a31af8b5498a79b1a3e7b6 = (I5139d8a7a099e3c619c60647c15b7420[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3a0a6f3d0141e8ad04d89c4bf306a96f;


Ic3da32f100a43f826b89a492544e7812 I4a725d3a4c90b94978ab59ce3cbf52db (
.flogtanh_sel( I6ccd2e11ebd5b2de80b120e20650a602[flogtanh_SEL-1:0]),
.flogtanh( I1c875571dd1be1bb28aa15554964b485),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie4f063eeaf7ee3f033e2a01ffaca623e = (I6ccd2e11ebd5b2de80b120e20650a602[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1c875571dd1be1bb28aa15554964b485;


Ic3da32f100a43f826b89a492544e7812 I3cdec5a824d31049ee8bfc11a6d0fecc (
.flogtanh_sel( Ie669cebe5fe39e1a841f8dd3c1f6bc57[flogtanh_SEL-1:0]),
.flogtanh( Ide5d5fdcf86b369b015890030a222a0a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibb3d57d510cad00064a331f61f6400a2 = (Ie669cebe5fe39e1a841f8dd3c1f6bc57[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ide5d5fdcf86b369b015890030a222a0a;


Ic3da32f100a43f826b89a492544e7812 Iee9c291e2aef4bb16f36cf96a339ece8 (
.flogtanh_sel( If32acb9fc212c4af34099acf6df2bc5a[flogtanh_SEL-1:0]),
.flogtanh( I7cf6e8d40e7bd7685a7260638523690c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I9485ae915474a31562ce358666d66245 = (If32acb9fc212c4af34099acf6df2bc5a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7cf6e8d40e7bd7685a7260638523690c;


Ic3da32f100a43f826b89a492544e7812 Idb21cd21d51ae816f45827dda58c63c7 (
.flogtanh_sel( I075ce236a181bf925c8ccce91d9bc8cd[flogtanh_SEL-1:0]),
.flogtanh( I52ccac771cc9a1c1797862bc781e1f58),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia54b6f7044a831020e49f1bf48bc063a = (I075ce236a181bf925c8ccce91d9bc8cd[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I52ccac771cc9a1c1797862bc781e1f58;


Ic3da32f100a43f826b89a492544e7812 Ie0766d36070d4c063601b1762bd8134f (
.flogtanh_sel( I541d4e422b999a0dfca44d275178e1d9[flogtanh_SEL-1:0]),
.flogtanh( I9db2090916f2535b14ed3292e78baa32),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie71c7babb5d17378d40444b6bbd4e7a6 = (I541d4e422b999a0dfca44d275178e1d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9db2090916f2535b14ed3292e78baa32;


Ic3da32f100a43f826b89a492544e7812 Ice445dd26ded3e46da2725577897197a (
.flogtanh_sel( I3e02657f3d9f79338cd083ed024bf96c[flogtanh_SEL-1:0]),
.flogtanh( I5b77a8ce7f495ae61315d1590bfd71b8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia0977b79857bdbf058535c30e338c38a = (I3e02657f3d9f79338cd083ed024bf96c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5b77a8ce7f495ae61315d1590bfd71b8;


Ic3da32f100a43f826b89a492544e7812 Ibab35e8130d66fd85afac3a72d7effa9 (
.flogtanh_sel( Ia5e5537405ab8edcc7cd43c86837d43d[flogtanh_SEL-1:0]),
.flogtanh( I4e4bb795cf09757c8ad3933c9ce4686f),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I600ea1371a2be66430ac9534583b512b = (Ia5e5537405ab8edcc7cd43c86837d43d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4e4bb795cf09757c8ad3933c9ce4686f;


Ic3da32f100a43f826b89a492544e7812 I80588561b3244853002de1cfe9c1ab55 (
.flogtanh_sel( I07ff388e3b6c7288f0f6c35a345023fe[flogtanh_SEL-1:0]),
.flogtanh( I78c29808e737dab48b5144b232dd02f6),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ife5b9afdbb30c122b84d5378f9cb366d = (I07ff388e3b6c7288f0f6c35a345023fe[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I78c29808e737dab48b5144b232dd02f6;


Ic3da32f100a43f826b89a492544e7812 I75aae9040c2cb58a397872fae81bcae1 (
.flogtanh_sel( I56cb3b3e193ca5068734417fd0ec4e02[flogtanh_SEL-1:0]),
.flogtanh( Ie2ae83a457d79fbddc640d49d626171c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I27556d599dd1a27ee8f49e819ccbf29a = (I56cb3b3e193ca5068734417fd0ec4e02[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie2ae83a457d79fbddc640d49d626171c;


Ic3da32f100a43f826b89a492544e7812 I0b17547d5a1120d61719d5f79881d07d (
.flogtanh_sel( I5bbf1765d8f81581d0cf31c0bc755fb3[flogtanh_SEL-1:0]),
.flogtanh( I3711e49a4eec517e47897fb731d75958),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icce595233ce089eafcca3eae5e71e5f8 = (I5bbf1765d8f81581d0cf31c0bc755fb3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3711e49a4eec517e47897fb731d75958;


Ic3da32f100a43f826b89a492544e7812 Ied9e089fca20b452bc0b69adb33d9722 (
.flogtanh_sel( Iaa1643095e518846cdede4d5a90dff84[flogtanh_SEL-1:0]),
.flogtanh( Ifda4e727eb6275266f583badb6d4a9ed),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icc3cadf40c09be1a8c2847caf0e3e63c = (Iaa1643095e518846cdede4d5a90dff84[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifda4e727eb6275266f583badb6d4a9ed;


Ic3da32f100a43f826b89a492544e7812 Icc5ce12ba2f3023af06d7465a59c65ea (
.flogtanh_sel( Iee6e12f4717a3279dd31b874eabae69e[flogtanh_SEL-1:0]),
.flogtanh( I2be66a82c7b58e3c14b5816522b46969),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib43886d923b8c683004713ff25b2f90d = (Iee6e12f4717a3279dd31b874eabae69e[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2be66a82c7b58e3c14b5816522b46969;


Ic3da32f100a43f826b89a492544e7812 Ib67fec8dc662f360a38b0723887d5484 (
.flogtanh_sel( Ic52a9edbbc5283844d2514ea142ca6e2[flogtanh_SEL-1:0]),
.flogtanh( I826fe7ad9e67061800d5d6543d779864),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I132d9671c582876568c0f7f5335f5227 = (Ic52a9edbbc5283844d2514ea142ca6e2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I826fe7ad9e67061800d5d6543d779864;


Ic3da32f100a43f826b89a492544e7812 I7958a073e758f1677a701f2a1ed5588b (
.flogtanh_sel( Ice3e978c8da2a7de5b28542a5589f0a2[flogtanh_SEL-1:0]),
.flogtanh( Ic0c9069041758b53f56a46da81dd2d60),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I0859c80b42a8c60dade8f05d58ee3701 = (Ice3e978c8da2a7de5b28542a5589f0a2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic0c9069041758b53f56a46da81dd2d60;


Ic3da32f100a43f826b89a492544e7812 I5272726ee65396592886d396d182ce4b (
.flogtanh_sel( I336a425aed221c85ca80b9a97d21d6b1[flogtanh_SEL-1:0]),
.flogtanh( I6f4c5a8de7690fec959861f43c134915),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib3690ec149adde94343d3e617931a287 = (I336a425aed221c85ca80b9a97d21d6b1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6f4c5a8de7690fec959861f43c134915;


Ic3da32f100a43f826b89a492544e7812 Ic6b5092bd1b6fa783bb3f5a6c109b8db (
.flogtanh_sel( Ie477c0f3b77bb299ba8b1a410d211ef7[flogtanh_SEL-1:0]),
.flogtanh( I14f1005a8c0fbdc5ca02c032b8891c2b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I41f2bf9ff00f983ad1298c8c83b041cb = (Ie477c0f3b77bb299ba8b1a410d211ef7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I14f1005a8c0fbdc5ca02c032b8891c2b;


Ic3da32f100a43f826b89a492544e7812 I230468305e3c4b09205ac4d54ca8ce78 (
.flogtanh_sel( Ie62920d089ae762603cd33fbf97d92bb[flogtanh_SEL-1:0]),
.flogtanh( Iacd30dfb96f6572ec56eff0a4094ec04),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib5414585cd6976cfce42e42190cc08d7 = (Ie62920d089ae762603cd33fbf97d92bb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Iacd30dfb96f6572ec56eff0a4094ec04;


Ic3da32f100a43f826b89a492544e7812 I61c630e438e3e38a56dca4be38bc10c8 (
.flogtanh_sel( I2ca952e4e676537fd5a8fc71ecfa10e9[flogtanh_SEL-1:0]),
.flogtanh( I1c748b8fe4979331bc3fe5aff4b6f9f4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1ca59325ff30db83df5bf0a2cd9706b6 = (I2ca952e4e676537fd5a8fc71ecfa10e9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1c748b8fe4979331bc3fe5aff4b6f9f4;


Ic3da32f100a43f826b89a492544e7812 Iea549632a9ba59a19cde8a0c56c23890 (
.flogtanh_sel( Iefd31e7ff3c829c88f60bc89d70afcf7[flogtanh_SEL-1:0]),
.flogtanh( I158c7973974f36c2793127964e50d1bd),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ie2f5b03f3b136e651b8aba92a30d298a = (Iefd31e7ff3c829c88f60bc89d70afcf7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I158c7973974f36c2793127964e50d1bd;


Ic3da32f100a43f826b89a492544e7812 I7f69bbf879c4c1bb0faffbd3ff7a11e7 (
.flogtanh_sel( Iafa987a413fd8fcacfe872bc0f5bc2d6[flogtanh_SEL-1:0]),
.flogtanh( Id5ea6ba2402275cb925a1848b31ec2e1),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I312ce79a8dd2ce3d37c930d42640509b = (Iafa987a413fd8fcacfe872bc0f5bc2d6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id5ea6ba2402275cb925a1848b31ec2e1;


Ic3da32f100a43f826b89a492544e7812 Ied6840820b1ec1047d2f2178bcf08919 (
.flogtanh_sel( I305c1ea420d666f258e38c5a65847367[flogtanh_SEL-1:0]),
.flogtanh( I3862f7017bc2bc69844b73f2a79f47f5),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I467d5e2554ef25873e0b44e947ee0011 = (I305c1ea420d666f258e38c5a65847367[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3862f7017bc2bc69844b73f2a79f47f5;


Ic3da32f100a43f826b89a492544e7812 Ica0b6384a76e23a71c66a9d0da8f1ab1 (
.flogtanh_sel( I9f040c4088bfab72d74e5332e9710d1a[flogtanh_SEL-1:0]),
.flogtanh( I4ed41fde5449b7112baf000a05484ac4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ice73b514709469fd21cd254bf4ceadd9 = (I9f040c4088bfab72d74e5332e9710d1a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4ed41fde5449b7112baf000a05484ac4;


Ic3da32f100a43f826b89a492544e7812 Idd0410d9a0c61943d37acafda9f6f549 (
.flogtanh_sel( Ia2f41f9778324a06daeb185c736516a4[flogtanh_SEL-1:0]),
.flogtanh( I40c4db2872b602bf9d6a4fc4ba5ac34d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I45ba06a6d6f00c174b1439a6f226a085 = (Ia2f41f9778324a06daeb185c736516a4[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I40c4db2872b602bf9d6a4fc4ba5ac34d;


Ic3da32f100a43f826b89a492544e7812 I7f3ee1368f93b7f9fe31333753dc88e4 (
.flogtanh_sel( Id9778ba5fbdbed4d33a092da6b68c414[flogtanh_SEL-1:0]),
.flogtanh( Ibe5ab52bd0f220f7a6aac244c0e3867e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic8a272f82736fd599fb3250e970edf9b = (Id9778ba5fbdbed4d33a092da6b68c414[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibe5ab52bd0f220f7a6aac244c0e3867e;


Ic3da32f100a43f826b89a492544e7812 I542d8156bf34653e118605d86f21a6ea (
.flogtanh_sel( I27c2c79d0d719c71c8e28218d1174a13[flogtanh_SEL-1:0]),
.flogtanh( I36668064f280c70f9143ee9f39973015),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5b9710b16effc8bf0695517c6e651836 = (I27c2c79d0d719c71c8e28218d1174a13[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I36668064f280c70f9143ee9f39973015;


Ic3da32f100a43f826b89a492544e7812 I19a302a8d0994bb4a7d9c1836f8c40d3 (
.flogtanh_sel( I2a9d6a774769b12ae20bc0cee0c36f5c[flogtanh_SEL-1:0]),
.flogtanh( Ief92462253c5a03a42d46ed7087caf9a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I038b42a83025f5eaebf45799d1ebe7b0 = (I2a9d6a774769b12ae20bc0cee0c36f5c[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ief92462253c5a03a42d46ed7087caf9a;


Ic3da32f100a43f826b89a492544e7812 I41aaf5ea46311cd142e89977231cdcb5 (
.flogtanh_sel( I2c567b75f1399c069b95284f4c36b6d1[flogtanh_SEL-1:0]),
.flogtanh( Idf196345491ff3290796ba7827d31c17),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I73ddd7cf9272ceab5a663e2244e72d7e = (I2c567b75f1399c069b95284f4c36b6d1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Idf196345491ff3290796ba7827d31c17;


Ic3da32f100a43f826b89a492544e7812 Iee41216450c0faedbed2ddb257e7328f (
.flogtanh_sel( If3d3eb609abfd6e315eec803d2e94490[flogtanh_SEL-1:0]),
.flogtanh( I2230f0e48899877bc2bcb3538be81bfa),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I16507fab8f9076bfeb419896fa7cdc1d = (If3d3eb609abfd6e315eec803d2e94490[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I2230f0e48899877bc2bcb3538be81bfa;


Ic3da32f100a43f826b89a492544e7812 Ib74a0ac782c0e0851b1503d88be5caa7 (
.flogtanh_sel( I9c58aea7ce986b1d28f5808b347c015d[flogtanh_SEL-1:0]),
.flogtanh( Ibc0ec83d6b8e6be89ddc88ef83f0b03d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3dd1f28cf199299aba54e47a429c9b11 = (I9c58aea7ce986b1d28f5808b347c015d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibc0ec83d6b8e6be89ddc88ef83f0b03d;


Ic3da32f100a43f826b89a492544e7812 I474fee670a1a5ab4fcd7e6f5ed1a711f (
.flogtanh_sel( Id139c7a783196941100003b6cb0cd1e7[flogtanh_SEL-1:0]),
.flogtanh( Ifc59c1b26ec09b3a7fe5a2b90511c93b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I49d9203dc6f8c17f17383e8f7e01f005 = (Id139c7a783196941100003b6cb0cd1e7[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifc59c1b26ec09b3a7fe5a2b90511c93b;


Ic3da32f100a43f826b89a492544e7812 Ibbe99afdefe88211d77485890c5eaba0 (
.flogtanh_sel( I524d7614b01460778da3ce98f6aaa3d9[flogtanh_SEL-1:0]),
.flogtanh( I9c6fc8e09cd63551f40accc98d784a44),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibeec86c75d950ee00dd63a2930f08a24 = (I524d7614b01460778da3ce98f6aaa3d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9c6fc8e09cd63551f40accc98d784a44;


Ic3da32f100a43f826b89a492544e7812 Ib43408e334d2438d3dc596bc50833e4a (
.flogtanh_sel( I8acda65f116d5c91cbe2662ac282aa31[flogtanh_SEL-1:0]),
.flogtanh( I26692a6aab1d81d71219a436bee5e10b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I47b2438c3680b2d816168df37d7c491c = (I8acda65f116d5c91cbe2662ac282aa31[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I26692a6aab1d81d71219a436bee5e10b;


Ic3da32f100a43f826b89a492544e7812 I0885b092568781505f8786acda74cd7c (
.flogtanh_sel( If67dbe22f8d22b3430215fb0deae8204[flogtanh_SEL-1:0]),
.flogtanh( Ieb50592e17305d0f74cbf216be947862),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5983bf2c6c90b872ee6cf58b5e520311 = (If67dbe22f8d22b3430215fb0deae8204[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieb50592e17305d0f74cbf216be947862;


Ic3da32f100a43f826b89a492544e7812 I14af4556909858c19f4582fdb963fc6b (
.flogtanh_sel( I9a35cd7512787263abedd6d9913cf507[flogtanh_SEL-1:0]),
.flogtanh( I0071f023f1be4400541c13bc68278417),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I6745cacecb7ee86cf3c7ad7eeee6048f = (I9a35cd7512787263abedd6d9913cf507[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0071f023f1be4400541c13bc68278417;


Ic3da32f100a43f826b89a492544e7812 Iae53a24e464bf8d721cf387df914eff7 (
.flogtanh_sel( If9cca23469c5e6001650f1f8b1360ae8[flogtanh_SEL-1:0]),
.flogtanh( Ib2f1635b38ca6090e5ff633cbfa13273),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib9672d20643d856ff31905ab14c0ac87 = (If9cca23469c5e6001650f1f8b1360ae8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib2f1635b38ca6090e5ff633cbfa13273;


Ic3da32f100a43f826b89a492544e7812 I34be2423dca79ec822a6b4db71f8a30d (
.flogtanh_sel( Icc2606ae8f9a3b425225ae7339112b9d[flogtanh_SEL-1:0]),
.flogtanh( Id2c0bc90fd26e82fe91b5aef7bdd3a29),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib9dfea1f34a120eda30d5bd919365a6a = (Icc2606ae8f9a3b425225ae7339112b9d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id2c0bc90fd26e82fe91b5aef7bdd3a29;


Ic3da32f100a43f826b89a492544e7812 Ibb723d8d375ff6f531f205a36407845d (
.flogtanh_sel( I34aa1802d24e074ae54563898929abfa[flogtanh_SEL-1:0]),
.flogtanh( If4a723ce836f5327b85e234ebd195bd9),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia7bf82c9e5ca4467b5e50beeaeb975e9 = (I34aa1802d24e074ae54563898929abfa[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If4a723ce836f5327b85e234ebd195bd9;


Ic3da32f100a43f826b89a492544e7812 I29b9b7bd378ed0e4c4bc0dd7818533a9 (
.flogtanh_sel( Icb85b3464dc40e8504c53c377e889c45[flogtanh_SEL-1:0]),
.flogtanh( If63dd5997e033817126a9ebaf38c1955),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I327c9acb8934729b4ea5486787afa2e8 = (Icb85b3464dc40e8504c53c377e889c45[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: If63dd5997e033817126a9ebaf38c1955;


Ic3da32f100a43f826b89a492544e7812 I02408e34541d748c107b16f4c974e3f0 (
.flogtanh_sel( Ie595a7d10b5ac84c0301fb55bebd3680[flogtanh_SEL-1:0]),
.flogtanh( Ie2ee6baf8ec357f6131dff92fb480e42),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ieddef08050c38d07e5d38f5bb7b099c0 = (Ie595a7d10b5ac84c0301fb55bebd3680[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie2ee6baf8ec357f6131dff92fb480e42;


Ic3da32f100a43f826b89a492544e7812 Ia42124b5528fdaa15431d0cc263861e1 (
.flogtanh_sel( I9c217a672cabc05efbdff218637123ba[flogtanh_SEL-1:0]),
.flogtanh( Ibff4d4fca3681fe10807414ed84e4157),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I39f9e8430db114991bfb27cc46ef3e39 = (I9c217a672cabc05efbdff218637123ba[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibff4d4fca3681fe10807414ed84e4157;


Ic3da32f100a43f826b89a492544e7812 I06aa4f71e36270bae01a1b3df5f0b54a (
.flogtanh_sel( If20f3780b4af857ffe8083056085517a[flogtanh_SEL-1:0]),
.flogtanh( I4540d74c919f50e9b6e40ef6b8cfd279),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I56aa548618a4a15e9a35e04f5eeb823f = (If20f3780b4af857ffe8083056085517a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4540d74c919f50e9b6e40ef6b8cfd279;


Ic3da32f100a43f826b89a492544e7812 Icbf90c5e62157ebb78cc42245533a57c (
.flogtanh_sel( Ic2e275bfa8ab3d2002d2aa374ac9bfe2[flogtanh_SEL-1:0]),
.flogtanh( I01637ffca829d72accbb5dcee48817ca),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I1908897b529ca04df7e7da395be4a8ce = (Ic2e275bfa8ab3d2002d2aa374ac9bfe2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I01637ffca829d72accbb5dcee48817ca;


Ic3da32f100a43f826b89a492544e7812 I73b2cbb8c6119d51ac07a1ea5b6db42c (
.flogtanh_sel( Iac5798fd9915b6778700da6a14f6a381[flogtanh_SEL-1:0]),
.flogtanh( I7e8af960e934c7cc3cb163d6f8e7d597),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib2bbd59cd6098608ed53ac556036534f = (Iac5798fd9915b6778700da6a14f6a381[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7e8af960e934c7cc3cb163d6f8e7d597;


Ic3da32f100a43f826b89a492544e7812 I484b5f5a8aed7a5e4925adda6278717c (
.flogtanh_sel( Ide3204bf317fdfb993410d338085b174[flogtanh_SEL-1:0]),
.flogtanh( Ifd80d371c8851b9e16193a3e62ddf79a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If004552b2047ab1cf23bb50375460b01 = (Ide3204bf317fdfb993410d338085b174[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifd80d371c8851b9e16193a3e62ddf79a;


Ic3da32f100a43f826b89a492544e7812 If5610dbdfd1b6a203d84c5c1be4ac7ab (
.flogtanh_sel( Ic3a95140fc1029efa17a6557bc977719[flogtanh_SEL-1:0]),
.flogtanh( I19d2c4bc969133fa59d22f7f2d8cfd4a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign If97092e1e2147de199c94a23831cf6b9 = (Ic3a95140fc1029efa17a6557bc977719[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I19d2c4bc969133fa59d22f7f2d8cfd4a;


Ic3da32f100a43f826b89a492544e7812 I6adee83776be48a034f8efd49058f45b (
.flogtanh_sel( I647d3a46bb2c7ed0f1ec08760b3858be[flogtanh_SEL-1:0]),
.flogtanh( I532326ad245909d441134296dae9a5d4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibf74a4dfaab7f7f538d2b5fac7394b63 = (I647d3a46bb2c7ed0f1ec08760b3858be[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I532326ad245909d441134296dae9a5d4;


Ic3da32f100a43f826b89a492544e7812 I590ce2649462d2b48875c2cfbfc42eac (
.flogtanh_sel( I4816747af9d9fc8dc85fd831336ec710[flogtanh_SEL-1:0]),
.flogtanh( I6ca7199e28b480ac5816bf5b4cfb1eef),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I991a7a7d562eb0a8b4b8d8f008ef2225 = (I4816747af9d9fc8dc85fd831336ec710[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I6ca7199e28b480ac5816bf5b4cfb1eef;


Ic3da32f100a43f826b89a492544e7812 I800be51fb0cb4ccded9a3fc790456adf (
.flogtanh_sel( I1f66c026a5437320bd1f4df2ff71663d[flogtanh_SEL-1:0]),
.flogtanh( I0d5b26d24fbce6b236120b5697d0db6b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I64c3d7be41abaa17d6992f9af8e72789 = (I1f66c026a5437320bd1f4df2ff71663d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0d5b26d24fbce6b236120b5697d0db6b;


Ic3da32f100a43f826b89a492544e7812 I74c0fe50913ae65ae65787eced04d41b (
.flogtanh_sel( If347c58c328193f420286ea27a4afa20[flogtanh_SEL-1:0]),
.flogtanh( I618d329f2b0f18617d80aa350b79601c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icb91e63ebabc7a75a54eb7c731df4fa0 = (If347c58c328193f420286ea27a4afa20[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I618d329f2b0f18617d80aa350b79601c;


Ic3da32f100a43f826b89a492544e7812 I17984729ee36ef800d16f9c734477932 (
.flogtanh_sel( I7a126c8304be920f2a920315dc61ba7f[flogtanh_SEL-1:0]),
.flogtanh( I58e3a5e842e14d09de91959839798a67),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I673d1d0d0daab99bd940c46cc14ef55a = (I7a126c8304be920f2a920315dc61ba7f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I58e3a5e842e14d09de91959839798a67;


Ic3da32f100a43f826b89a492544e7812 I64b3bbbe7bb8d13e7e92c2ab57368fcc (
.flogtanh_sel( I237327d6a74df1fb05537dc3691ebf11[flogtanh_SEL-1:0]),
.flogtanh( Icdecd5095ef818a0915ff3fcb395db5b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I62cadbd70b07a6a7a2974c7c392696b3 = (I237327d6a74df1fb05537dc3691ebf11[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Icdecd5095ef818a0915ff3fcb395db5b;


Ic3da32f100a43f826b89a492544e7812 I1f722d7ad9bb3b31da74bdbfa8818bac (
.flogtanh_sel( I64a3e8bb4c87b066806d33a5306a2c53[flogtanh_SEL-1:0]),
.flogtanh( I236f843994d3065b6ee70c41f390a3d0),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icd8257d7f53d93db989eb56eaeb7e593 = (I64a3e8bb4c87b066806d33a5306a2c53[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I236f843994d3065b6ee70c41f390a3d0;


Ic3da32f100a43f826b89a492544e7812 I98f966db853a11ffc1315494ce32395f (
.flogtanh_sel( Ibbca6ec39234473fb517447a8beacafc[flogtanh_SEL-1:0]),
.flogtanh( I7a9001d6c1d1aa8af79d9b152e596b70),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I05931ceae6eff26e5a66a44a54d628ae = (Ibbca6ec39234473fb517447a8beacafc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7a9001d6c1d1aa8af79d9b152e596b70;


Ic3da32f100a43f826b89a492544e7812 Ifdff296113f028882cd9e18e5578fe0d (
.flogtanh_sel( I78327356176a16fc996188b83b058cbc[flogtanh_SEL-1:0]),
.flogtanh( I56a43a072d463792d9e676c4907b3e76),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I306fec0aa68a0396053a6e0fa1cda38f = (I78327356176a16fc996188b83b058cbc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I56a43a072d463792d9e676c4907b3e76;


Ic3da32f100a43f826b89a492544e7812 Ie057aed9b8d76278f08c087868f09c4b (
.flogtanh_sel( Ifec496c87a7a2474855067305ac8cba3[flogtanh_SEL-1:0]),
.flogtanh( I336a86e85d3a8a42c4b6458ccb92ae05),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Idee8c8144207d676d1f2f9064bbdff45 = (Ifec496c87a7a2474855067305ac8cba3[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I336a86e85d3a8a42c4b6458ccb92ae05;


Ic3da32f100a43f826b89a492544e7812 Ia018b862c11a378b644bf40310b72df2 (
.flogtanh_sel( I41584165a62caaa37ddebbf79bb8b617[flogtanh_SEL-1:0]),
.flogtanh( Id97f66b78f1e3b6bf0b962b85ca1cde7),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5855124d566af739caa6511f8598f2c5 = (I41584165a62caaa37ddebbf79bb8b617[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id97f66b78f1e3b6bf0b962b85ca1cde7;


Ic3da32f100a43f826b89a492544e7812 I47230e65145ef951045032cce4c551cc (
.flogtanh_sel( Idf0916d6b025aad6eccb98ada5ba3aca[flogtanh_SEL-1:0]),
.flogtanh( I52c7f0a8f9b4533052b5acd1b5bd5e17),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I50729db4a8e04f18979707df14cb2419 = (Idf0916d6b025aad6eccb98ada5ba3aca[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I52c7f0a8f9b4533052b5acd1b5bd5e17;


Ic3da32f100a43f826b89a492544e7812 I77e98518151a4480bab54df6712c8b3d (
.flogtanh_sel( I00ef133d5a53f8f99f35b50327e5272b[flogtanh_SEL-1:0]),
.flogtanh( I3b1db672b1a94502b90451260062a274),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia3cb3ea64576a3e7332e1fb55953aa3e = (I00ef133d5a53f8f99f35b50327e5272b[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I3b1db672b1a94502b90451260062a274;


Ic3da32f100a43f826b89a492544e7812 Iccf5cb35860f9ebea1366f27ddc4983b (
.flogtanh_sel( I6f0e302d38d75982d0761e306ce9f146[flogtanh_SEL-1:0]),
.flogtanh( I1a83f91eb1262911ae8d99e305294bf8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I3cb1f233951d49f985b0deac6e052bfd = (I6f0e302d38d75982d0761e306ce9f146[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I1a83f91eb1262911ae8d99e305294bf8;


Ic3da32f100a43f826b89a492544e7812 I0ac462f33956122486bc7b6ae9a730dc (
.flogtanh_sel( I127eed5de00e10a020717e796de76c7d[flogtanh_SEL-1:0]),
.flogtanh( Id01bfbd86b6321a843e239ca97cec514),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7015def91103398e54f446ce3e43af01 = (I127eed5de00e10a020717e796de76c7d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Id01bfbd86b6321a843e239ca97cec514;


Ic3da32f100a43f826b89a492544e7812 Ib0b64a4b4d9899bdb008b5a24f321373 (
.flogtanh_sel( If9aad73aefb1b225f35e8c813b85fe87[flogtanh_SEL-1:0]),
.flogtanh( I26b769b58e1c21b68dd95c9f38c0362b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I04874bd1bf257f205b5189c8c20e5a12 = (If9aad73aefb1b225f35e8c813b85fe87[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I26b769b58e1c21b68dd95c9f38c0362b;


Ic3da32f100a43f826b89a492544e7812 Iea9fd1dae1f890f371990759b117ed16 (
.flogtanh_sel( I00a89ac37676521a081a21b1ec1a0798[flogtanh_SEL-1:0]),
.flogtanh( Ic86f9988281398adfe43152beb722c1b),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I937e3a8ede2305ea7c1750283224a870 = (I00a89ac37676521a081a21b1ec1a0798[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic86f9988281398adfe43152beb722c1b;


Ic3da32f100a43f826b89a492544e7812 Ifbeaf32038f3cf22265f0bc1fef1ffd6 (
.flogtanh_sel( I06f3a34f2b1770ef82ddc2a732b3d4fb[flogtanh_SEL-1:0]),
.flogtanh( I9d8ac6c29c2f5df7c2d124dface59e35),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia7206430a739a11af4d860096eedd6c3 = (I06f3a34f2b1770ef82ddc2a732b3d4fb[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9d8ac6c29c2f5df7c2d124dface59e35;


Ic3da32f100a43f826b89a492544e7812 Ic8da88c0920636e001dd2138f21ec58f (
.flogtanh_sel( I4744d64a746f16004e3bedaaa41465f1[flogtanh_SEL-1:0]),
.flogtanh( I56b46c426895409b40c3be9b79365a8a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ibf4c2c00f8e012e9498361bfd3c5b06e = (I4744d64a746f16004e3bedaaa41465f1[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I56b46c426895409b40c3be9b79365a8a;


Ic3da32f100a43f826b89a492544e7812 I3653f33d698a22202ee2975e51101454 (
.flogtanh_sel( Ifae0cc6cc1c65d24bbe84c4ba938e2ea[flogtanh_SEL-1:0]),
.flogtanh( Ic63de8464f79ae05f27f05c935dbf495),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I899e5f03cd1d52d11f898959559aaeea = (Ifae0cc6cc1c65d24bbe84c4ba938e2ea[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ic63de8464f79ae05f27f05c935dbf495;


Ic3da32f100a43f826b89a492544e7812 Ic1c122d700eb5e9fa61c842b1336e9a6 (
.flogtanh_sel( I1223c21129382d41e4f38ef4bbe60c2f[flogtanh_SEL-1:0]),
.flogtanh( I4d21ee443e5921532d5bf1db7ef93f82),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I59c80c7ec26f43308b1a646c47160568 = (I1223c21129382d41e4f38ef4bbe60c2f[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I4d21ee443e5921532d5bf1db7ef93f82;


Ic3da32f100a43f826b89a492544e7812 Iba5c6c5ca1c5d08b54928848ef1fa8a4 (
.flogtanh_sel( I14e36e16df00adcd7dc1973d3852d2d9[flogtanh_SEL-1:0]),
.flogtanh( Ieb5fa20abbdb29a7f75021b7afafea31),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8a954a331d36266465a0813d2e8b319b = (I14e36e16df00adcd7dc1973d3852d2d9[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ieb5fa20abbdb29a7f75021b7afafea31;


Ic3da32f100a43f826b89a492544e7812 I09feb8ce383e6bab74488a905cd089b2 (
.flogtanh_sel( I0d05ae27b53fb6939e4c2f862a8d20b2[flogtanh_SEL-1:0]),
.flogtanh( I16a12326344aadf4226bd149424a53a8),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ib49e53ca8efd9564ee9572eb3089bb51 = (I0d05ae27b53fb6939e4c2f862a8d20b2[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I16a12326344aadf4226bd149424a53a8;


Ic3da32f100a43f826b89a492544e7812 I19213cf4ab1c0a3ad1ed011733930a4c (
.flogtanh_sel( I97a6fcc08929c3b7d15e36d7706ed13d[flogtanh_SEL-1:0]),
.flogtanh( I07f36b533b48344c13dbb133739712f4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icbde2c6230e9cc67ef12031e38bb344f = (I97a6fcc08929c3b7d15e36d7706ed13d[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I07f36b533b48344c13dbb133739712f4;


Ic3da32f100a43f826b89a492544e7812 Ie1d3b883db1f997cc3af7579b482a0bc (
.flogtanh_sel( I1f04e86bf27596718836d0a09adbe120[flogtanh_SEL-1:0]),
.flogtanh( I7a0072bf1e5fb0c4de85c6e4447878a4),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I2e22e867f6f84a7807b82f64a147022e = (I1f04e86bf27596718836d0a09adbe120[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I7a0072bf1e5fb0c4de85c6e4447878a4;


Ic3da32f100a43f826b89a492544e7812 I8e6a22f10221bcce6f782c111c5f099e (
.flogtanh_sel( Ie40873cfd6d10a61a94a761becf588a8[flogtanh_SEL-1:0]),
.flogtanh( I320bafc5a1775d6933bcb9f2d2c84576),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id9704e1d8096cd28577c5c357d30b7a4 = (Ie40873cfd6d10a61a94a761becf588a8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I320bafc5a1775d6933bcb9f2d2c84576;


Ic3da32f100a43f826b89a492544e7812 I18a4d6265272844e1a82ecca75149855 (
.flogtanh_sel( I61960ed74fee948cc12bd1fd8384559a[flogtanh_SEL-1:0]),
.flogtanh( I5ec61756ff7237146f2d83f17eb5bb3a),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I4b8554cab486a4fc1e14884a6495016e = (I61960ed74fee948cc12bd1fd8384559a[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I5ec61756ff7237146f2d83f17eb5bb3a;


Ic3da32f100a43f826b89a492544e7812 Ia36e6aef2ad801d0706f3626ba2ad29d (
.flogtanh_sel( I8533a3ec4be4c49166184c94761eaebc[flogtanh_SEL-1:0]),
.flogtanh( I382008a17338641e68fa859ac2af1d20),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Iaa235d085a5916a3b0814c3ed2a9026f = (I8533a3ec4be4c49166184c94761eaebc[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I382008a17338641e68fa859ac2af1d20;


Ic3da32f100a43f826b89a492544e7812 If338259da548afa8039e769b4f9fece0 (
.flogtanh_sel( I00be319b5bdb85ffaf3bb0eca0b348b6[flogtanh_SEL-1:0]),
.flogtanh( Ifd375ad8038ea2455c0e3b1463b83b7e),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I5d86ce0b58c0b281d747116a9069ef33 = (I00be319b5bdb85ffaf3bb0eca0b348b6[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ifd375ad8038ea2455c0e3b1463b83b7e;


Ic3da32f100a43f826b89a492544e7812 Ic0ec1dc21242d0b4f2eb446ea5bf4ac9 (
.flogtanh_sel( Ie889c916b5af185b52ff5e2e3cc23045[flogtanh_SEL-1:0]),
.flogtanh( I0b75763235278d8eca6ca72fc97fb83c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Id20394136fb036435bb4680aac64581f = (Ie889c916b5af185b52ff5e2e3cc23045[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I0b75763235278d8eca6ca72fc97fb83c;


Ic3da32f100a43f826b89a492544e7812 Idd47130227196af1c07824f261960777 (
.flogtanh_sel( I89697be6dcb2e7f972db498c1b1dea71[flogtanh_SEL-1:0]),
.flogtanh( I9bc4c3b77a9635bb77ad31527d961952),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I8a16afac6e470ca69634d7fe9656387a = (I89697be6dcb2e7f972db498c1b1dea71[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I9bc4c3b77a9635bb77ad31527d961952;


Ic3da32f100a43f826b89a492544e7812 Ica2c981f339f1837ef80d00ff8719f8d (
.flogtanh_sel( If13dfbfff7cd8e197bb44006a3db73bf[flogtanh_SEL-1:0]),
.flogtanh( Ief93f4a7eaaa1f43ea1788dc4629c093),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic4e7f690bc050f1d1f84eae7ca193e1c = (If13dfbfff7cd8e197bb44006a3db73bf[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ief93f4a7eaaa1f43ea1788dc4629c093;


Ic3da32f100a43f826b89a492544e7812 I68832efe84de3f0982aef3f0350d39a2 (
.flogtanh_sel( I87ed6c3e172c7a06bf6aefe7bf718d70[flogtanh_SEL-1:0]),
.flogtanh( I34b86fbc3949cb2083931ad8edd2444d),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ia60421aa427236540b4d0d08d52ff507 = (I87ed6c3e172c7a06bf6aefe7bf718d70[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I34b86fbc3949cb2083931ad8edd2444d;


Ic3da32f100a43f826b89a492544e7812 Ib918e22f494b7c6cbcc11de46b4ea7c5 (
.flogtanh_sel( I0db87adc849839fab3a4c9884d5a4882[flogtanh_SEL-1:0]),
.flogtanh( I560c163fb55aa4b56da25f96e9b8ef6c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Icace650ee3865bd7bbddd2d9435c5561 = (I0db87adc849839fab3a4c9884d5a4882[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: I560c163fb55aa4b56da25f96e9b8ef6c;


Ic3da32f100a43f826b89a492544e7812 I73aa7f9c7931e07bafbeb5d388fe5cb8 (
.flogtanh_sel( I535e01a6c35fd7b455e4b79b1d4bb414[flogtanh_SEL-1:0]),
.flogtanh( Ib3c46d34c5bc3d2651147b3e764d9786),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I7d27d070b96b7810f667e1d1845342d3 = (I535e01a6c35fd7b455e4b79b1d4bb414[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ib3c46d34c5bc3d2651147b3e764d9786;


Ic3da32f100a43f826b89a492544e7812 Ib53b3683f37f4f1bf8f229753614a4be (
.flogtanh_sel( Ia2d1c752cc4b405adb97a815e90a7b96[flogtanh_SEL-1:0]),
.flogtanh( Ie5e2ba4fe22870afc81d6cfc708570be),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ida7ec09c913caa0e78a2c4cbaae517c8 = (Ia2d1c752cc4b405adb97a815e90a7b96[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ie5e2ba4fe22870afc81d6cfc708570be;


Ic3da32f100a43f826b89a492544e7812 Ib17b7f7a1fa4c71953f2144b8d877ed4 (
.flogtanh_sel( I9ac12eb3878f6fc7dc428fe5e7f35d97[flogtanh_SEL-1:0]),
.flogtanh( Ibf3bde181da4f960537516d6c0b2a72c),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign Ic5eba898858be1f768841ead792d6d86 = (I9ac12eb3878f6fc7dc428fe5e7f35d97[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ibf3bde181da4f960537516d6c0b2a72c;


Ic3da32f100a43f826b89a492544e7812 I11e8ec581a95e2705add61f3afefebb1 (
.flogtanh_sel( If46fa11dfadb0691eaaa0a40836e08d8[flogtanh_SEL-1:0]),
.flogtanh( Ia93f96aa0718f8755e9ebb8cc5d8f405),
.start_in(I699819696b0299ab80e7233d054ec590),
.start_out(),
.rstn(rstn),
.clk(clk)
);

assign I72197797a307c611fa8952533e63d7bf = (If46fa11dfadb0691eaaa0a40836e08d8[MAX_SUM_WDTH:0] > flogtanh_LEN ) ? 'h0: Ia93f96aa0718f8755e9ebb8cc5d8f405;





Ic9c2f173881d25f8976d723957809f51 Ied1ef1f3c0fd7afaae5baa9cfe2a2535 (
.fgallag_sel( I97afe24956b7f87cd431f048202bab67[fgallag_SEL-1:0]),
.fgallag( Ic188ebb37ff178022c61400613f4f3dc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(I92354deea988f3beb25bfba90735c6ac),
.rstn(rstn),
.clk(clk)
);


assign I5a11c8e7d2b7d4c0253df9015b7f3ab5 = (I97afe24956b7f87cd431f048202bab67[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic188ebb37ff178022c61400613f4f3dc ;

Ic9c2f173881d25f8976d723957809f51 Ibc2fcc821b2425084cbdd233159fc006 (
.fgallag_sel( I117235e3ac8e68e4c1ab34db1612aba0[fgallag_SEL-1:0]),
.fgallag( I3f80921fd94cff373648fa34fcadd4d2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib0740d8c9ab158e682432a0e3ec89798 = (I117235e3ac8e68e4c1ab34db1612aba0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3f80921fd94cff373648fa34fcadd4d2 ;

Ic9c2f173881d25f8976d723957809f51 I5806029f24210308e5ef5f73b9b8bcac (
.fgallag_sel( Ifd700cc9d18f99b63f1947f3ae631976[fgallag_SEL-1:0]),
.fgallag( I229f7430f590d86a323b48806beec48c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibb6505392d5b3be76542bb0303d46876 = (Ifd700cc9d18f99b63f1947f3ae631976[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I229f7430f590d86a323b48806beec48c ;

Ic9c2f173881d25f8976d723957809f51 Ic8daf8ffe06d27a0c84083675507c938 (
.fgallag_sel( Ifffbe3d1007fb07a20d3b37902b3ec95[fgallag_SEL-1:0]),
.fgallag( I26fa0a5f87600d9535e8f83fa1a11136 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If23edf1bc3801016b24252fbc3d33508 = (Ifffbe3d1007fb07a20d3b37902b3ec95[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I26fa0a5f87600d9535e8f83fa1a11136 ;

Ic9c2f173881d25f8976d723957809f51 I3cc84bed6b0b1ac3206b3ee03f637fd2 (
.fgallag_sel( If5443777169422ea6e1e3f709b970e05[fgallag_SEL-1:0]),
.fgallag( Id87360986474c9bfa5266a90b59a9a8b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I47478ccbfc4c3b944d130a192fb4fb5a = (If5443777169422ea6e1e3f709b970e05[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id87360986474c9bfa5266a90b59a9a8b ;

Ic9c2f173881d25f8976d723957809f51 I3abcbe1f5f69abcfd50f7e9b4c6faa74 (
.fgallag_sel( Ifaf9fc93e4609d818aa46751754c17f1[fgallag_SEL-1:0]),
.fgallag( Id63daaeb52208682533b5f136480a29c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I40b126fdab110e58eac80ea13bcc699d = (Ifaf9fc93e4609d818aa46751754c17f1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id63daaeb52208682533b5f136480a29c ;

Ic9c2f173881d25f8976d723957809f51 I1152f0e84d9368eebc9b2c8770ff87c2 (
.fgallag_sel( I419caf964986c655df84d043badc37c9[fgallag_SEL-1:0]),
.fgallag( I1e9d5c2338b6f89e43c30c0ad71f675c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib12b389fb2603e428b72d1e712975e40 = (I419caf964986c655df84d043badc37c9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1e9d5c2338b6f89e43c30c0ad71f675c ;

Ic9c2f173881d25f8976d723957809f51 I8b9fe3036e2359699b0a458ba95a3ca9 (
.fgallag_sel( I3095214ac0e6c1323e75ee4ec85e6821[fgallag_SEL-1:0]),
.fgallag( I11cce7dd119eb0e3acafc12dbc6d3536 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I22b0cc5517631526be6455fc60dd5323 = (I3095214ac0e6c1323e75ee4ec85e6821[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I11cce7dd119eb0e3acafc12dbc6d3536 ;

Ic9c2f173881d25f8976d723957809f51 I4278d8aa5885a75a34ad1408d5ca8702 (
.fgallag_sel( Ided9739bf63937933250a6d0c37535f9[fgallag_SEL-1:0]),
.fgallag( I934b111c08439d3797cb8928c7238f23 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib8aba28214fb9ee1693cafe9175831e1 = (Ided9739bf63937933250a6d0c37535f9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I934b111c08439d3797cb8928c7238f23 ;

Ic9c2f173881d25f8976d723957809f51 I65e82922c9e54f9b79654d55a0900b47 (
.fgallag_sel( Id0f139b9f3848b45554ac8429230eea2[fgallag_SEL-1:0]),
.fgallag( I508cb12fa71441b216fd7c1899d00e24 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia03282a7ed4a337981d4f5b01f564a1d = (Id0f139b9f3848b45554ac8429230eea2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I508cb12fa71441b216fd7c1899d00e24 ;

Ic9c2f173881d25f8976d723957809f51 Ib5c646ad9dd6fee826088018930d8c50 (
.fgallag_sel( Id9feed58cf9565255abfd0bf7e3ec068[fgallag_SEL-1:0]),
.fgallag( Ic69c6ea6b4f360efae87611c00b00fdb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icf75bf863d8867b0fe354017921aeae1 = (Id9feed58cf9565255abfd0bf7e3ec068[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic69c6ea6b4f360efae87611c00b00fdb ;

Ic9c2f173881d25f8976d723957809f51 Ifee02b093e011b8bcd51f9c8a8829aa6 (
.fgallag_sel( I30a3be3b5f6ad1880a917eb35659a1bf[fgallag_SEL-1:0]),
.fgallag( Ifccbe59b7ebe3f692f5b7e7564ca50ba ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia65c174738acf41b82f75be972e9022e = (I30a3be3b5f6ad1880a917eb35659a1bf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifccbe59b7ebe3f692f5b7e7564ca50ba ;

Ic9c2f173881d25f8976d723957809f51 Ia8fa310f0c568cf154b2b8f559820f2a (
.fgallag_sel( Ie8148d9aa962a733eb65877b902a187d[fgallag_SEL-1:0]),
.fgallag( Ifd7275bc534fe9da81b12b25ed218e91 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I587a0e70cecf4d054cc0ab53150876e0 = (Ie8148d9aa962a733eb65877b902a187d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifd7275bc534fe9da81b12b25ed218e91 ;

Ic9c2f173881d25f8976d723957809f51 I5440a65550974852174a86b5e70cee47 (
.fgallag_sel( I69e98cf3e679183aef6005bb582b18dc[fgallag_SEL-1:0]),
.fgallag( I01a99ac2a3f919f4fc1680edb11c576b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7dc71f64f9b3940721569574db6e18d0 = (I69e98cf3e679183aef6005bb582b18dc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I01a99ac2a3f919f4fc1680edb11c576b ;

Ic9c2f173881d25f8976d723957809f51 I14093343f32180181772e04daefd0a13 (
.fgallag_sel( I7f42a504fc61c9548acebdd8b1858eaa[fgallag_SEL-1:0]),
.fgallag( I322b3879383d75c43c55535f01fdfdd6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I935ba9f8f6e9c68f75a7cb576655cab5 = (I7f42a504fc61c9548acebdd8b1858eaa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I322b3879383d75c43c55535f01fdfdd6 ;

Ic9c2f173881d25f8976d723957809f51 I2b9c5d47f848188a8010a80c74e9b86d (
.fgallag_sel( I08b1b4639b5a9ca509b943b977f6d4bb[fgallag_SEL-1:0]),
.fgallag( I1adc689464e0b81fa165eb17e71310fa ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibdc981a062c989ada978f733ddff0f71 = (I08b1b4639b5a9ca509b943b977f6d4bb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1adc689464e0b81fa165eb17e71310fa ;

Ic9c2f173881d25f8976d723957809f51 Ic93034cd51979700d51babca220be23f (
.fgallag_sel( I8d7296627d886566783e79c01b9fa423[fgallag_SEL-1:0]),
.fgallag( I2bdc0908c3d365d25f8026263dc4a258 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibcbc5e2720516c24359870ac790373f4 = (I8d7296627d886566783e79c01b9fa423[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2bdc0908c3d365d25f8026263dc4a258 ;

Ic9c2f173881d25f8976d723957809f51 I2e95bba468c48cceb71f006dbf06eece (
.fgallag_sel( I4fc4c97229a8b1f631a3b505941159e4[fgallag_SEL-1:0]),
.fgallag( Icf6c6fcfa42c48f16a1b30cd325c139f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I11fdefe51f8f028fba7698870d198df6 = (I4fc4c97229a8b1f631a3b505941159e4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Icf6c6fcfa42c48f16a1b30cd325c139f ;

Ic9c2f173881d25f8976d723957809f51 I7b2eed1152ba088b207fba7450885f43 (
.fgallag_sel( Ib9b16bf51891c328dba2699eb9bcef95[fgallag_SEL-1:0]),
.fgallag( Ife8337f33629521c096d4dcfde96e879 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I10f17104471f87c53a589926534fc9fe = (Ib9b16bf51891c328dba2699eb9bcef95[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ife8337f33629521c096d4dcfde96e879 ;

Ic9c2f173881d25f8976d723957809f51 I29a34e3f98c0bd69e7aa9204f49033a9 (
.fgallag_sel( I6c30501ec81fce286817788d614a7824[fgallag_SEL-1:0]),
.fgallag( I8afa93d48ae589bb90cc74897defe4de ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8fdaa3f282af2d5f053d77216c659146 = (I6c30501ec81fce286817788d614a7824[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8afa93d48ae589bb90cc74897defe4de ;

Ic9c2f173881d25f8976d723957809f51 Ic9617b2e89efcaa4c8249a287af21871 (
.fgallag_sel( Ia4d4f37baec48121a88808075dd655ef[fgallag_SEL-1:0]),
.fgallag( I56d0b4df55f7f4181a51f58187d399e4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I167ee185ac7beee082544897898b27fa = (Ia4d4f37baec48121a88808075dd655ef[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I56d0b4df55f7f4181a51f58187d399e4 ;

Ic9c2f173881d25f8976d723957809f51 I98ce0bdc7e2b3a205ed054ce747546bf (
.fgallag_sel( I385495ea2bf6442a95ab7561456254ac[fgallag_SEL-1:0]),
.fgallag( I8ae9260d2a5dd6c2ed4b6157946e38d4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5264a25f96edda24a763298d92cdf8c1 = (I385495ea2bf6442a95ab7561456254ac[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8ae9260d2a5dd6c2ed4b6157946e38d4 ;

Ic9c2f173881d25f8976d723957809f51 I4f99d5a9644e17aca23a8d33e54ba1b8 (
.fgallag_sel( I5128e03d383c226befa6f7422f3a6f04[fgallag_SEL-1:0]),
.fgallag( Ie405c3459c9caf16c0a257a059a9fa96 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If7d5260450e23711760a6f9e5f7aa820 = (I5128e03d383c226befa6f7422f3a6f04[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie405c3459c9caf16c0a257a059a9fa96 ;

Ic9c2f173881d25f8976d723957809f51 Ibe41e6cd8796984537c236df29203e77 (
.fgallag_sel( Ib208908bab4c20713cd17e20139c8db3[fgallag_SEL-1:0]),
.fgallag( Ie76a46f18cbb52a93a4fad65462da3e8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id1265b30a8ed85169b1837aa1b656aa2 = (Ib208908bab4c20713cd17e20139c8db3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie76a46f18cbb52a93a4fad65462da3e8 ;

Ic9c2f173881d25f8976d723957809f51 I5a98b7e432b5508f70b55fdcb502e832 (
.fgallag_sel( Id939992b99a11c09f4688c10ca1a34d1[fgallag_SEL-1:0]),
.fgallag( I0445dbe40692ef21353aacc7b4f7a4c9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I84e6c5099aaef8094f4c2bbc82989c4c = (Id939992b99a11c09f4688c10ca1a34d1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0445dbe40692ef21353aacc7b4f7a4c9 ;

Ic9c2f173881d25f8976d723957809f51 I4833867123384374e5fd034e6629c018 (
.fgallag_sel( I823453ccb90d5b2b2d9dfc6e8358224d[fgallag_SEL-1:0]),
.fgallag( Ie3be0f770c8ddbdf301ae23881499e9d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibf4bfa16424f7051e80b2947ff7f5533 = (I823453ccb90d5b2b2d9dfc6e8358224d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie3be0f770c8ddbdf301ae23881499e9d ;

Ic9c2f173881d25f8976d723957809f51 Iab4ce39770acfed571965352cae92c10 (
.fgallag_sel( I279c5c00b92eb1b872b5afa168b0306e[fgallag_SEL-1:0]),
.fgallag( I3a4d175e3b015a17f7a49cc6bacbd12f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0e138642d8ed7e30cc254d4e259e3d51 = (I279c5c00b92eb1b872b5afa168b0306e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3a4d175e3b015a17f7a49cc6bacbd12f ;

Ic9c2f173881d25f8976d723957809f51 I59fe58ec0aa6b1d27afa73271aa0983b (
.fgallag_sel( I66f25b1c3c0eb226295179adcca2c3d2[fgallag_SEL-1:0]),
.fgallag( Id85473220f4909f9182711939cf6a978 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If1c79ab7bbf50d343ba3f758a31d6786 = (I66f25b1c3c0eb226295179adcca2c3d2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id85473220f4909f9182711939cf6a978 ;

Ic9c2f173881d25f8976d723957809f51 I82ed432dbb156e795df7eb7edddbc6ac (
.fgallag_sel( I3068627e91b667d14cd3e55a9371931a[fgallag_SEL-1:0]),
.fgallag( If77ecdb29d692c01752be0908c4f4392 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic2d209d919c7e43f467c3f2d093c9a8c = (I3068627e91b667d14cd3e55a9371931a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If77ecdb29d692c01752be0908c4f4392 ;

Ic9c2f173881d25f8976d723957809f51 I0fa2411ae78a94b20b3cce85ab19110d (
.fgallag_sel( I44c4e0a2d8a7289f8660b81a9ecfa19b[fgallag_SEL-1:0]),
.fgallag( Ia188482ea4a2696f188f637912aa6f3b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6c59651ae65c67edfa963ce797b98234 = (I44c4e0a2d8a7289f8660b81a9ecfa19b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia188482ea4a2696f188f637912aa6f3b ;

Ic9c2f173881d25f8976d723957809f51 If89e681d9340e16014cdf269d3eb81e5 (
.fgallag_sel( Ibe868e258dc87f0dd1460ba6b8354671[fgallag_SEL-1:0]),
.fgallag( Ibd0c9231ee029200ca39013c839bc4ae ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If4b95101c6d8670411a018ed1ae697d3 = (Ibe868e258dc87f0dd1460ba6b8354671[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibd0c9231ee029200ca39013c839bc4ae ;

Ic9c2f173881d25f8976d723957809f51 Idbad8b20599f8ec1979606226040e4de (
.fgallag_sel( Idc3083c3021200345e3edd35a9d4725a[fgallag_SEL-1:0]),
.fgallag( I0fed2eb07a75f701ff7b7ca9dbcddb81 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib1e406a5bb0569ac2c25e7021ec58edb = (Idc3083c3021200345e3edd35a9d4725a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0fed2eb07a75f701ff7b7ca9dbcddb81 ;

Ic9c2f173881d25f8976d723957809f51 I16ce3220cd54730858727d5693dfd447 (
.fgallag_sel( I320d4f19a5b18c23ff407508d47caa77[fgallag_SEL-1:0]),
.fgallag( I96140f2ad00cb9a1249b5135ea251bc8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8198f75286b8c817d3b69cf7537b1c38 = (I320d4f19a5b18c23ff407508d47caa77[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I96140f2ad00cb9a1249b5135ea251bc8 ;

Ic9c2f173881d25f8976d723957809f51 Ie59e1b18dcb4f2d35a9c7c9238743f1b (
.fgallag_sel( I16becf3c92615d98d5ec51ee9641cc0a[fgallag_SEL-1:0]),
.fgallag( I34fecbd6c558b25e7f8d08fb10b224f4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9431b10311eda8240d91bed96a969523 = (I16becf3c92615d98d5ec51ee9641cc0a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I34fecbd6c558b25e7f8d08fb10b224f4 ;

Ic9c2f173881d25f8976d723957809f51 I81035565ff539fd780f9c7c8c8597463 (
.fgallag_sel( Ifbfacc3b3a0128119943bcbf80176612[fgallag_SEL-1:0]),
.fgallag( I8df49bd85a846a4c4c32af63798f3e0e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib623d99c3d272f39c518b6a41dd03e8d = (Ifbfacc3b3a0128119943bcbf80176612[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8df49bd85a846a4c4c32af63798f3e0e ;

Ic9c2f173881d25f8976d723957809f51 I64f946de094aaf688c4cb8c8e73d5c90 (
.fgallag_sel( I6b4f670c9e8e25984e8891f2440322ab[fgallag_SEL-1:0]),
.fgallag( I05be7b5c657867c4331ed3df72a1aec5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I388b66a7b7e9225f7aef4699521e9250 = (I6b4f670c9e8e25984e8891f2440322ab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I05be7b5c657867c4331ed3df72a1aec5 ;

Ic9c2f173881d25f8976d723957809f51 I977ee6c9fa86dddbfcd2f944fc40a0af (
.fgallag_sel( I19bf0990a30c72421f231772b8627e8e[fgallag_SEL-1:0]),
.fgallag( Id47eecb4e17f799da48d80451cb47b5d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I532db075ab1b0a5a37a2085ecd0611c3 = (I19bf0990a30c72421f231772b8627e8e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id47eecb4e17f799da48d80451cb47b5d ;

Ic9c2f173881d25f8976d723957809f51 Iee4a23ecb4c40c373f84bbb4554db60e (
.fgallag_sel( I3ec3eb096ebe3ee8a47e1cba6487b997[fgallag_SEL-1:0]),
.fgallag( Iedabb8b1ffd46b983fd74b9f6010dcca ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I357c21c29061134ed6e5c872836f4759 = (I3ec3eb096ebe3ee8a47e1cba6487b997[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iedabb8b1ffd46b983fd74b9f6010dcca ;

Ic9c2f173881d25f8976d723957809f51 I458334bece48070d9cc3926b2e7a87a3 (
.fgallag_sel( I7379ef16405c461ac44b66c4315df831[fgallag_SEL-1:0]),
.fgallag( Ib032a08190a75ceb242a9dc8272b4a02 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5a1d671b8b8877192d2c129be7f149c0 = (I7379ef16405c461ac44b66c4315df831[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib032a08190a75ceb242a9dc8272b4a02 ;

Ic9c2f173881d25f8976d723957809f51 I3be4f1a4643508e1855f0a2585cfcb4c (
.fgallag_sel( I79db45b23d21d533a1f9a6e8f94d403d[fgallag_SEL-1:0]),
.fgallag( Ia870db84a0411e463b6e15f502323810 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4d1c830053fedd74930d9992732e9542 = (I79db45b23d21d533a1f9a6e8f94d403d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia870db84a0411e463b6e15f502323810 ;

Ic9c2f173881d25f8976d723957809f51 Id996909c05c3e6244ab67893f03f9bdd (
.fgallag_sel( I0979534730cc2b53547d413dbb6b75f4[fgallag_SEL-1:0]),
.fgallag( I8105600a0847cabdb96310074840bdb7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie53c31ded4a5c8977f956e968dd5a9a7 = (I0979534730cc2b53547d413dbb6b75f4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8105600a0847cabdb96310074840bdb7 ;

Ic9c2f173881d25f8976d723957809f51 I50be605a6015a779d5fc652a3833aad0 (
.fgallag_sel( I5aa2f9c0667d1a6e871efbd4d2bad3a8[fgallag_SEL-1:0]),
.fgallag( I7d6591184fd95d3f288f481734e85c02 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id5355c3ed75d1aed52250f6f0d00b1a0 = (I5aa2f9c0667d1a6e871efbd4d2bad3a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7d6591184fd95d3f288f481734e85c02 ;

Ic9c2f173881d25f8976d723957809f51 Ib5a6232daf646272f8fa545a8762473b (
.fgallag_sel( Iadb28dc990ccf2dd3099544de16b8f16[fgallag_SEL-1:0]),
.fgallag( I69c3d2866b040d67900eeb991b7c2981 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib43ca9d864e41a89bec5344ece17fd10 = (Iadb28dc990ccf2dd3099544de16b8f16[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I69c3d2866b040d67900eeb991b7c2981 ;

Ic9c2f173881d25f8976d723957809f51 I602e86d151abd3248add4b18a4047f4c (
.fgallag_sel( I1f71aebf698788d6ada66891e9ea756f[fgallag_SEL-1:0]),
.fgallag( Ice61d34abe5e2a9593bfb911da54e959 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6c7b0be00e8302794aa3a79fb2acf100 = (I1f71aebf698788d6ada66891e9ea756f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ice61d34abe5e2a9593bfb911da54e959 ;

Ic9c2f173881d25f8976d723957809f51 I9667284df1deac69373fc5e85e49fe76 (
.fgallag_sel( Ib234e9cf7e7616a1ebc6ab99df2a7ccb[fgallag_SEL-1:0]),
.fgallag( I7dfe4eb1588a68b8a35dec39978d06eb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I144843095a5e8952e26bb5c9943f0cad = (Ib234e9cf7e7616a1ebc6ab99df2a7ccb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7dfe4eb1588a68b8a35dec39978d06eb ;

Ic9c2f173881d25f8976d723957809f51 I335d0c659ee1d77669565d6c8d702258 (
.fgallag_sel( I297d1edcc583ea4d69da780150f0620c[fgallag_SEL-1:0]),
.fgallag( Ica59cc444ecf8f8700bf1ce16a254b89 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0b6cd5372e2cc6a72c1c8f984279cb69 = (I297d1edcc583ea4d69da780150f0620c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ica59cc444ecf8f8700bf1ce16a254b89 ;

Ic9c2f173881d25f8976d723957809f51 I5dd2edd850e50fb4cafeabf124c7354d (
.fgallag_sel( Ib0a717cbb4fe38a3fc85520ca0826fd9[fgallag_SEL-1:0]),
.fgallag( I0d69f1eb92a8b30d86ffbe0c153197f2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icd143823913eb777c0cba42d8a5802e9 = (Ib0a717cbb4fe38a3fc85520ca0826fd9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0d69f1eb92a8b30d86ffbe0c153197f2 ;

Ic9c2f173881d25f8976d723957809f51 I1b4d968802db0e9dcd2916ac527315ea (
.fgallag_sel( I037ecd5945b1f1280b4469d73fe1c7ff[fgallag_SEL-1:0]),
.fgallag( I5a48ea253b357c8e6441be01918bc57c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I02a575305a6112f734bc3ebf6b883b90 = (I037ecd5945b1f1280b4469d73fe1c7ff[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5a48ea253b357c8e6441be01918bc57c ;

Ic9c2f173881d25f8976d723957809f51 I334836058139b9a1cba37870d575f50a (
.fgallag_sel( I367ff6b11b884e02a3065fc7fe811e15[fgallag_SEL-1:0]),
.fgallag( Ic3c81f609bf98f2ded891b55bacbd453 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I20f0ea42718bdd84caf3da4a1b32c5a1 = (I367ff6b11b884e02a3065fc7fe811e15[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic3c81f609bf98f2ded891b55bacbd453 ;

Ic9c2f173881d25f8976d723957809f51 I8de2106c56422d321688ab977b4fa94b (
.fgallag_sel( I6fab19692b512166fe9c74b5e987788d[fgallag_SEL-1:0]),
.fgallag( Ie38b3f5ad91f2c983d519c9b1200559c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I11489ad40e6ff10933319784981fe59f = (I6fab19692b512166fe9c74b5e987788d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie38b3f5ad91f2c983d519c9b1200559c ;

Ic9c2f173881d25f8976d723957809f51 I6c34047a2fd5dad74e011767d9798b23 (
.fgallag_sel( I04dd73af505f618ccdb209b3cf97ceec[fgallag_SEL-1:0]),
.fgallag( I1e5e2679a0e75104cc0be107ecadd01c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I10fe1f517735fad803f3d5d75fa3d406 = (I04dd73af505f618ccdb209b3cf97ceec[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1e5e2679a0e75104cc0be107ecadd01c ;

Ic9c2f173881d25f8976d723957809f51 Icd7fe5c0f3b70f53602597e7faa083a3 (
.fgallag_sel( If8c559905d4120488d431719c4e8ce24[fgallag_SEL-1:0]),
.fgallag( I903e174feff2be7109cdb19fa15a63ec ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifed41503f4acb3625530d3c74b5ccb52 = (If8c559905d4120488d431719c4e8ce24[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I903e174feff2be7109cdb19fa15a63ec ;

Ic9c2f173881d25f8976d723957809f51 I01f58ef489c66c43d57def8bd9d7fe64 (
.fgallag_sel( I20ed4f6f14e20ce3f0e106d1b7782fcd[fgallag_SEL-1:0]),
.fgallag( I6893d09bc4fca46b4ad33c42d1950790 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic9550361e9ae769b5095df4857041e60 = (I20ed4f6f14e20ce3f0e106d1b7782fcd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6893d09bc4fca46b4ad33c42d1950790 ;

Ic9c2f173881d25f8976d723957809f51 I8c2019e6158fd6dc644fe0bc8647d895 (
.fgallag_sel( Ib10626ffa126188c5bf1fc8399107b26[fgallag_SEL-1:0]),
.fgallag( I4ec84e063fb84d278ae90b84751b1bcc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I29cedb22eb565264529effcf107e167f = (Ib10626ffa126188c5bf1fc8399107b26[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4ec84e063fb84d278ae90b84751b1bcc ;

Ic9c2f173881d25f8976d723957809f51 I776d0f5a5c8001f5e2b57d5c54c4356d (
.fgallag_sel( I29007c52357ac7afbda39d72a5bb60af[fgallag_SEL-1:0]),
.fgallag( I33998829023b087dbfa2e568d77291b3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I229b8819c94a612ca986936c96ffa9a9 = (I29007c52357ac7afbda39d72a5bb60af[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I33998829023b087dbfa2e568d77291b3 ;

Ic9c2f173881d25f8976d723957809f51 I7ecc8bea9a08d1e90dcbe59a557f757b (
.fgallag_sel( I66d367c046611f145e607a90911cf499[fgallag_SEL-1:0]),
.fgallag( I5bc68432bc0a9ea8cd024d7fc3d3fdc8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I62c0db0621c1a71960770d14c332dc0d = (I66d367c046611f145e607a90911cf499[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5bc68432bc0a9ea8cd024d7fc3d3fdc8 ;

Ic9c2f173881d25f8976d723957809f51 I6baa0bd6664b5e59451def4a2e76f699 (
.fgallag_sel( I9c4c2556f6170a8df61d909855a846ed[fgallag_SEL-1:0]),
.fgallag( Ib84e5271ffa3584148ce87dcf2a4f2a2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id94e17f3fb5b4fe7a5fbe8e25d02ec27 = (I9c4c2556f6170a8df61d909855a846ed[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib84e5271ffa3584148ce87dcf2a4f2a2 ;

Ic9c2f173881d25f8976d723957809f51 I3860ef61824e279cf9bce7712ac534ff (
.fgallag_sel( I6fadc3e8d995bb4317bf7b4377c3c2c5[fgallag_SEL-1:0]),
.fgallag( Ib633998a5fd0df508b47ba9c2f7c390a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I10cb83fe0a939bf2784eb93ca1d7b3c5 = (I6fadc3e8d995bb4317bf7b4377c3c2c5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib633998a5fd0df508b47ba9c2f7c390a ;

Ic9c2f173881d25f8976d723957809f51 I5829b006644b9595232c977a7b7f671f (
.fgallag_sel( I99b20e911c189e0616f02376ab736e91[fgallag_SEL-1:0]),
.fgallag( Ie36cfd3519810d325d5cdc5150380fe0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8f8b2e93ca65e789d13d66ecea733894 = (I99b20e911c189e0616f02376ab736e91[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie36cfd3519810d325d5cdc5150380fe0 ;

Ic9c2f173881d25f8976d723957809f51 Ibc026eb2937785ddbc10a1798e068191 (
.fgallag_sel( I5793c12f5dbdd8245dbb202d550ca960[fgallag_SEL-1:0]),
.fgallag( I6ac3755ff9de4d43d0493891b2a5758d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2527b288272a0ee2127436252a47a6aa = (I5793c12f5dbdd8245dbb202d550ca960[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6ac3755ff9de4d43d0493891b2a5758d ;

Ic9c2f173881d25f8976d723957809f51 I2d276ef7f8e35da9d708148e584cc110 (
.fgallag_sel( Id0660e9637cad1ce1a73d37188060154[fgallag_SEL-1:0]),
.fgallag( I5f0212d2ffe8f85614891882390bbc25 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I743dd733d1c20868da7a802ea99b23bb = (Id0660e9637cad1ce1a73d37188060154[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5f0212d2ffe8f85614891882390bbc25 ;

Ic9c2f173881d25f8976d723957809f51 I8989b306578253ca1ecd8254bf9b9538 (
.fgallag_sel( If5a7af7ca023e1393526e888f4220a44[fgallag_SEL-1:0]),
.fgallag( I1e009fcbec9031954637f055cb9cfe01 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5dacf7fba8d457b393930fcc76135b39 = (If5a7af7ca023e1393526e888f4220a44[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1e009fcbec9031954637f055cb9cfe01 ;

Ic9c2f173881d25f8976d723957809f51 I9618d610b0cfa33e2a1a04e589f313d1 (
.fgallag_sel( Id043eb50634e803e53adc1168379a5d0[fgallag_SEL-1:0]),
.fgallag( Ia6caeb0fcc8e7486e4d55b72a0d499a5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic50ab0fdec011923b02c0c0d717befa5 = (Id043eb50634e803e53adc1168379a5d0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia6caeb0fcc8e7486e4d55b72a0d499a5 ;

Ic9c2f173881d25f8976d723957809f51 Icd9a35d18d152c94cb60edfa57e773b0 (
.fgallag_sel( I1f866dd0b129267550aea1a267d9c91e[fgallag_SEL-1:0]),
.fgallag( I631e31da7dccd5b9311a4fa73e6a0227 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3afc7e76861fb1fa36291ac8d5508483 = (I1f866dd0b129267550aea1a267d9c91e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I631e31da7dccd5b9311a4fa73e6a0227 ;

Ic9c2f173881d25f8976d723957809f51 Id1380e6738e0783bf9e286acf90e861d (
.fgallag_sel( I8c4da05c08210fe33139c3d3e5d75d58[fgallag_SEL-1:0]),
.fgallag( Ib152eea9af905931ab45c4f9d89fa50b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7c06d7efe631bc01f98ca137df06876e = (I8c4da05c08210fe33139c3d3e5d75d58[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib152eea9af905931ab45c4f9d89fa50b ;

Ic9c2f173881d25f8976d723957809f51 I785b4074e8532eaf78443142553d4988 (
.fgallag_sel( Ib41f7b823681fdd084b6d8436a407aa8[fgallag_SEL-1:0]),
.fgallag( I94118c50e80e5fed4294d16358d41579 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifd5f5f8f7ac4238cdb3a5fb2e86eecad = (Ib41f7b823681fdd084b6d8436a407aa8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I94118c50e80e5fed4294d16358d41579 ;

Ic9c2f173881d25f8976d723957809f51 Ie0de093dc3cc1d194c2e0e7ff19bd5b2 (
.fgallag_sel( Ic5b50a785b7acac7e3be4095aa92e50a[fgallag_SEL-1:0]),
.fgallag( I1269d97f8ab4f5dddc002acf38b4a189 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I17e9d58c80d0da6e6093836deecfa743 = (Ic5b50a785b7acac7e3be4095aa92e50a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1269d97f8ab4f5dddc002acf38b4a189 ;

Ic9c2f173881d25f8976d723957809f51 If9c3f5b87787afc8e25e225e35c591a9 (
.fgallag_sel( I3ffbe03796b66d00d47fd918be60ab89[fgallag_SEL-1:0]),
.fgallag( I89a793ddaf4887ddb8dbaaba13225d08 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icd18edbcc227111c037023bf2b57ee5a = (I3ffbe03796b66d00d47fd918be60ab89[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I89a793ddaf4887ddb8dbaaba13225d08 ;

Ic9c2f173881d25f8976d723957809f51 I035a19d490c19fbb1eaaa6673fb01a58 (
.fgallag_sel( Ifc92a916da938ef6164db250be635f88[fgallag_SEL-1:0]),
.fgallag( I2b4fe952791866aecbbbcf01257d527b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id22f8eb74ec1e8499e150278e438359d = (Ifc92a916da938ef6164db250be635f88[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2b4fe952791866aecbbbcf01257d527b ;

Ic9c2f173881d25f8976d723957809f51 I0a2ee30a89a2254461e1b7679a4490fa (
.fgallag_sel( I8ccd42508ce7d5bd897c2cf0c54caeb3[fgallag_SEL-1:0]),
.fgallag( I797321bb9e3c2d7d3727af9a4cf5418b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id10ed140128d500e98d984a15b479fb4 = (I8ccd42508ce7d5bd897c2cf0c54caeb3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I797321bb9e3c2d7d3727af9a4cf5418b ;

Ic9c2f173881d25f8976d723957809f51 Ib700045c49f1212c46ffed81f1787daf (
.fgallag_sel( I4920e7e82749cc036b58a7cd0a03e327[fgallag_SEL-1:0]),
.fgallag( I5eeb78b1511aa7b76765d82328323a4c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If89f8e436166d9beeca9937c45b2c7d5 = (I4920e7e82749cc036b58a7cd0a03e327[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5eeb78b1511aa7b76765d82328323a4c ;

Ic9c2f173881d25f8976d723957809f51 I7527ff564b5a3c4be2ba599acfedccdd (
.fgallag_sel( Ie1040b2aa91f272e4449c4b5f9f8f575[fgallag_SEL-1:0]),
.fgallag( I55f8232fcfcb929a35717f724f44eb4c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idfd24573e271b5cdd6f051496cb6ba8f = (Ie1040b2aa91f272e4449c4b5f9f8f575[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I55f8232fcfcb929a35717f724f44eb4c ;

Ic9c2f173881d25f8976d723957809f51 I01fb6c8bfe9eaa892e9fd0e89a5bae28 (
.fgallag_sel( I65968fb0f63d52ad96cd8fa270126a1b[fgallag_SEL-1:0]),
.fgallag( I7a7705607e93fca1cf1e7b1c92c4e3cc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I145c31d89636b936f18a19bf50966bbe = (I65968fb0f63d52ad96cd8fa270126a1b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7a7705607e93fca1cf1e7b1c92c4e3cc ;

Ic9c2f173881d25f8976d723957809f51 I8f71a60b9546637d6f947757d3015b4b (
.fgallag_sel( I839ac8ee59f51d4c3de92ba5cb26e788[fgallag_SEL-1:0]),
.fgallag( I7e2e0ffb2b5622ba6e03a47755a9a1dc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I15cae93770d041e2ef681a81e8256059 = (I839ac8ee59f51d4c3de92ba5cb26e788[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7e2e0ffb2b5622ba6e03a47755a9a1dc ;

Ic9c2f173881d25f8976d723957809f51 I5debfc999dfca9187b236439b51947cf (
.fgallag_sel( I33cd95f1919318a0f3df5df7310d64c6[fgallag_SEL-1:0]),
.fgallag( I5f50e835526833015a2087dbdb77686e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6a86457e1b16bfc515084fe599281818 = (I33cd95f1919318a0f3df5df7310d64c6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5f50e835526833015a2087dbdb77686e ;

Ic9c2f173881d25f8976d723957809f51 I02f3bb6429030161631cd0286e61f838 (
.fgallag_sel( I4933e8d16fba26cd797b25a9ac2a2de8[fgallag_SEL-1:0]),
.fgallag( I98f32439ec64d796ebb157815b259aa2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2453c39e5805313c3a8fd0d074058916 = (I4933e8d16fba26cd797b25a9ac2a2de8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I98f32439ec64d796ebb157815b259aa2 ;

Ic9c2f173881d25f8976d723957809f51 I103ecc8bd400c9590ee9df342a34629d (
.fgallag_sel( I218f7578eb748e31d0002052f30c5842[fgallag_SEL-1:0]),
.fgallag( Id59ca1b1cff93a8544c54c6d4ee22b2f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I34636cc42b16776295078bd349a76ac6 = (I218f7578eb748e31d0002052f30c5842[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id59ca1b1cff93a8544c54c6d4ee22b2f ;

Ic9c2f173881d25f8976d723957809f51 I046bae774c128788dfcad9a0a5f9c812 (
.fgallag_sel( I2a808d1c42ad758ae3baaaee8129dfb2[fgallag_SEL-1:0]),
.fgallag( I726538434626c5202d53d29faedddd56 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I48f8d5589f772fbb4b3923fbd213e7f7 = (I2a808d1c42ad758ae3baaaee8129dfb2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I726538434626c5202d53d29faedddd56 ;

Ic9c2f173881d25f8976d723957809f51 I5d0280a20c165388e6a95d083ff7d754 (
.fgallag_sel( I4e851fd3c114af87f5e8c68c02594e3a[fgallag_SEL-1:0]),
.fgallag( I8ea236c734f7b96620a37750134d3872 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I83e4b71b0a0a3a82fc0a9fb56f803fa9 = (I4e851fd3c114af87f5e8c68c02594e3a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8ea236c734f7b96620a37750134d3872 ;

Ic9c2f173881d25f8976d723957809f51 I22fa2882526275e8b20d4d7289285a3c (
.fgallag_sel( I0da40f88adc46e90f616acdcdb8e0e2c[fgallag_SEL-1:0]),
.fgallag( I259d7244226dbcbd1d02df5ca164afdc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2abd0942d4d5e3aff2d24db9656c025f = (I0da40f88adc46e90f616acdcdb8e0e2c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I259d7244226dbcbd1d02df5ca164afdc ;

Ic9c2f173881d25f8976d723957809f51 Idf82769f4d0db7093e82d42f13c4b3ca (
.fgallag_sel( I0dee7767e472a5fd71250ae6c57cc8b5[fgallag_SEL-1:0]),
.fgallag( I086375f289b769938edfc8b9b5146714 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0fa19f52fef5a583890e3096eb23f1db = (I0dee7767e472a5fd71250ae6c57cc8b5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I086375f289b769938edfc8b9b5146714 ;

Ic9c2f173881d25f8976d723957809f51 I86d5b425f6a3f5fbcfd5148b7fbdc478 (
.fgallag_sel( I9f40be7552b3dd625e5bce0befc5a548[fgallag_SEL-1:0]),
.fgallag( Icb82f8092f14511d62f7cbe821af9faf ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0e4a9bf26a9df3551a69edced6128e30 = (I9f40be7552b3dd625e5bce0befc5a548[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Icb82f8092f14511d62f7cbe821af9faf ;

Ic9c2f173881d25f8976d723957809f51 Icc597684dd6471072d87ef841d2f48be (
.fgallag_sel( I8fdf98ffd757c8845ed6ffa4ddd1a16b[fgallag_SEL-1:0]),
.fgallag( I7e8df00362c29bd3924ecbe3dd1db23c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icd359ef9d3a983f4258cc4441110cc97 = (I8fdf98ffd757c8845ed6ffa4ddd1a16b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7e8df00362c29bd3924ecbe3dd1db23c ;

Ic9c2f173881d25f8976d723957809f51 I4014408b9ff9d90c7323cc66ea362b40 (
.fgallag_sel( I8103b777314a4fa471e0898fde9cde08[fgallag_SEL-1:0]),
.fgallag( If1014cbbd6e267aaacbcf3c8ba33a98b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I31d6000373f248b1dde9fc0108bfd280 = (I8103b777314a4fa471e0898fde9cde08[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If1014cbbd6e267aaacbcf3c8ba33a98b ;

Ic9c2f173881d25f8976d723957809f51 I6322eba8be2a8a3d10083745d6bf0e88 (
.fgallag_sel( If6c3ee8e0d7dea58043d5be0f4630873[fgallag_SEL-1:0]),
.fgallag( Iae4dfe3ede67923e8b740dd575b216b6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I445cd3125f69b7e29d582a4803709c8f = (If6c3ee8e0d7dea58043d5be0f4630873[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iae4dfe3ede67923e8b740dd575b216b6 ;

Ic9c2f173881d25f8976d723957809f51 I62906715977232c418942cdd1799aa92 (
.fgallag_sel( I711a5171f591f472cdbfc9a0f5e1aa17[fgallag_SEL-1:0]),
.fgallag( Iccfddf46ea48242ca751b5d53f98d270 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2a8dcc8d3db0d8b5bb54bc7fae5e6ca7 = (I711a5171f591f472cdbfc9a0f5e1aa17[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iccfddf46ea48242ca751b5d53f98d270 ;

Ic9c2f173881d25f8976d723957809f51 I946e9fec0507e526fdd99cdac1e033de (
.fgallag_sel( Ic30bc38184dfbbd694af52640692709d[fgallag_SEL-1:0]),
.fgallag( I804705ac9a613b4107c8ceaac4127386 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibbf4549a33d4916489e7e325a811add1 = (Ic30bc38184dfbbd694af52640692709d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I804705ac9a613b4107c8ceaac4127386 ;

Ic9c2f173881d25f8976d723957809f51 I77c1c299bea377ba2ae6e113969f786a (
.fgallag_sel( I422f6fd1d273a3834d04b04ab8e2812d[fgallag_SEL-1:0]),
.fgallag( I8f40972503fbfdab92676a32f351dfe6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9a2d80bf2bbc2101c8e426cfc1c8277b = (I422f6fd1d273a3834d04b04ab8e2812d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8f40972503fbfdab92676a32f351dfe6 ;

Ic9c2f173881d25f8976d723957809f51 I27c934da26f862be210aad00f7ec7eb6 (
.fgallag_sel( Ia0fdc60b90ad18b6585ec1ad4e89e80b[fgallag_SEL-1:0]),
.fgallag( I8fc9ec077c7c6ce5e2660a4530a234ae ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I71c9904d29e88f0a5e6d7f8ec88de592 = (Ia0fdc60b90ad18b6585ec1ad4e89e80b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8fc9ec077c7c6ce5e2660a4530a234ae ;

Ic9c2f173881d25f8976d723957809f51 I2b258bde38b47625ccd6f4e5fee0b610 (
.fgallag_sel( I7809fe7a30d041a7e569ffe890242df8[fgallag_SEL-1:0]),
.fgallag( I3e3bf3c2155f584784863ae41cb73c7d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic6c8869890916818213809df90b52856 = (I7809fe7a30d041a7e569ffe890242df8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3e3bf3c2155f584784863ae41cb73c7d ;

Ic9c2f173881d25f8976d723957809f51 I2ac45958d5493d6b92ec6fac9e7a96fb (
.fgallag_sel( I672b14ec1b3c4797545f266727505a85[fgallag_SEL-1:0]),
.fgallag( I9cc24d95a0ddbe4145d144003778eebc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3c61b092287e1f2c446aa7346b3dfcfb = (I672b14ec1b3c4797545f266727505a85[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9cc24d95a0ddbe4145d144003778eebc ;

Ic9c2f173881d25f8976d723957809f51 I1b062f157cee8fe91e61dd48c5dc2b8d (
.fgallag_sel( If9620d20ebaae6245a2c386d9bf5fdb1[fgallag_SEL-1:0]),
.fgallag( Ib9b96de1e217660c2ac9f7815249c6a2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8f94e1fe9df14c5dd75421cdfe8b1efe = (If9620d20ebaae6245a2c386d9bf5fdb1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib9b96de1e217660c2ac9f7815249c6a2 ;

Ic9c2f173881d25f8976d723957809f51 Idb90b29bee5f73787888e40b65292d5a (
.fgallag_sel( Ic74e22bffd88f32eefe499cde0fafa8a[fgallag_SEL-1:0]),
.fgallag( I2cc498e11d3d487d1e8319df8521ff6d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie2a432bd8429925297936c8aebf7282f = (Ic74e22bffd88f32eefe499cde0fafa8a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2cc498e11d3d487d1e8319df8521ff6d ;

Ic9c2f173881d25f8976d723957809f51 I5ca084a426c39605ae76b7fee1d434fb (
.fgallag_sel( I76d38ce67387bd76ab45c9cba7d18b31[fgallag_SEL-1:0]),
.fgallag( Iae3d8158d13c8179719cbe12fdd7f9ab ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I309c99cc023e0c7804b2574821d63f10 = (I76d38ce67387bd76ab45c9cba7d18b31[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iae3d8158d13c8179719cbe12fdd7f9ab ;

Ic9c2f173881d25f8976d723957809f51 I921198366330c15b64ed56a0667ed038 (
.fgallag_sel( I44413c6f6f6493f8a86abf6eb32604f6[fgallag_SEL-1:0]),
.fgallag( Ieadf1b0e427ecddd261297ae4054a0bd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5806c65240e9ce9f9d0804d063c2674e = (I44413c6f6f6493f8a86abf6eb32604f6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ieadf1b0e427ecddd261297ae4054a0bd ;

Ic9c2f173881d25f8976d723957809f51 Id6303dc54850b16c0b6d5b8832e2c411 (
.fgallag_sel( I67f632fca617fe06565ddcaaee8fa8b8[fgallag_SEL-1:0]),
.fgallag( I8dbe4e03db655e1f691254835fb58798 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib73d05919f3373f122b121be5a038f4b = (I67f632fca617fe06565ddcaaee8fa8b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8dbe4e03db655e1f691254835fb58798 ;

Ic9c2f173881d25f8976d723957809f51 I674f492f5570a8650f53521ceb348141 (
.fgallag_sel( I3fd38a71ce6aa3db1d7a5a9f8a991e12[fgallag_SEL-1:0]),
.fgallag( I14b22818be28bc385f91920399012555 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I84136dfec9c8ab98228801deffbe8c19 = (I3fd38a71ce6aa3db1d7a5a9f8a991e12[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I14b22818be28bc385f91920399012555 ;

Ic9c2f173881d25f8976d723957809f51 Ibd0522c32e0095fdd4e4b00327da3023 (
.fgallag_sel( I63e5718bf7d8771ef90b91be73d73264[fgallag_SEL-1:0]),
.fgallag( Id2878a17128a23eee2272c7e39743bd3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I09e9850f90a7f073169e66c9e2339f51 = (I63e5718bf7d8771ef90b91be73d73264[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id2878a17128a23eee2272c7e39743bd3 ;

Ic9c2f173881d25f8976d723957809f51 I0cb97ba4591f86695e53b3e4dcd071bd (
.fgallag_sel( Ie385e1aeb2b0dcf6d2454be3d7708b27[fgallag_SEL-1:0]),
.fgallag( I3701d2d2e74c43b3ae347902c0efff20 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1260922a3e6cd464e43f215299d70ef1 = (Ie385e1aeb2b0dcf6d2454be3d7708b27[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3701d2d2e74c43b3ae347902c0efff20 ;

Ic9c2f173881d25f8976d723957809f51 I25e7839c15678fbceba9348701eb0f3b (
.fgallag_sel( Ib2d1b7e105b25b492b45da72536d7578[fgallag_SEL-1:0]),
.fgallag( Id6487b559b7ebad725aa43382f09bab3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I97cf4612b19722d7f5f4cf9a867a9b22 = (Ib2d1b7e105b25b492b45da72536d7578[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id6487b559b7ebad725aa43382f09bab3 ;

Ic9c2f173881d25f8976d723957809f51 I16774b96670d829cfe7720bd7f3e821e (
.fgallag_sel( I588abf5ef4c583f0fec422736a0ce6a0[fgallag_SEL-1:0]),
.fgallag( Ib6ea830665d44628aef5041b2fa46328 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4856ddf90e056e12eb6ec14d66f776b3 = (I588abf5ef4c583f0fec422736a0ce6a0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib6ea830665d44628aef5041b2fa46328 ;

Ic9c2f173881d25f8976d723957809f51 I3a13ded4b9783619a18e4a1b0f339601 (
.fgallag_sel( I58bb95c56c7be17c263a2161210d7d8d[fgallag_SEL-1:0]),
.fgallag( Ia6181e1acc2ea46a85626a22983e2662 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I370986beb4c411ce7154bb1c7045c5d8 = (I58bb95c56c7be17c263a2161210d7d8d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia6181e1acc2ea46a85626a22983e2662 ;

Ic9c2f173881d25f8976d723957809f51 If7530f5b730ac2d11cfdd58c941e52a5 (
.fgallag_sel( Ifaf0e1f21b3bd7393c475b5126540a72[fgallag_SEL-1:0]),
.fgallag( I8b38fb1f95f036393933d07e0a60b875 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0b22c5487df5e2b47d2ac3e16ca195b9 = (Ifaf0e1f21b3bd7393c475b5126540a72[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8b38fb1f95f036393933d07e0a60b875 ;

Ic9c2f173881d25f8976d723957809f51 I16a31de65046934872600db782c63bbb (
.fgallag_sel( I7027db9e0450724a6d417d708f1043f2[fgallag_SEL-1:0]),
.fgallag( I33d76ad1185bbf80de5e8ff0ad52b15f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic7437fa32ca344b6eaa895d35d335e57 = (I7027db9e0450724a6d417d708f1043f2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I33d76ad1185bbf80de5e8ff0ad52b15f ;

Ic9c2f173881d25f8976d723957809f51 Ib0f31439087a976b322adcd6c2946f27 (
.fgallag_sel( Iebcb7206d8860b5094459c5d10b4efed[fgallag_SEL-1:0]),
.fgallag( If2c522a90684b77b18f0058d1d2b14d8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1dcfffaaabc223ae08cd9d08d6e968d2 = (Iebcb7206d8860b5094459c5d10b4efed[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If2c522a90684b77b18f0058d1d2b14d8 ;

Ic9c2f173881d25f8976d723957809f51 I67a4b9edd8a15693944d7ecf83504396 (
.fgallag_sel( I6bbf2b47a7dc50e66a3d8d258d6e31fb[fgallag_SEL-1:0]),
.fgallag( I869e040de179572cdfd9373a4de8b31c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I16bb10e8ddda86c2c8a1df7b0ec4c133 = (I6bbf2b47a7dc50e66a3d8d258d6e31fb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I869e040de179572cdfd9373a4de8b31c ;

Ic9c2f173881d25f8976d723957809f51 I183de27fe84e629fbf41ce15613a6fff (
.fgallag_sel( I8459abaa907f5afcd11884b1ec8c06c5[fgallag_SEL-1:0]),
.fgallag( I3fb8890ee1f1cb30ecdf50d69e4ac0fa ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I50ab3193dde101b550b508744be5a775 = (I8459abaa907f5afcd11884b1ec8c06c5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3fb8890ee1f1cb30ecdf50d69e4ac0fa ;

Ic9c2f173881d25f8976d723957809f51 Ie125844167090094359a499e4ff84205 (
.fgallag_sel( Ia16ae2f6ef5000d47b6b84ed058252aa[fgallag_SEL-1:0]),
.fgallag( I6b60e2478c009889776de20209929ee0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I022ed4e5e55e9c3cd418bca5475beb82 = (Ia16ae2f6ef5000d47b6b84ed058252aa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6b60e2478c009889776de20209929ee0 ;

Ic9c2f173881d25f8976d723957809f51 Ifd0a5a99f85260cf3da5d23e8defd5af (
.fgallag_sel( Ica32690dbc9ea110fefdce92260b125c[fgallag_SEL-1:0]),
.fgallag( Ie6b559c2f0bd388d072b660341eebe31 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie44afe129f71022f34e9f9cb5ac4eb3d = (Ica32690dbc9ea110fefdce92260b125c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie6b559c2f0bd388d072b660341eebe31 ;

Ic9c2f173881d25f8976d723957809f51 Ie60decf00039f8d036a69d931da76641 (
.fgallag_sel( Ic431d9383cce30b1889c92e2be4cb9d0[fgallag_SEL-1:0]),
.fgallag( Ia46aa3a3e6a01d4690dfe0e7f1eab548 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I38c8f2c90a4d997e5597b462e7e8c613 = (Ic431d9383cce30b1889c92e2be4cb9d0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia46aa3a3e6a01d4690dfe0e7f1eab548 ;

Ic9c2f173881d25f8976d723957809f51 Ia1d603b65db534d8f996f302b15df27a (
.fgallag_sel( Ib9cca4c0e58373c26d5fd9f51f793898[fgallag_SEL-1:0]),
.fgallag( Idb7244908662bcd97fe8fe0db4b1abdc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib38a5e546fdc5837a97c4ff3a627777d = (Ib9cca4c0e58373c26d5fd9f51f793898[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idb7244908662bcd97fe8fe0db4b1abdc ;

Ic9c2f173881d25f8976d723957809f51 I3996ab9886309f0f84f9b6c29ddd804e (
.fgallag_sel( I99bf0bc8ac20832b3724b2753f6ca449[fgallag_SEL-1:0]),
.fgallag( If570b3495ea5b3f250cf4873f5dd0bb9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iaebf3465f121a3c054c87227d7e9e167 = (I99bf0bc8ac20832b3724b2753f6ca449[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If570b3495ea5b3f250cf4873f5dd0bb9 ;

Ic9c2f173881d25f8976d723957809f51 I87909992668f40e30f720eb45760724d (
.fgallag_sel( Ie701008f3c60c51ed72c5f964a8fc36e[fgallag_SEL-1:0]),
.fgallag( I50bbcccc40af5e9700b97e682953c8c9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6fd1108c6ac90f5c69db5aca76055a32 = (Ie701008f3c60c51ed72c5f964a8fc36e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I50bbcccc40af5e9700b97e682953c8c9 ;

Ic9c2f173881d25f8976d723957809f51 I1c31cdc3d8551f893a8391bbb8ca1612 (
.fgallag_sel( I3e2d78f8307a1787f8b2eccba94c7557[fgallag_SEL-1:0]),
.fgallag( I5422f11a7e0b646dd4fa254602f91b34 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If6f92d3b43974c88963a188a26bc3009 = (I3e2d78f8307a1787f8b2eccba94c7557[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5422f11a7e0b646dd4fa254602f91b34 ;

Ic9c2f173881d25f8976d723957809f51 I1a13684b6014ae4d686a25a7dd3df995 (
.fgallag_sel( Ic1b4444ab0df9745d29bf893d9b83168[fgallag_SEL-1:0]),
.fgallag( Ic5c34f86b03fffdcf723ff4116822e3f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I19fb6cacc6841dec5653ef273676f18f = (Ic1b4444ab0df9745d29bf893d9b83168[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic5c34f86b03fffdcf723ff4116822e3f ;

Ic9c2f173881d25f8976d723957809f51 I39d6ac57ceb46bbf9013a67ae84d3f93 (
.fgallag_sel( I5f52dbf600656a8f5dc6b6b8a45ccebe[fgallag_SEL-1:0]),
.fgallag( I2ebd72fb063702a7c36b4b546f4b94b8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia0abbf270f98b4bf4f29b56611db23b6 = (I5f52dbf600656a8f5dc6b6b8a45ccebe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2ebd72fb063702a7c36b4b546f4b94b8 ;

Ic9c2f173881d25f8976d723957809f51 I91acc92a6e9c029331b75b3d30385864 (
.fgallag_sel( I7f307af79f45ad4b9511e3961c917078[fgallag_SEL-1:0]),
.fgallag( I6328eca7325eea20ccf30adf8b928edb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I38ad3c494c777f3985d61eef7cab8fb6 = (I7f307af79f45ad4b9511e3961c917078[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6328eca7325eea20ccf30adf8b928edb ;

Ic9c2f173881d25f8976d723957809f51 Ide58f30cc36825833f3a0e2b9113fd3c (
.fgallag_sel( Ie17a5be2a16d2efb98c976d7ee882535[fgallag_SEL-1:0]),
.fgallag( Ica13fd6daec896ddb0fa6be797edf6bb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ieb8d87fc8ecfad97cb9840b3739d6ea4 = (Ie17a5be2a16d2efb98c976d7ee882535[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ica13fd6daec896ddb0fa6be797edf6bb ;

Ic9c2f173881d25f8976d723957809f51 I3f894a76006a293eae83dde7699a69f7 (
.fgallag_sel( I5f19d2adff2f34a4bebe03f929a09c49[fgallag_SEL-1:0]),
.fgallag( I970c832cf68b5178f3d8111c9fed3b5a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic1087bae156ef4dd5fe218537432b0ed = (I5f19d2adff2f34a4bebe03f929a09c49[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I970c832cf68b5178f3d8111c9fed3b5a ;

Ic9c2f173881d25f8976d723957809f51 I7ac46b6d57f07f4c5f0b00c34819501c (
.fgallag_sel( I3cd69aeed9e869a2096d6dced5c209a0[fgallag_SEL-1:0]),
.fgallag( I65f78ccc122f96f97fee54955d370288 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6655118cfe24b706e6557438ffa1711a = (I3cd69aeed9e869a2096d6dced5c209a0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I65f78ccc122f96f97fee54955d370288 ;

Ic9c2f173881d25f8976d723957809f51 I5bc071af22c22c2283ef60a34fbd6f6f (
.fgallag_sel( I359b6a22c9568a13b81670c741281393[fgallag_SEL-1:0]),
.fgallag( I5f77d7804a3e4adb641908be74f3ea19 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia12b8e62d6e1d52861589818deb6a851 = (I359b6a22c9568a13b81670c741281393[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5f77d7804a3e4adb641908be74f3ea19 ;

Ic9c2f173881d25f8976d723957809f51 I72a88a5d0350eb125ad88ca4861bea27 (
.fgallag_sel( I24ba99614df383c38bbac50ae8b4487e[fgallag_SEL-1:0]),
.fgallag( I9263e4ab78ca05f93ff921c4fd9ff787 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I59260857d96064096680b8361521b588 = (I24ba99614df383c38bbac50ae8b4487e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9263e4ab78ca05f93ff921c4fd9ff787 ;

Ic9c2f173881d25f8976d723957809f51 I8bbb846a8d8b0b5348d52c915b2fc3bf (
.fgallag_sel( I7498bee46de6b1c946ce95fdcc89f6e5[fgallag_SEL-1:0]),
.fgallag( I6f8f253cfb1fe1c2254e557f732a9b22 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iee39a5d6276b276729abd14472262ed1 = (I7498bee46de6b1c946ce95fdcc89f6e5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6f8f253cfb1fe1c2254e557f732a9b22 ;

Ic9c2f173881d25f8976d723957809f51 Ie3a715f0fd86beedb2b36e6dbe22f0d2 (
.fgallag_sel( I0f644f42cabf871b71e5a82871bc7b5d[fgallag_SEL-1:0]),
.fgallag( I3f247e74edd47e346d3bbb5dc3408844 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I20aa2879f47abd3c368f7494d944222d = (I0f644f42cabf871b71e5a82871bc7b5d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3f247e74edd47e346d3bbb5dc3408844 ;

Ic9c2f173881d25f8976d723957809f51 I5224853b7e9d431d0eaa6076dd492253 (
.fgallag_sel( I71f9e059726a6cac8bdf0efcc0eadd2b[fgallag_SEL-1:0]),
.fgallag( Ie0b33e2c1def11ccdaaae4ed2b042df6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If0192b9580e5fdb8d71b422ccb28666f = (I71f9e059726a6cac8bdf0efcc0eadd2b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie0b33e2c1def11ccdaaae4ed2b042df6 ;

Ic9c2f173881d25f8976d723957809f51 I336d4422917abebf910f1e4e298844f9 (
.fgallag_sel( I0c9b2c1da30bfab514bbb556ae7bd4c4[fgallag_SEL-1:0]),
.fgallag( I39448514454c92ce93c3b0bc1d0e5d50 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5095a3f4dd1c3bca218d17f5c609b667 = (I0c9b2c1da30bfab514bbb556ae7bd4c4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I39448514454c92ce93c3b0bc1d0e5d50 ;

Ic9c2f173881d25f8976d723957809f51 I051db3a777b48cd31280a285a2fd1d04 (
.fgallag_sel( I7918b2e37e96aee94fbccca7e0f75fc4[fgallag_SEL-1:0]),
.fgallag( I677e9047c3ede581db9512b4fe072ea9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iea2a2368935757fe57b3d283fdccdb3e = (I7918b2e37e96aee94fbccca7e0f75fc4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I677e9047c3ede581db9512b4fe072ea9 ;

Ic9c2f173881d25f8976d723957809f51 I73937b440876c63c6c0e4651c18b1d13 (
.fgallag_sel( I76eebd77eb77e0abcbc727d2c511370a[fgallag_SEL-1:0]),
.fgallag( Ief6fbe6927f26b7a037f8e0bcb7751d8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I36cd8882960099f242551ff3cbf8e4bd = (I76eebd77eb77e0abcbc727d2c511370a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ief6fbe6927f26b7a037f8e0bcb7751d8 ;

Ic9c2f173881d25f8976d723957809f51 Ia96d424c061446fdb4bca919359b11d4 (
.fgallag_sel( Ibb2288e62110bae5b2d3fe901974e5c7[fgallag_SEL-1:0]),
.fgallag( Ie1e5c12afad8f2d8c2abef26473b7d9c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3ac47b1ac8e31b0082c7acfab65e222c = (Ibb2288e62110bae5b2d3fe901974e5c7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie1e5c12afad8f2d8c2abef26473b7d9c ;

Ic9c2f173881d25f8976d723957809f51 I08f59b74433f85cb5aaa33f996dcd038 (
.fgallag_sel( I080f931dfef9d8adfb1dc1ee073eb64c[fgallag_SEL-1:0]),
.fgallag( Ic8f2ae80147ee27c548de195dfefa382 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2a4914c71690073767e6f5fe13f26178 = (I080f931dfef9d8adfb1dc1ee073eb64c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic8f2ae80147ee27c548de195dfefa382 ;

Ic9c2f173881d25f8976d723957809f51 Ia3505842f370f07297eb60ad7f4c87c8 (
.fgallag_sel( Ide1106431e3565158bd81ccd6b18f3a1[fgallag_SEL-1:0]),
.fgallag( I533eb0729cc85339e2fcd1847930adc9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I99903b3dad6af712c1148c2f43194da0 = (Ide1106431e3565158bd81ccd6b18f3a1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I533eb0729cc85339e2fcd1847930adc9 ;

Ic9c2f173881d25f8976d723957809f51 I4f88744cf95346d7e5304ade8d31c4de (
.fgallag_sel( I63df19931e8d28666cccd79922cbd418[fgallag_SEL-1:0]),
.fgallag( Ic68fd0a9ea4b641913aadb7fe011d8ab ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icccc370bf2f48ce93f479d13fa7075e9 = (I63df19931e8d28666cccd79922cbd418[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic68fd0a9ea4b641913aadb7fe011d8ab ;

Ic9c2f173881d25f8976d723957809f51 Iec535cb175233622735018e39dd64ec0 (
.fgallag_sel( I9a7e4a59447048de90446f877eb06627[fgallag_SEL-1:0]),
.fgallag( Ica1f13759a67176573842e56bcdf09bd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5b5a0ccc2f5f9a7554d6d55b0dc61d76 = (I9a7e4a59447048de90446f877eb06627[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ica1f13759a67176573842e56bcdf09bd ;

Ic9c2f173881d25f8976d723957809f51 I15091ee4cdbc4c1f9eb3b034e56f9194 (
.fgallag_sel( I0917e92ed84363ca92fd2074acd74eba[fgallag_SEL-1:0]),
.fgallag( Ifed30886099cbeb5da64d1d0696bb5de ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0cd3d6b7cb85a87bfbebc1982c5fddf7 = (I0917e92ed84363ca92fd2074acd74eba[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifed30886099cbeb5da64d1d0696bb5de ;

Ic9c2f173881d25f8976d723957809f51 I6d1278a14ade7356523bfb25e20f628f (
.fgallag_sel( Ie3eefdf7b5561a90a6ddd9e6aa432509[fgallag_SEL-1:0]),
.fgallag( I317b34a0f6e16550b4a3e887cdd0c250 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I38a9b558c3289d954fe0de802b473be4 = (Ie3eefdf7b5561a90a6ddd9e6aa432509[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I317b34a0f6e16550b4a3e887cdd0c250 ;

Ic9c2f173881d25f8976d723957809f51 I6e49777493eed9b55477815e7d00be9d (
.fgallag_sel( I56eeb10d11e886cff629457a640a1c76[fgallag_SEL-1:0]),
.fgallag( I39fa2bacef89a2f523f91b1e7f3cbe90 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iacadd2fc2b7446edd7c45341a0670cb7 = (I56eeb10d11e886cff629457a640a1c76[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I39fa2bacef89a2f523f91b1e7f3cbe90 ;

Ic9c2f173881d25f8976d723957809f51 I0be8508e992282e94d48eb707a43ed89 (
.fgallag_sel( I7a9eea89c4e76d856df44b6bdc332840[fgallag_SEL-1:0]),
.fgallag( Id01272140c18ae29a8c75e493cf01268 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I316810ae743e5626556ad8f3176849bc = (I7a9eea89c4e76d856df44b6bdc332840[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id01272140c18ae29a8c75e493cf01268 ;

Ic9c2f173881d25f8976d723957809f51 Iaef181cab0b8c58fef92ff35c455c444 (
.fgallag_sel( If8d8f4333e893788fcb9ec54256e5b7a[fgallag_SEL-1:0]),
.fgallag( I4d981fbbadbaa97ef98429ac12ca6710 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib9d5224a4d0b87aeb65cd6cf030ee52e = (If8d8f4333e893788fcb9ec54256e5b7a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4d981fbbadbaa97ef98429ac12ca6710 ;

Ic9c2f173881d25f8976d723957809f51 Ib09322f890f417bfa739971d0b40040a (
.fgallag_sel( Ie4af0e7e04778d85f5dee73da33376a8[fgallag_SEL-1:0]),
.fgallag( I2a1672224d3a3c513f2f04bb4dc123e0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I92246b941db36e725ce7cbb1c9b4a0b5 = (Ie4af0e7e04778d85f5dee73da33376a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2a1672224d3a3c513f2f04bb4dc123e0 ;

Ic9c2f173881d25f8976d723957809f51 I9065816af419fcb1b35fab2fe9221d0d (
.fgallag_sel( I019a4e997adf54f5f5ca651f80b7901b[fgallag_SEL-1:0]),
.fgallag( I364afb3546858e133a2bb541798e7886 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I62b8229b8e21a4bfd043c23450ff50e5 = (I019a4e997adf54f5f5ca651f80b7901b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I364afb3546858e133a2bb541798e7886 ;

Ic9c2f173881d25f8976d723957809f51 I44ac6b42b40b59272875bad6f519921e (
.fgallag_sel( I10294667f09abbfd4e2f757c414072fc[fgallag_SEL-1:0]),
.fgallag( I9908671d65856b8714d43d83f0811a17 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I49266ae645036370bba4d99a1a85bc6f = (I10294667f09abbfd4e2f757c414072fc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9908671d65856b8714d43d83f0811a17 ;

Ic9c2f173881d25f8976d723957809f51 If3994abeefefff274c4ef13f079134bb (
.fgallag_sel( Id4e8ab8f15b36bd27d1e4ebc5cbe1495[fgallag_SEL-1:0]),
.fgallag( I3e3f06cade9b6c8ea10e45996449e405 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I242c35248366a124753da854841595a7 = (Id4e8ab8f15b36bd27d1e4ebc5cbe1495[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3e3f06cade9b6c8ea10e45996449e405 ;

Ic9c2f173881d25f8976d723957809f51 I3c72cc8cb0b0973962c1a4e817d6a2c0 (
.fgallag_sel( I6c93588ca9e7c623d75314da39e89a91[fgallag_SEL-1:0]),
.fgallag( I9525b42d4dc80c42608cfa0ea10b8b2d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I347dd57356eb6e025dada067d0f661b9 = (I6c93588ca9e7c623d75314da39e89a91[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9525b42d4dc80c42608cfa0ea10b8b2d ;

Ic9c2f173881d25f8976d723957809f51 Iabbbe8e3f8d6deb5c142a17d6c5587ad (
.fgallag_sel( I1020412efc78d12a9ebcbaeb83e5dcea[fgallag_SEL-1:0]),
.fgallag( I94361c7eb9f16c4b20dfcdb7b8ad8cf3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6bb3031e93da171fac995de3e23c8b71 = (I1020412efc78d12a9ebcbaeb83e5dcea[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I94361c7eb9f16c4b20dfcdb7b8ad8cf3 ;

Ic9c2f173881d25f8976d723957809f51 Ibf6f5867a95bf2289280401e3641058c (
.fgallag_sel( Id0b574f35a83dcfd4481a10043cd1884[fgallag_SEL-1:0]),
.fgallag( Idc043493a919ec50417594df96f4d669 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I88cede4b89eb0f3917530d0ce2468c3a = (Id0b574f35a83dcfd4481a10043cd1884[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idc043493a919ec50417594df96f4d669 ;

Ic9c2f173881d25f8976d723957809f51 Ia06321b5ea2f80034cbe4fbf224367c9 (
.fgallag_sel( Ifc577e5c2c7288373a8c5e3969ac1589[fgallag_SEL-1:0]),
.fgallag( I9e051ecfe79c36a913b15a0c7fe27f4d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3a590077bea5f1023ac006b321083554 = (Ifc577e5c2c7288373a8c5e3969ac1589[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9e051ecfe79c36a913b15a0c7fe27f4d ;

Ic9c2f173881d25f8976d723957809f51 Ia308b6206fdcfb6bd85ce805d5775d46 (
.fgallag_sel( Id18a1a17c1cf6e8a2492aa73b62898f2[fgallag_SEL-1:0]),
.fgallag( I5479857f4f724aaea25ba124c9edb232 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2bac571cd0d32e8a1bd527245a76f11b = (Id18a1a17c1cf6e8a2492aa73b62898f2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5479857f4f724aaea25ba124c9edb232 ;

Ic9c2f173881d25f8976d723957809f51 I9c3f5975bdbeb13129733c80b3b81416 (
.fgallag_sel( Id8ce8f636723b9f119bb86c25017e6b3[fgallag_SEL-1:0]),
.fgallag( Id2ed64cae3cb1e0ada8e3fb4ebb2dc78 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic1c911bc20d03275c7d20ab993e9a54d = (Id8ce8f636723b9f119bb86c25017e6b3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id2ed64cae3cb1e0ada8e3fb4ebb2dc78 ;

Ic9c2f173881d25f8976d723957809f51 Id8ba768211ca86d53bc4c586d4c12338 (
.fgallag_sel( Ic29a18d8d504a2d5280c1d7771346518[fgallag_SEL-1:0]),
.fgallag( I16b9849d3f2edd7f9ed7accb138d2c02 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iff207077a60c0196ac33f68e37d7d824 = (Ic29a18d8d504a2d5280c1d7771346518[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I16b9849d3f2edd7f9ed7accb138d2c02 ;

Ic9c2f173881d25f8976d723957809f51 I61dbd7b1f858e6643e9becbe40bd2401 (
.fgallag_sel( I96a79193aa2956b8f901d5fcc9cf65cf[fgallag_SEL-1:0]),
.fgallag( Ibcfe38455aa7aa33ae950172fb915dc5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0980811a7928bd72e415daf24b41137f = (I96a79193aa2956b8f901d5fcc9cf65cf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibcfe38455aa7aa33ae950172fb915dc5 ;

Ic9c2f173881d25f8976d723957809f51 I43812a122da4a767c14a2622f4153bab (
.fgallag_sel( I8c97a246c749fbef029f8b1671c772bd[fgallag_SEL-1:0]),
.fgallag( Ic9d9832294a3707b4041b2c4d8f92615 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie5a8e0e3d35d27fbb680552444f2ae65 = (I8c97a246c749fbef029f8b1671c772bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic9d9832294a3707b4041b2c4d8f92615 ;

Ic9c2f173881d25f8976d723957809f51 Ib150fbd0120b2bb9b532b1306cf5e2df (
.fgallag_sel( If9ba9d221909ce7499725f6fd7d519f8[fgallag_SEL-1:0]),
.fgallag( I3ef9641c53e7aa6a588481b57b865aa3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I91e4dd08f282857ab4c275bb1441c9d7 = (If9ba9d221909ce7499725f6fd7d519f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3ef9641c53e7aa6a588481b57b865aa3 ;

Ic9c2f173881d25f8976d723957809f51 I11266d7179f7f0f311d8432a3a691d0b (
.fgallag_sel( I53a7878f44253f0f1a82d9d27b1a44c3[fgallag_SEL-1:0]),
.fgallag( Ie838f76c6fc041e4fa66441094ae477c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iea26a1265fd6c48c038993b2038d2747 = (I53a7878f44253f0f1a82d9d27b1a44c3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie838f76c6fc041e4fa66441094ae477c ;

Ic9c2f173881d25f8976d723957809f51 If97f66f5e16bba57e0fb9f9a1dd042e5 (
.fgallag_sel( Ie0e928125f9d3d17d123d97e00f1fc34[fgallag_SEL-1:0]),
.fgallag( Ice9f8149ed08f537da5e146b417085e0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7920256f397f35450287256339769d4b = (Ie0e928125f9d3d17d123d97e00f1fc34[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ice9f8149ed08f537da5e146b417085e0 ;

Ic9c2f173881d25f8976d723957809f51 Ic00396f526a70c0975a4aa272b151cdd (
.fgallag_sel( I2bd0f77efeca09eebe82ea234e9fe638[fgallag_SEL-1:0]),
.fgallag( I71f6bd2fe34731aab306cfb89a3335ca ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibad06757b56b14755f0e50620a53dc6c = (I2bd0f77efeca09eebe82ea234e9fe638[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I71f6bd2fe34731aab306cfb89a3335ca ;

Ic9c2f173881d25f8976d723957809f51 Ie3e81cc439ad0e00e7107a9ce94b5d69 (
.fgallag_sel( I94f2e7ef9b3463bd598dc9049f6fb0ef[fgallag_SEL-1:0]),
.fgallag( I5dd57cfd0d7ce83fcbdb3f560ac713fb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id76592cbf9ad537e9cab20469c5e5861 = (I94f2e7ef9b3463bd598dc9049f6fb0ef[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5dd57cfd0d7ce83fcbdb3f560ac713fb ;

Ic9c2f173881d25f8976d723957809f51 If1c59b70218adcc4229f1440ef552cf7 (
.fgallag_sel( I6dc16510af6b61b79b339d0fce77ac24[fgallag_SEL-1:0]),
.fgallag( I239498228bdcb1c2a8b2cbef48e850a6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibc80d98586cca13a6849ae053b68e5fb = (I6dc16510af6b61b79b339d0fce77ac24[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I239498228bdcb1c2a8b2cbef48e850a6 ;

Ic9c2f173881d25f8976d723957809f51 I31769faff97b38b0f7004868f0888951 (
.fgallag_sel( Ic655e213ab81f5d61a018d3ed7016b12[fgallag_SEL-1:0]),
.fgallag( I82fc4233a3d2840670eb9b9adf6c9215 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I257237e7bef8b0e4cb27bc9a3a93aba6 = (Ic655e213ab81f5d61a018d3ed7016b12[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I82fc4233a3d2840670eb9b9adf6c9215 ;

Ic9c2f173881d25f8976d723957809f51 Ied7a4789cf3b2d3e8a96b5c39c0c75c5 (
.fgallag_sel( I2ffc4a604025a2f5c4e273c1d070a725[fgallag_SEL-1:0]),
.fgallag( Ieb08f6a94aa827632606608d014e26d3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1980cdd5ecb000134e55f507f369af66 = (I2ffc4a604025a2f5c4e273c1d070a725[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ieb08f6a94aa827632606608d014e26d3 ;

Ic9c2f173881d25f8976d723957809f51 I14c7ec0bc342b579a7e818f9298aa10d (
.fgallag_sel( I1c76818a9a3b688ca897aa479f7d807f[fgallag_SEL-1:0]),
.fgallag( Ifdbb9947713ac574738236fcb5c6ae07 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id0efde1d7f80f8848613c26fa4637c37 = (I1c76818a9a3b688ca897aa479f7d807f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifdbb9947713ac574738236fcb5c6ae07 ;

Ic9c2f173881d25f8976d723957809f51 I2777190ac4dfdcd2f0b0e1d5a94071eb (
.fgallag_sel( I3bfee9d3d88f0569010a4e0101200c19[fgallag_SEL-1:0]),
.fgallag( Ia737ee8f2c01feba1db87fe3e1a2388c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I76952d4ed281844c1c1795290b1ddc05 = (I3bfee9d3d88f0569010a4e0101200c19[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia737ee8f2c01feba1db87fe3e1a2388c ;

Ic9c2f173881d25f8976d723957809f51 I4a6224c8841532de975d2d596c83d26d (
.fgallag_sel( I5d4738755a26beb6d0f61dd3dec0f804[fgallag_SEL-1:0]),
.fgallag( I5d8e065dba640832d9d8db3e4338fbb5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7fa89ba905b099ebafe001878c4f0bed = (I5d4738755a26beb6d0f61dd3dec0f804[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5d8e065dba640832d9d8db3e4338fbb5 ;

Ic9c2f173881d25f8976d723957809f51 Ib1b5bff1b96263da86083441dca298e4 (
.fgallag_sel( I2f3c800091275bcb72d1a2a38fba53f3[fgallag_SEL-1:0]),
.fgallag( I3b3e36ffb1cff2c07bc9a61afdde10c1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icd841b02588f755a3133b72f8c625897 = (I2f3c800091275bcb72d1a2a38fba53f3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3b3e36ffb1cff2c07bc9a61afdde10c1 ;

Ic9c2f173881d25f8976d723957809f51 Ib553c63f670a9ce1c4140682da9ecec9 (
.fgallag_sel( I378e67cca7c4ff6325683f8346963210[fgallag_SEL-1:0]),
.fgallag( I2c8137e5ee04a1067858d7bb8d09d65b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I52945b9d986280c3dab4248e69247005 = (I378e67cca7c4ff6325683f8346963210[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2c8137e5ee04a1067858d7bb8d09d65b ;

Ic9c2f173881d25f8976d723957809f51 I97b41184507ef0d2d15409b9c9a7e317 (
.fgallag_sel( I04c8915a7f4bbde003f7facc84435c1a[fgallag_SEL-1:0]),
.fgallag( I38eb22d29ad9f4192499980fc17898b4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia0319e76fc112b3457f20662a7a51603 = (I04c8915a7f4bbde003f7facc84435c1a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I38eb22d29ad9f4192499980fc17898b4 ;

Ic9c2f173881d25f8976d723957809f51 Ib5b7012b5f65fe1e946a3617e1fc7bcc (
.fgallag_sel( I3f50b10072f38b6addee6845e6df9118[fgallag_SEL-1:0]),
.fgallag( Ib714941df0aaca40e7573e030d97b3f1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7a82bbf1146a3c68f01abf488a2e3c8f = (I3f50b10072f38b6addee6845e6df9118[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib714941df0aaca40e7573e030d97b3f1 ;

Ic9c2f173881d25f8976d723957809f51 I8475df925c5d296ba5b5b9be32079563 (
.fgallag_sel( Icc60eb18ba740036d2a17f98f15cfb98[fgallag_SEL-1:0]),
.fgallag( I47bcab5b082a8ce6312244224c162d39 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I05b26dca2316a9d527da24deb63c4756 = (Icc60eb18ba740036d2a17f98f15cfb98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I47bcab5b082a8ce6312244224c162d39 ;

Ic9c2f173881d25f8976d723957809f51 I9f45a1e89a686cd30228644e489f0d31 (
.fgallag_sel( I1677daa18aa8b226753b1a887b9420d1[fgallag_SEL-1:0]),
.fgallag( I68ded74f52dbd02ceb1da62a79d619d2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I256d84c23de18bd9a03cb41c0e3e4b8e = (I1677daa18aa8b226753b1a887b9420d1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I68ded74f52dbd02ceb1da62a79d619d2 ;

Ic9c2f173881d25f8976d723957809f51 I27da45a97528db12fa8d2626286ac0e2 (
.fgallag_sel( I36bc2d4c9a4480daa9b0944c08b50738[fgallag_SEL-1:0]),
.fgallag( Iaa113fd5f1e0c51d9f47240fe81b5604 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I619aafd5767c45229765838152161b71 = (I36bc2d4c9a4480daa9b0944c08b50738[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaa113fd5f1e0c51d9f47240fe81b5604 ;

Ic9c2f173881d25f8976d723957809f51 Ice02caf7ee55112718cb0149270298b3 (
.fgallag_sel( I38419a6905f50135a6783aacca0384dd[fgallag_SEL-1:0]),
.fgallag( I907bf413f65fad54303751c054687b29 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4bbb9f6eb1d79d41c7b5d61df854bd16 = (I38419a6905f50135a6783aacca0384dd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I907bf413f65fad54303751c054687b29 ;

Ic9c2f173881d25f8976d723957809f51 I5c3fa29765b477c8a995f2e1e8c2b1a4 (
.fgallag_sel( Ib48892dcb0715987289662a14672611e[fgallag_SEL-1:0]),
.fgallag( I7b727f2e9454f90d4fa4ef2cf69ddf23 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I997c88ff27fe957ec35a2b7146dd56f0 = (Ib48892dcb0715987289662a14672611e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7b727f2e9454f90d4fa4ef2cf69ddf23 ;

Ic9c2f173881d25f8976d723957809f51 I2634c19e4e8a043866fcf0d1e4e84476 (
.fgallag_sel( Icd9c94f929dbc71c9b836fda3019630b[fgallag_SEL-1:0]),
.fgallag( I6fc1f37134064dd7514b46ce7d27ceaa ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ide7fdb7a17f3d99a7840a648e0873bec = (Icd9c94f929dbc71c9b836fda3019630b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6fc1f37134064dd7514b46ce7d27ceaa ;

Ic9c2f173881d25f8976d723957809f51 I60a417a83848a27de2fda7a4a155b889 (
.fgallag_sel( I5d0249d9a772805b3fba3f3c7f5d35bd[fgallag_SEL-1:0]),
.fgallag( I7856585e0374651fc5f9921f69706a0b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I93dc025ca2d2cc3002c62c5d2e13d45b = (I5d0249d9a772805b3fba3f3c7f5d35bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7856585e0374651fc5f9921f69706a0b ;

Ic9c2f173881d25f8976d723957809f51 I31540e175158f7ea0e4ccbe8d03ae73e (
.fgallag_sel( Ie97341deb6fb24d49eb8b96bd0fd3f35[fgallag_SEL-1:0]),
.fgallag( I79b1967c2128c611ee4fe0d14bced1f4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9c656300bb176deba4be8400371f0ef2 = (Ie97341deb6fb24d49eb8b96bd0fd3f35[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I79b1967c2128c611ee4fe0d14bced1f4 ;

Ic9c2f173881d25f8976d723957809f51 I99824346afc8254abad0d1f534acaca9 (
.fgallag_sel( I17dd788f9d8e91307b6b1ab7488f9ce2[fgallag_SEL-1:0]),
.fgallag( Ib8aeaf62789d1d7a5a23d7492ff551b2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I141a53fdaada1994dc38d694fd03b5e3 = (I17dd788f9d8e91307b6b1ab7488f9ce2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib8aeaf62789d1d7a5a23d7492ff551b2 ;

Ic9c2f173881d25f8976d723957809f51 I80c48cdcf3a520d4b63cff1efa99f02f (
.fgallag_sel( I92ae370022ed107b152b10fd0aa3d2b7[fgallag_SEL-1:0]),
.fgallag( I9a8e8c3ce2c6323acee0877d445a2268 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1d81174ecfb84b8c906126d13900178e = (I92ae370022ed107b152b10fd0aa3d2b7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9a8e8c3ce2c6323acee0877d445a2268 ;

Ic9c2f173881d25f8976d723957809f51 Icb3b859203f402007b525e1f5b907b34 (
.fgallag_sel( Iebb39f0d19ec1208bbfba6cf67a3bfc7[fgallag_SEL-1:0]),
.fgallag( I701a3c05ad8e6ac5cea30b78707e77d1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I92ab5c30a7bfae4e698a74d2e48cde1a = (Iebb39f0d19ec1208bbfba6cf67a3bfc7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I701a3c05ad8e6ac5cea30b78707e77d1 ;

Ic9c2f173881d25f8976d723957809f51 I39529ea984c07211e313289db95ad0e9 (
.fgallag_sel( I81861f6bb8bbbab6e93407cfb4a852b8[fgallag_SEL-1:0]),
.fgallag( I75fefd09122859510021931c16051262 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifd41e7ed8ef5fa870c1abf043b5d5f2d = (I81861f6bb8bbbab6e93407cfb4a852b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I75fefd09122859510021931c16051262 ;

Ic9c2f173881d25f8976d723957809f51 Ic49849a1655995525aaa95764929269c (
.fgallag_sel( I217b2e3ca0a534fc5b1910adf3c1b57d[fgallag_SEL-1:0]),
.fgallag( I2779af0ff280ea511af850df795d1fb6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I983825ee77db3cbd86c937e5fe4707fd = (I217b2e3ca0a534fc5b1910adf3c1b57d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2779af0ff280ea511af850df795d1fb6 ;

Ic9c2f173881d25f8976d723957809f51 I9e1d70715a325f2b502187700938220b (
.fgallag_sel( I8429b08891dc56af24c72ce1b7725457[fgallag_SEL-1:0]),
.fgallag( I2eb84b0b6b12b9269bb791ae03e5094d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I715efc0ca41f678f8c582aaa3f255767 = (I8429b08891dc56af24c72ce1b7725457[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2eb84b0b6b12b9269bb791ae03e5094d ;

Ic9c2f173881d25f8976d723957809f51 I592bc17b3ae75c561b4c3ae06ec6832e (
.fgallag_sel( If96747262303f6c5c6b129e39224bd23[fgallag_SEL-1:0]),
.fgallag( Ie42cb87efb2b87d88eed6139132bb23e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I764815deb8bceeb1b9929de2dfd46235 = (If96747262303f6c5c6b129e39224bd23[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie42cb87efb2b87d88eed6139132bb23e ;

Ic9c2f173881d25f8976d723957809f51 I4fd87d2f96e137b5ba7c1c708db58b8b (
.fgallag_sel( If7012457af15c405baeaa1710319b541[fgallag_SEL-1:0]),
.fgallag( Id2e2722999e300df1bc7ea89dbf5689d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1b869d6b94307bc9bea28db11161e61e = (If7012457af15c405baeaa1710319b541[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id2e2722999e300df1bc7ea89dbf5689d ;

Ic9c2f173881d25f8976d723957809f51 I0501d0cc5dc53d5d943c1ce545fd215a (
.fgallag_sel( Ia0a0229ef71b85195352bb664ea4e4e3[fgallag_SEL-1:0]),
.fgallag( I2b7e1a65c52821f3f7e194a443b0117d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idf695c6735d8d8aafa37ad4cbd5a5872 = (Ia0a0229ef71b85195352bb664ea4e4e3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2b7e1a65c52821f3f7e194a443b0117d ;

Ic9c2f173881d25f8976d723957809f51 Iadb8d540e77d09f8c1d03c26d995d449 (
.fgallag_sel( I42aeb7c23accc2ca874c7f8221c3af93[fgallag_SEL-1:0]),
.fgallag( I8b31aa4edbc800c99628c5851cad8770 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib9114ddde15c1908595081b52ba00c48 = (I42aeb7c23accc2ca874c7f8221c3af93[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8b31aa4edbc800c99628c5851cad8770 ;

Ic9c2f173881d25f8976d723957809f51 I47952c07f1118a0f3273d7e61aed15c9 (
.fgallag_sel( I7df6a95bf51f40693c439c6df36510d4[fgallag_SEL-1:0]),
.fgallag( Id40d461c28ecc2017d9b7d2eadf5ea44 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3d52a609547a0ac3cd6d0481f09d00f2 = (I7df6a95bf51f40693c439c6df36510d4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id40d461c28ecc2017d9b7d2eadf5ea44 ;

Ic9c2f173881d25f8976d723957809f51 Idf8e5464571f598b08988067d8c43e9f (
.fgallag_sel( I8fe65f9c344d7ec8657f192abefc3fb6[fgallag_SEL-1:0]),
.fgallag( I4b8f58440e6848610f2e7e06efbc64fe ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I45abcbcdc3951ebaef039e6cb2562d4d = (I8fe65f9c344d7ec8657f192abefc3fb6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4b8f58440e6848610f2e7e06efbc64fe ;

Ic9c2f173881d25f8976d723957809f51 Idc11ca5ea4dadb092c48dbeb9b2f8e31 (
.fgallag_sel( I4d75c95d34d8d8aeeb528456bbe136e1[fgallag_SEL-1:0]),
.fgallag( Ica1d5cc8dc277e91787ec1bf0f2ed65c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5bed8ad020614972a82bf3ad66300f12 = (I4d75c95d34d8d8aeeb528456bbe136e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ica1d5cc8dc277e91787ec1bf0f2ed65c ;

Ic9c2f173881d25f8976d723957809f51 Ie27de266f957d347c02bcf708d4e342f (
.fgallag_sel( I43746054a38c9521f8da9db9d0e91f99[fgallag_SEL-1:0]),
.fgallag( Ie5d481ac7a371e1fd3c48c5cf9649a67 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic7ec84d03001998a8504a79afb1f0d5c = (I43746054a38c9521f8da9db9d0e91f99[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie5d481ac7a371e1fd3c48c5cf9649a67 ;

Ic9c2f173881d25f8976d723957809f51 I7c2a4aded3c855f2e4102a5039ef1841 (
.fgallag_sel( I0430ac2a4b2b2e2fc7f8154bf946553c[fgallag_SEL-1:0]),
.fgallag( I9786bf468ba8540d7e75d762fc832709 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I43cfed51e8dec917304dff4f44a984c6 = (I0430ac2a4b2b2e2fc7f8154bf946553c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9786bf468ba8540d7e75d762fc832709 ;

Ic9c2f173881d25f8976d723957809f51 I50db012203a53a2a4724ea1ab3b987d8 (
.fgallag_sel( I25dc807fd55b81c9f24fd0d1edcaa758[fgallag_SEL-1:0]),
.fgallag( Ib093fabefab0a1b46d2199c1c948abc8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If34baa3a92291d91308582e9c268ccaf = (I25dc807fd55b81c9f24fd0d1edcaa758[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib093fabefab0a1b46d2199c1c948abc8 ;

Ic9c2f173881d25f8976d723957809f51 If72140e2897efa05621361021f538352 (
.fgallag_sel( I7881184f1779b9fd4fdf329c5f7664da[fgallag_SEL-1:0]),
.fgallag( I9b53bbb22003297175c6c4655ef83c93 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8c00e1f1c7faa04600505a6f30e32ccc = (I7881184f1779b9fd4fdf329c5f7664da[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9b53bbb22003297175c6c4655ef83c93 ;

Ic9c2f173881d25f8976d723957809f51 Ieff640e15923eb02a7ee48e957838466 (
.fgallag_sel( I8e6de2d692a307ee8a5a4b2a9265a633[fgallag_SEL-1:0]),
.fgallag( I9df2a441fadba7dc49effc5eecf4b0e8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I225a03b34b73fee071973985a66f9213 = (I8e6de2d692a307ee8a5a4b2a9265a633[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9df2a441fadba7dc49effc5eecf4b0e8 ;

Ic9c2f173881d25f8976d723957809f51 Ie3e8e5a8f8eacdb842398d334d2ae443 (
.fgallag_sel( I54b2b18ab051b468808a3d0fc4bc893f[fgallag_SEL-1:0]),
.fgallag( I102372ac8a06119e5d827d83f172bbd2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4b819b7da7ced2a32e77b3b26682168f = (I54b2b18ab051b468808a3d0fc4bc893f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I102372ac8a06119e5d827d83f172bbd2 ;

Ic9c2f173881d25f8976d723957809f51 I9e26ebc8a526bfd31a6126445a3b2c59 (
.fgallag_sel( I37ee86e2ca32832862cb57efe76bbedf[fgallag_SEL-1:0]),
.fgallag( I5cad4cd564b0956b08f22cd42d594b01 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3d1050efa384172a3af1fa5f259a3877 = (I37ee86e2ca32832862cb57efe76bbedf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5cad4cd564b0956b08f22cd42d594b01 ;

Ic9c2f173881d25f8976d723957809f51 I07694564445cf74dfc16c7e61e4c472c (
.fgallag_sel( Ic95f2fc697574803c0f7fa35c2609f0c[fgallag_SEL-1:0]),
.fgallag( Id685ced1c37d97c75b49b2f790dbabad ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I66de52bc354a661ccda6f4d6d744bfdf = (Ic95f2fc697574803c0f7fa35c2609f0c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id685ced1c37d97c75b49b2f790dbabad ;

Ic9c2f173881d25f8976d723957809f51 Ie273f846f8e27fbc9e1f9b4182b58494 (
.fgallag_sel( I933a30c52c9bec5172530b2d739a3b63[fgallag_SEL-1:0]),
.fgallag( I219e400c87948e7b2bf715745a4b152c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib9a88f5ea722553569167ca7b186fd50 = (I933a30c52c9bec5172530b2d739a3b63[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I219e400c87948e7b2bf715745a4b152c ;

Ic9c2f173881d25f8976d723957809f51 I44178ef2909991a576dda469f29c121b (
.fgallag_sel( I7bbd7df18f85197c22fe8cfe37312af6[fgallag_SEL-1:0]),
.fgallag( I3372567dacc350adf991928753209605 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I68904155ce7e8d722b67725f81af7f06 = (I7bbd7df18f85197c22fe8cfe37312af6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3372567dacc350adf991928753209605 ;

Ic9c2f173881d25f8976d723957809f51 Ic7a05ac13da7b88422ab1fffc4d2eebc (
.fgallag_sel( I50d5ada7c91c7af16492c6b41151b68f[fgallag_SEL-1:0]),
.fgallag( Ibf50476ac553bceaedcb121b28093394 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7bc807d9f1b67d68e11c8a064b218963 = (I50d5ada7c91c7af16492c6b41151b68f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibf50476ac553bceaedcb121b28093394 ;

Ic9c2f173881d25f8976d723957809f51 I6c9939132719e67e6576c4181ed5ab56 (
.fgallag_sel( I32c8e7996b3473d4906c40018799a16b[fgallag_SEL-1:0]),
.fgallag( I5d20fcccde5844e36b83d7fd7034c413 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id1b5740fd8ce883d3cf724bd7410f27e = (I32c8e7996b3473d4906c40018799a16b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5d20fcccde5844e36b83d7fd7034c413 ;

Ic9c2f173881d25f8976d723957809f51 I8a00e756b6f25c9085a1b27a9191b0d3 (
.fgallag_sel( Ic0eacd5a4812ad7ae3fa251ab2db4694[fgallag_SEL-1:0]),
.fgallag( I47e720341773b3a11f4c71b4e9644525 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I12c6efa1dbc88f222ebcb8866946eea1 = (Ic0eacd5a4812ad7ae3fa251ab2db4694[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I47e720341773b3a11f4c71b4e9644525 ;

Ic9c2f173881d25f8976d723957809f51 I0b58788fb0deda5447289fd246c03bb3 (
.fgallag_sel( Ideecf8ab87d28a840cd93851169ab05b[fgallag_SEL-1:0]),
.fgallag( I0251d8ecec82a24878ce494f0b417ce3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9c9d28abad8610fa2cecb74d18a1c9e3 = (Ideecf8ab87d28a840cd93851169ab05b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0251d8ecec82a24878ce494f0b417ce3 ;

Ic9c2f173881d25f8976d723957809f51 Id973fd1b3cd14f4e7a331627682a5ebd (
.fgallag_sel( I1ac6775eb38457b7962241d2e7336b0d[fgallag_SEL-1:0]),
.fgallag( Ibeef795b2235c98439628da8d7c094e0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I21af49923adfeca8b24188a7bba54b1d = (I1ac6775eb38457b7962241d2e7336b0d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibeef795b2235c98439628da8d7c094e0 ;

Ic9c2f173881d25f8976d723957809f51 I292915f604600a834b060bf6c72e41d5 (
.fgallag_sel( I2ecaa89698604fddd863d7e28d643a57[fgallag_SEL-1:0]),
.fgallag( I61769f7c08a0b9cf78068455410b6bb2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I46c921b6dbb398813ad0d6c06e2eb33a = (I2ecaa89698604fddd863d7e28d643a57[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I61769f7c08a0b9cf78068455410b6bb2 ;

Ic9c2f173881d25f8976d723957809f51 Ia77ffed02e5c6f5303b63432baba7dd3 (
.fgallag_sel( I273e0fe9c51c8549c8dfff393ca2e4e1[fgallag_SEL-1:0]),
.fgallag( I77fe52c685b1075c294ac3c0a5b0d63a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifa087dd71378f388142d351fa18806b5 = (I273e0fe9c51c8549c8dfff393ca2e4e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I77fe52c685b1075c294ac3c0a5b0d63a ;

Ic9c2f173881d25f8976d723957809f51 I20e7b39d7d91ba3d04dd395b00e0f868 (
.fgallag_sel( Ifb1fc76002f6920a1f44c7b1bbcd0020[fgallag_SEL-1:0]),
.fgallag( Ia688029a35b4a62417906c9aa1cd7719 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3f3c345d02438bc96a1f7b162315ea43 = (Ifb1fc76002f6920a1f44c7b1bbcd0020[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia688029a35b4a62417906c9aa1cd7719 ;

Ic9c2f173881d25f8976d723957809f51 I7cd22d14fb985f7b77d8a5376841d6e0 (
.fgallag_sel( Idf6d4e3aa753aa396a9bffb27732f851[fgallag_SEL-1:0]),
.fgallag( Ifaaab2c6f368b133936a7295eeb9b45d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7577c4409a32ebf50e5a187f71c84b1e = (Idf6d4e3aa753aa396a9bffb27732f851[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifaaab2c6f368b133936a7295eeb9b45d ;

Ic9c2f173881d25f8976d723957809f51 I6f1b479a2d953e6e7531bf736e9519f6 (
.fgallag_sel( If14ca1f5d1c2977f9da79eaebaad1bf9[fgallag_SEL-1:0]),
.fgallag( Ifbe064ac0a5f4bbf6caae486064a983d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iec97b82162ff77d0b123feeb5b5904e6 = (If14ca1f5d1c2977f9da79eaebaad1bf9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifbe064ac0a5f4bbf6caae486064a983d ;

Ic9c2f173881d25f8976d723957809f51 I59d1fc4a759ba792b85159a90048ff75 (
.fgallag_sel( If8f1505d9f10e30bd3320f500d34932f[fgallag_SEL-1:0]),
.fgallag( I439ac39c831e0ca87a40f49e439ce24f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2206f864d477e44a18769ea9cc01d8ee = (If8f1505d9f10e30bd3320f500d34932f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I439ac39c831e0ca87a40f49e439ce24f ;

Ic9c2f173881d25f8976d723957809f51 I3f83d4605c6ba082c674649ee057d7b3 (
.fgallag_sel( Id32aa77c6406b35a00168bb5452b12fb[fgallag_SEL-1:0]),
.fgallag( I5c616021ebd98fc8e0fcf5b19732175c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9b67c7138cc6e8c9ef36b5cb28932c9e = (Id32aa77c6406b35a00168bb5452b12fb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5c616021ebd98fc8e0fcf5b19732175c ;

Ic9c2f173881d25f8976d723957809f51 I707c4c77d2ec237be5a2de561a2029c5 (
.fgallag_sel( I9a73686acefeb361337511f6943b036b[fgallag_SEL-1:0]),
.fgallag( Id3a6c8114a92efaf5f6c280f897bef71 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic295c2717dcc256113776b8d39368802 = (I9a73686acefeb361337511f6943b036b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id3a6c8114a92efaf5f6c280f897bef71 ;

Ic9c2f173881d25f8976d723957809f51 I7a9baa4356bc69441b6c68acbbbb1d3f (
.fgallag_sel( Ib6eb7ce5a070f3a87bcf0e18be8c855d[fgallag_SEL-1:0]),
.fgallag( I854d4e2867b459da2e2fc06c438e6077 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4875abaa409c919efee2cde0c90e1e7d = (Ib6eb7ce5a070f3a87bcf0e18be8c855d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I854d4e2867b459da2e2fc06c438e6077 ;

Ic9c2f173881d25f8976d723957809f51 I0cf4be14e112d7f7622eb6d5a4f52a5f (
.fgallag_sel( If69b0b717c35d33fc8c0e59b07eb9edc[fgallag_SEL-1:0]),
.fgallag( I3b334e8064cbfe97e70a0f4055496f04 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0bcc0953acf369ba9571d11e68511af4 = (If69b0b717c35d33fc8c0e59b07eb9edc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3b334e8064cbfe97e70a0f4055496f04 ;

Ic9c2f173881d25f8976d723957809f51 I9ed910ce6d1d77c8c99875d1f63ef0b6 (
.fgallag_sel( Ibb0d73078b779585e6b0e228391ecb96[fgallag_SEL-1:0]),
.fgallag( Iff92d12470884efa033800c88e1983e3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4d92612c245b6ebb246d2f41b3dd4107 = (Ibb0d73078b779585e6b0e228391ecb96[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iff92d12470884efa033800c88e1983e3 ;

Ic9c2f173881d25f8976d723957809f51 Ia2ef95c545fda7b113c6ce231371c3ec (
.fgallag_sel( I2894546e399fe3e33d7579772a1310df[fgallag_SEL-1:0]),
.fgallag( I3d167f5af41902dc0a6477d55cf0abfd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I53a8be01a8f8067f67e0498c48cfa2a8 = (I2894546e399fe3e33d7579772a1310df[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3d167f5af41902dc0a6477d55cf0abfd ;

Ic9c2f173881d25f8976d723957809f51 I397873aa72d2a1d103a44e752afc1898 (
.fgallag_sel( I97f99a266267859aed199b278a430417[fgallag_SEL-1:0]),
.fgallag( Iaa7edba3767735cad1ec76479b5548b0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I036d8ab76c1f8c3b52ddcad50c6c8a6c = (I97f99a266267859aed199b278a430417[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaa7edba3767735cad1ec76479b5548b0 ;

Ic9c2f173881d25f8976d723957809f51 I89288af78822fa4fb393507ca87844d5 (
.fgallag_sel( Ie18cc792329941a3654322376a937d8d[fgallag_SEL-1:0]),
.fgallag( Ifaa7aff0fb2af9d3e04b2641b13cf884 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idaffa51af26a79990b50e9422da6074c = (Ie18cc792329941a3654322376a937d8d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifaa7aff0fb2af9d3e04b2641b13cf884 ;

Ic9c2f173881d25f8976d723957809f51 I8d10e837b2579ba62aa9c6009a7bfc71 (
.fgallag_sel( Ie914a99f08d60b74c3c36a632a4ca9b0[fgallag_SEL-1:0]),
.fgallag( Ia78b9e9a1faddb38b4a1472f5eea3939 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia17748dd92434f8658e49a3f7ed682e8 = (Ie914a99f08d60b74c3c36a632a4ca9b0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia78b9e9a1faddb38b4a1472f5eea3939 ;

Ic9c2f173881d25f8976d723957809f51 Ibdfae7538c74199abf96b1eae8fe465c (
.fgallag_sel( I82916e9dc3894ad88e12de01a68d6aa5[fgallag_SEL-1:0]),
.fgallag( I367d25430d8ec417123931f9534f3eba ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1ecdfded32659bd57c752928f0cc12eb = (I82916e9dc3894ad88e12de01a68d6aa5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I367d25430d8ec417123931f9534f3eba ;

Ic9c2f173881d25f8976d723957809f51 I9926e290e9960c698b1cc0cbc1e211b8 (
.fgallag_sel( I6cbf576b3d652e34c0221f8316b5a392[fgallag_SEL-1:0]),
.fgallag( I38a19bd51c6ee4fcb38493d869b7808a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If7bcd20651da485996362af6b633fec3 = (I6cbf576b3d652e34c0221f8316b5a392[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I38a19bd51c6ee4fcb38493d869b7808a ;

Ic9c2f173881d25f8976d723957809f51 I87631d8fbfc6f9af74a9233c82012aa6 (
.fgallag_sel( I9141b2516d7f855cd186472780af7b67[fgallag_SEL-1:0]),
.fgallag( I0fe662c7d5cce9cf3cac56b6125852ff ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7a04a2c4768a6703cb98c2adfd53088f = (I9141b2516d7f855cd186472780af7b67[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0fe662c7d5cce9cf3cac56b6125852ff ;

Ic9c2f173881d25f8976d723957809f51 I25ec622096b17f98ea417bc352f76130 (
.fgallag_sel( I07bf32ed72de9c02abf700c64853af61[fgallag_SEL-1:0]),
.fgallag( I6867bb41ee0a7f4c6ae0071e7975526d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iebc9456956b29940df3df4dddae0619f = (I07bf32ed72de9c02abf700c64853af61[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6867bb41ee0a7f4c6ae0071e7975526d ;

Ic9c2f173881d25f8976d723957809f51 Iedf384e273bee58a4a46675012959213 (
.fgallag_sel( I52663a2999fb9571834d517538691b6f[fgallag_SEL-1:0]),
.fgallag( I74d3dc7b6116f47b27dbfd112d7afd5d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iefb9092502c1c93656c9050bf74e6849 = (I52663a2999fb9571834d517538691b6f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I74d3dc7b6116f47b27dbfd112d7afd5d ;

Ic9c2f173881d25f8976d723957809f51 Id6772788be394846f0ec6df8a6838f45 (
.fgallag_sel( I8dcb88c94506367aabe8d7ed62cc56c2[fgallag_SEL-1:0]),
.fgallag( I13440021cb8441969d3242de4fc6a0b5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I42edf14a24cb1e19924e0f5531f97ed9 = (I8dcb88c94506367aabe8d7ed62cc56c2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I13440021cb8441969d3242de4fc6a0b5 ;

Ic9c2f173881d25f8976d723957809f51 If6845ac23c6b7a49e789cd8abf8fa507 (
.fgallag_sel( Ie676a4bee61154145391d9cc473fe91d[fgallag_SEL-1:0]),
.fgallag( Id3c71879c307df1390bbc60c55a5f249 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia332b7b61c57cee58ef4a1733da2afc6 = (Ie676a4bee61154145391d9cc473fe91d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id3c71879c307df1390bbc60c55a5f249 ;

Ic9c2f173881d25f8976d723957809f51 I8587d6b1627320e856a97de564f6ba9e (
.fgallag_sel( I9502c8fbf6b48749bf9f84a89a937dfe[fgallag_SEL-1:0]),
.fgallag( I2e1fa8e49bf48184e6a669d18f5c8ced ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib4450f5e900229ff87baede34be883b4 = (I9502c8fbf6b48749bf9f84a89a937dfe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2e1fa8e49bf48184e6a669d18f5c8ced ;

Ic9c2f173881d25f8976d723957809f51 Ibcc5a23109092b34dc5f8ba28ae14d0c (
.fgallag_sel( I0c91e540e7106f32ae59491d8ed1853e[fgallag_SEL-1:0]),
.fgallag( Ibc9c9339a0bcbc6addcce833051a8cd0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie7d8f527db720e17a73a57400a5360a5 = (I0c91e540e7106f32ae59491d8ed1853e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibc9c9339a0bcbc6addcce833051a8cd0 ;

Ic9c2f173881d25f8976d723957809f51 I8d131dfac0789022816bf35243812482 (
.fgallag_sel( Iddfb8a8e261389eb4a2a10880c19446a[fgallag_SEL-1:0]),
.fgallag( I2c0a2ad9eef6e84c60d1a6503aa836db ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7c420e9724fd4bc31071a57ac1ba5293 = (Iddfb8a8e261389eb4a2a10880c19446a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2c0a2ad9eef6e84c60d1a6503aa836db ;

Ic9c2f173881d25f8976d723957809f51 I460c7247611c77e6db33ac20f44831da (
.fgallag_sel( If0d55f861d4b3f0970c529024ca142d5[fgallag_SEL-1:0]),
.fgallag( I3b06c3a23b2068e8f45870524c4af870 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5a38174a83eaebe2678ca70fe5915c02 = (If0d55f861d4b3f0970c529024ca142d5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3b06c3a23b2068e8f45870524c4af870 ;

Ic9c2f173881d25f8976d723957809f51 I39993aec2352bdb693485fe6417f58c8 (
.fgallag_sel( Ib054f5d3f5cbb29a053d0e50c23cb3a8[fgallag_SEL-1:0]),
.fgallag( I87d44c01b261e9c13add415e6b3cc5ba ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib3639c700fe97648415fd4dfc8a6466b = (Ib054f5d3f5cbb29a053d0e50c23cb3a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I87d44c01b261e9c13add415e6b3cc5ba ;

Ic9c2f173881d25f8976d723957809f51 I7ad151742feaa8b0b5cf9611ccd62bc8 (
.fgallag_sel( I1d65e9f97e93de8cc2a5dd532f8e482a[fgallag_SEL-1:0]),
.fgallag( Ifc15e0dd91741676f23cc20fc542ec14 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5228b59565a0ae5f56237e5332ddefa1 = (I1d65e9f97e93de8cc2a5dd532f8e482a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifc15e0dd91741676f23cc20fc542ec14 ;

Ic9c2f173881d25f8976d723957809f51 I162b760665dabb5fcd40572a2e8db68d (
.fgallag_sel( I3bdeab8c87325d46e45d9e2d44756934[fgallag_SEL-1:0]),
.fgallag( I50fdfffb4e2dbcf33282b3653f595ad0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I87188c070d52012c107a5b37e718a5d4 = (I3bdeab8c87325d46e45d9e2d44756934[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I50fdfffb4e2dbcf33282b3653f595ad0 ;

Ic9c2f173881d25f8976d723957809f51 I4c0f0e7da97042b9b52f5dc70cba3d7d (
.fgallag_sel( If9228f7ecf19c41f4bbd8dabd0d5816c[fgallag_SEL-1:0]),
.fgallag( I4e9786ec39d388cdce110c86bb436ae3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7d0ebb3f7a7e77362b41f9ec9b98c9af = (If9228f7ecf19c41f4bbd8dabd0d5816c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4e9786ec39d388cdce110c86bb436ae3 ;

Ic9c2f173881d25f8976d723957809f51 I42894dc8979482b884c79acdcc6dd17f (
.fgallag_sel( I9e3edee214c4937d2aa462d3cffa624b[fgallag_SEL-1:0]),
.fgallag( I47cb30eb341ae7ce99042a16cd109f26 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1c2e01ba53fb12e4c3e44e4a9ef97888 = (I9e3edee214c4937d2aa462d3cffa624b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I47cb30eb341ae7ce99042a16cd109f26 ;

Ic9c2f173881d25f8976d723957809f51 I7f093686b1cb09ab8d26de12f771332f (
.fgallag_sel( I9fcbbd2e81b006b50e2d35ed2627bf83[fgallag_SEL-1:0]),
.fgallag( If004fa1c4e6bbe1f458c2d2a4f1f6e03 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icf7e609c4a537e6f2a7b86b7035717d3 = (I9fcbbd2e81b006b50e2d35ed2627bf83[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If004fa1c4e6bbe1f458c2d2a4f1f6e03 ;

Ic9c2f173881d25f8976d723957809f51 I9077205993ae3077102d5b0b12ccd573 (
.fgallag_sel( Ie16f3d50ad5e5581ca099549db7232d2[fgallag_SEL-1:0]),
.fgallag( I7c9910ade59c54e170c4f10822b5aff4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I39d74e21fb67539c0d310571b99a3e22 = (Ie16f3d50ad5e5581ca099549db7232d2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7c9910ade59c54e170c4f10822b5aff4 ;

Ic9c2f173881d25f8976d723957809f51 I9cdc8da954611d4c1849c93dd7f7af57 (
.fgallag_sel( I6345e93f3fa7f5eb2008dd41742afc2d[fgallag_SEL-1:0]),
.fgallag( I98939499dd98e583a4788cacc66c7fc4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I395b85e88acd203dd93e519710aea79b = (I6345e93f3fa7f5eb2008dd41742afc2d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I98939499dd98e583a4788cacc66c7fc4 ;

Ic9c2f173881d25f8976d723957809f51 Ied01a8add32e337bf27ca4f7be313487 (
.fgallag_sel( I698b93e10073b5d29357cde4bcac9dbe[fgallag_SEL-1:0]),
.fgallag( Ic530781e13180026815873e12550e405 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I850e5fd50416aaad26283152c4a49ddc = (I698b93e10073b5d29357cde4bcac9dbe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic530781e13180026815873e12550e405 ;

Ic9c2f173881d25f8976d723957809f51 Ia4f45373c924cec1e13e8e918bc4f741 (
.fgallag_sel( Ie7ced910d84655790823e6173a5a314a[fgallag_SEL-1:0]),
.fgallag( Iba43927cdbcb6a80953fced163686073 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ide38f5cac19b1bc82b26bfa12e5f9d8c = (Ie7ced910d84655790823e6173a5a314a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iba43927cdbcb6a80953fced163686073 ;

Ic9c2f173881d25f8976d723957809f51 I354ccd98ab7afe04839399551959e7bb (
.fgallag_sel( If6e3b6fd1810f6964e9024329d7cb3e3[fgallag_SEL-1:0]),
.fgallag( I29aefee3f95a7d2838ec5068515f69b0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib2d8874232a27b78a8c664e0fa2af512 = (If6e3b6fd1810f6964e9024329d7cb3e3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I29aefee3f95a7d2838ec5068515f69b0 ;

Ic9c2f173881d25f8976d723957809f51 I76e0eced0640a9508929678b7021a98e (
.fgallag_sel( If1045908c6d7476bd5507e57d08c406c[fgallag_SEL-1:0]),
.fgallag( Ib964c4dd0a0ce2553766251b73018699 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id002a482b2a09d2d17b9fa903882e8e0 = (If1045908c6d7476bd5507e57d08c406c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib964c4dd0a0ce2553766251b73018699 ;

Ic9c2f173881d25f8976d723957809f51 I6c676c51742a36f111ce2276513e093a (
.fgallag_sel( I4d4f6705ed77a16ff31b34bae0d8b6d9[fgallag_SEL-1:0]),
.fgallag( Ifd870cf74e7e3e5b348ad55af7242c27 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I359451948e89283ee89d89cebf689445 = (I4d4f6705ed77a16ff31b34bae0d8b6d9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifd870cf74e7e3e5b348ad55af7242c27 ;

Ic9c2f173881d25f8976d723957809f51 I4f8464d5a75dfd152fa59ff2173e6b0f (
.fgallag_sel( I70a492396580ac1143d8a2f4b181e873[fgallag_SEL-1:0]),
.fgallag( Ic4ba744721cdd747affca302b2b926d4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifffc8f779e22eedf06f7d1c24da411cb = (I70a492396580ac1143d8a2f4b181e873[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic4ba744721cdd747affca302b2b926d4 ;

Ic9c2f173881d25f8976d723957809f51 Ica65be9dae22def47ae9bbf3ffe9cba0 (
.fgallag_sel( I2fade32b5bdf245fa15289620dae2670[fgallag_SEL-1:0]),
.fgallag( Id381e35622a3ac2c549a8c9b702ec020 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3ccf7fbf7a13aef5daa7905b485d6e3a = (I2fade32b5bdf245fa15289620dae2670[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id381e35622a3ac2c549a8c9b702ec020 ;

Ic9c2f173881d25f8976d723957809f51 I04c5ca7b4cd3a0f8dd7b61a80d24e9ff (
.fgallag_sel( Ie0dc166f57fea074496241a32cdb6015[fgallag_SEL-1:0]),
.fgallag( If49e3943165e2782c928a7da86847145 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9deead4d27ef61f468a1bac90adfa27e = (Ie0dc166f57fea074496241a32cdb6015[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If49e3943165e2782c928a7da86847145 ;

Ic9c2f173881d25f8976d723957809f51 Ie267dd02019576044df476a137c52fd2 (
.fgallag_sel( If6a2518891412caa6d6d507082501f1e[fgallag_SEL-1:0]),
.fgallag( Ie4d85aa4951d1a918d698c9e411b1ab2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6c050a19b5031493dcc7163509b00012 = (If6a2518891412caa6d6d507082501f1e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie4d85aa4951d1a918d698c9e411b1ab2 ;

Ic9c2f173881d25f8976d723957809f51 Ic3210fe154f05486e7a3a188b5bea12e (
.fgallag_sel( Ic9912e5a838a377b26a19d22148a64df[fgallag_SEL-1:0]),
.fgallag( Iff6a8d4bc8f5f37d0ccc2d41f469ca86 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If74b57fb1d88f063bfef26ae6b74ff2d = (Ic9912e5a838a377b26a19d22148a64df[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iff6a8d4bc8f5f37d0ccc2d41f469ca86 ;

Ic9c2f173881d25f8976d723957809f51 Ib2f0d64b01274fd6a5763ffdd8eb12d5 (
.fgallag_sel( Ibc0fca22d16444bc17877106ca772c31[fgallag_SEL-1:0]),
.fgallag( I6bed9b6e8b499c11d719f869467d2322 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9fc7952b3920da1adf39777e9a1cd13f = (Ibc0fca22d16444bc17877106ca772c31[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6bed9b6e8b499c11d719f869467d2322 ;

Ic9c2f173881d25f8976d723957809f51 If652fad353e018a8af7cfd060f20194c (
.fgallag_sel( Ie4291d233597d5d676a80fd62d9bd208[fgallag_SEL-1:0]),
.fgallag( Id1db54a136ab42fe675fa77b2b7fd2de ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic013de8383ced83cb6cb368e54cd0f43 = (Ie4291d233597d5d676a80fd62d9bd208[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id1db54a136ab42fe675fa77b2b7fd2de ;

Ic9c2f173881d25f8976d723957809f51 If98d34e0cacd1bfaeb43d40f410ae1e0 (
.fgallag_sel( Ifc13b798d76aa70ec1877c275fb31d36[fgallag_SEL-1:0]),
.fgallag( Ia6ed9442d22d3228ce14749ffdacfab2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If71eac564bbca0cf2967a8803a24f586 = (Ifc13b798d76aa70ec1877c275fb31d36[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia6ed9442d22d3228ce14749ffdacfab2 ;

Ic9c2f173881d25f8976d723957809f51 I3dfe0c63f256569e12f3dded2454abee (
.fgallag_sel( I57d6637f0bdab578a790e4a12ccaa16b[fgallag_SEL-1:0]),
.fgallag( I32e0c22a86e88cadc6a956c213ff992c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib19bf2920a5486af62d38fa181293a47 = (I57d6637f0bdab578a790e4a12ccaa16b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I32e0c22a86e88cadc6a956c213ff992c ;

Ic9c2f173881d25f8976d723957809f51 Icb58911f3d1955e6931fd5a7a3c2dbe9 (
.fgallag_sel( If8ea04fe685b4f20cdaf9a84984d56fe[fgallag_SEL-1:0]),
.fgallag( I1b0dcddcb3e0a398857f038d3a52e719 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I92a94b468b025e5c1d103b2f8c92709e = (If8ea04fe685b4f20cdaf9a84984d56fe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1b0dcddcb3e0a398857f038d3a52e719 ;

Ic9c2f173881d25f8976d723957809f51 I0c2948b2874bdb26600e196dd96b6dc9 (
.fgallag_sel( Ie0c86f20c28bcbe410b191b90d29bf76[fgallag_SEL-1:0]),
.fgallag( I8c6bcabb8814607901102aca5f820293 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I76fe38786c53eb9f57d6512adb920d5b = (Ie0c86f20c28bcbe410b191b90d29bf76[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8c6bcabb8814607901102aca5f820293 ;

Ic9c2f173881d25f8976d723957809f51 I6adaf9688e4c4370c8c6acc63a5795c3 (
.fgallag_sel( I3dc5d3f66726e15968a70cbf3d3b656a[fgallag_SEL-1:0]),
.fgallag( I731089de22b5becf3621097ed7a81b7e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7878eb8ad885ea4193b8534015a445bb = (I3dc5d3f66726e15968a70cbf3d3b656a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I731089de22b5becf3621097ed7a81b7e ;

Ic9c2f173881d25f8976d723957809f51 Ibe99fbd7273bfc60e9728e9e60b0c75d (
.fgallag_sel( Id674686e7ac37fd6f63846f9a9cede19[fgallag_SEL-1:0]),
.fgallag( Ifb3674681315fa8cf6739996b823a7aa ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5b26270d07cd79afa7019dac72898e3c = (Id674686e7ac37fd6f63846f9a9cede19[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifb3674681315fa8cf6739996b823a7aa ;

Ic9c2f173881d25f8976d723957809f51 If98d73fbfab90ac514a4963a2e270f78 (
.fgallag_sel( Ie2ed9668d13d219c60f2e0614488cd42[fgallag_SEL-1:0]),
.fgallag( I2d5ef5bf9c28065a2a4ab718fbc8ba3e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I167dccb5e632afc0686602b35f9dea42 = (Ie2ed9668d13d219c60f2e0614488cd42[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2d5ef5bf9c28065a2a4ab718fbc8ba3e ;

Ic9c2f173881d25f8976d723957809f51 I0bc2ab815da6800d1e8b997a4b561815 (
.fgallag_sel( I98abc995ff89934534543be93c6e3ffa[fgallag_SEL-1:0]),
.fgallag( I7c5f9c301a0bdbf642f7b3f33e9bfc66 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3cb81e29fa5d50fadebe311acca6d090 = (I98abc995ff89934534543be93c6e3ffa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7c5f9c301a0bdbf642f7b3f33e9bfc66 ;

Ic9c2f173881d25f8976d723957809f51 I4b8ef74eb75ae916e024034f7bd88415 (
.fgallag_sel( I579cf9386ab7b08efa204d735335e462[fgallag_SEL-1:0]),
.fgallag( I7bde3bcef8556c1b1e4c7d2192196e00 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia25c11794a51c0937e0600032133a6dd = (I579cf9386ab7b08efa204d735335e462[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7bde3bcef8556c1b1e4c7d2192196e00 ;

Ic9c2f173881d25f8976d723957809f51 Ib380ffba08d50671a2d7973ce23e4326 (
.fgallag_sel( I9efa4d729d10a6b7cc335fb765ed032c[fgallag_SEL-1:0]),
.fgallag( Id13f3a39b334d8a80b7c8286b09bd1e1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I95b38f00928726b7b701405baf74f66a = (I9efa4d729d10a6b7cc335fb765ed032c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id13f3a39b334d8a80b7c8286b09bd1e1 ;

Ic9c2f173881d25f8976d723957809f51 I1584b70121c614eb778a24ebab16879d (
.fgallag_sel( If9191ebc8e88d4e75f0f35897ebb1421[fgallag_SEL-1:0]),
.fgallag( Ie6443f42260e0a2983927d0940c82a06 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I32c90cfef12eece5e90200ef79c7231f = (If9191ebc8e88d4e75f0f35897ebb1421[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie6443f42260e0a2983927d0940c82a06 ;

Ic9c2f173881d25f8976d723957809f51 I2780caaddcfe90e3169a03f34d78b9fb (
.fgallag_sel( I3511287cfe69d5cedc5a8fbcad708437[fgallag_SEL-1:0]),
.fgallag( I43003b2ef41b34363169f004a6668a59 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0b27fcbbc4514fa212fe3d023bdb526c = (I3511287cfe69d5cedc5a8fbcad708437[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I43003b2ef41b34363169f004a6668a59 ;

Ic9c2f173881d25f8976d723957809f51 I1a00eb4908b4bb2fdbbdd88f719c624a (
.fgallag_sel( I91812179d44cb675b90d477f33ec48ad[fgallag_SEL-1:0]),
.fgallag( Ic385923d90d69cd387eb9fb5f62fd9ba ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic420c6e4d3748dafd05197706f316f62 = (I91812179d44cb675b90d477f33ec48ad[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic385923d90d69cd387eb9fb5f62fd9ba ;

Ic9c2f173881d25f8976d723957809f51 If35314531f646278f5b327c89debd4ad (
.fgallag_sel( Idb04a1aae91fdc477ca38ed66789ee88[fgallag_SEL-1:0]),
.fgallag( I2f642acd0cb0bd30177bc0d65751ed99 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifd760e2ecefe198d6f583146e8cbe9fc = (Idb04a1aae91fdc477ca38ed66789ee88[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2f642acd0cb0bd30177bc0d65751ed99 ;

Ic9c2f173881d25f8976d723957809f51 I4c2171381c32c243ec85b2cbbc5f67cb (
.fgallag_sel( I566054aece562960590ee28b157e4a3e[fgallag_SEL-1:0]),
.fgallag( If1064670adff5b00cbf7809e2621cfd5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8078293bd2540592bffc91383fa5ad38 = (I566054aece562960590ee28b157e4a3e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If1064670adff5b00cbf7809e2621cfd5 ;

Ic9c2f173881d25f8976d723957809f51 Iee5286d12d53728f3ef52fd64632a80f (
.fgallag_sel( I7b2ffb762cd9ef7aa8ba224efb75c46c[fgallag_SEL-1:0]),
.fgallag( I72311a2c7557be2b6cb95b3bc6f511a5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1c0777b46bd3a7e2126f614d55703204 = (I7b2ffb762cd9ef7aa8ba224efb75c46c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I72311a2c7557be2b6cb95b3bc6f511a5 ;

Ic9c2f173881d25f8976d723957809f51 Ic3a697526d0421a6a24ae95ecba110da (
.fgallag_sel( Id90bbb642b0f4434d8a148a28b6b2f65[fgallag_SEL-1:0]),
.fgallag( I79ee4c7277f713aa710ae8cf7c470aa1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2a719cff60bf0985e451a32aa71c82fe = (Id90bbb642b0f4434d8a148a28b6b2f65[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I79ee4c7277f713aa710ae8cf7c470aa1 ;

Ic9c2f173881d25f8976d723957809f51 I9c7a05690c17ecbe726c08745c5d8611 (
.fgallag_sel( Ia4e297e35d484b15adce7e1d67f582b0[fgallag_SEL-1:0]),
.fgallag( I32bfef7a7ecaa533e3bf92fb560e657b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia1af17b99a087b22fecb7ff79a370363 = (Ia4e297e35d484b15adce7e1d67f582b0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I32bfef7a7ecaa533e3bf92fb560e657b ;

Ic9c2f173881d25f8976d723957809f51 Ibc0a202042a593794957c79a9ee8fb2f (
.fgallag_sel( I84996b1d03b692f6f736fb04c7f91e83[fgallag_SEL-1:0]),
.fgallag( If4a6b6a8b44d2c55c93b111d20525ec6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id75247b073a7993bff1992cfe1874ff6 = (I84996b1d03b692f6f736fb04c7f91e83[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If4a6b6a8b44d2c55c93b111d20525ec6 ;

Ic9c2f173881d25f8976d723957809f51 Ib7145e3b0c3fdd57349d77ca37425df5 (
.fgallag_sel( I83078cc7857fc17b30f640854a4d6be5[fgallag_SEL-1:0]),
.fgallag( I7d41f27ff64d549b7e5df6b172969d8a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I63a6ad22f067ea29cf79e51ebc011f8d = (I83078cc7857fc17b30f640854a4d6be5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7d41f27ff64d549b7e5df6b172969d8a ;

Ic9c2f173881d25f8976d723957809f51 I0b0895d7d86b2f3d0f4d7a9fdb53e110 (
.fgallag_sel( I94bb467129904032736fb13dd636c600[fgallag_SEL-1:0]),
.fgallag( Ie3a2d4d85d4e4ac011887cbd329bd9b7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic3b5918c230369180edc94c5b01046e7 = (I94bb467129904032736fb13dd636c600[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie3a2d4d85d4e4ac011887cbd329bd9b7 ;

Ic9c2f173881d25f8976d723957809f51 I10553709e5053d2974d3a13b14a05f1f (
.fgallag_sel( Ifa76758b50f439170ecd6d86ff898bc4[fgallag_SEL-1:0]),
.fgallag( I3bc9fcec69ab6a1efb2d86e03804415c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifdf2c8ac7eb668b49ed3cf950d08c179 = (Ifa76758b50f439170ecd6d86ff898bc4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3bc9fcec69ab6a1efb2d86e03804415c ;

Ic9c2f173881d25f8976d723957809f51 I4a42c4ddcd3ea434cbce7c5cc1249af0 (
.fgallag_sel( I9d831dd976e8cd5d8f6a6818601e6424[fgallag_SEL-1:0]),
.fgallag( I9ee16e46a399d1445fcdf251757a5e43 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I644ff86dfecc5a20a1431f9cc67ee6f9 = (I9d831dd976e8cd5d8f6a6818601e6424[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9ee16e46a399d1445fcdf251757a5e43 ;

Ic9c2f173881d25f8976d723957809f51 Idc009094d22e5e31bdb1dd2daf616475 (
.fgallag_sel( I474774ae149804412ed4aaf1cdcaba88[fgallag_SEL-1:0]),
.fgallag( I45cf986a60a429a68051f76beb8188fb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I56a7bd438035251cd67dfb97b3a345d7 = (I474774ae149804412ed4aaf1cdcaba88[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I45cf986a60a429a68051f76beb8188fb ;

Ic9c2f173881d25f8976d723957809f51 Ibd31a1c0943170d3b4c37b18e5fe18ff (
.fgallag_sel( I964cdcb4e6b49a62d30c2a2540851317[fgallag_SEL-1:0]),
.fgallag( I4e48461fcd58a133a09d856852887a4f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I00c294596fc87af7f1b8377260232832 = (I964cdcb4e6b49a62d30c2a2540851317[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4e48461fcd58a133a09d856852887a4f ;

Ic9c2f173881d25f8976d723957809f51 I9f272d1007b196c58847fbcbfe88e6eb (
.fgallag_sel( I6df268bc9f85ce88674a9165664ea84a[fgallag_SEL-1:0]),
.fgallag( I901714025da5b89ee929ea2859f3e6c7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7af09468b60d8e594a1aa85ad74911d5 = (I6df268bc9f85ce88674a9165664ea84a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I901714025da5b89ee929ea2859f3e6c7 ;

Ic9c2f173881d25f8976d723957809f51 I1da0acdc523e7e4d559b501a09c98ee8 (
.fgallag_sel( I74fdcbe9f49f7bce1f5e31d956c5883c[fgallag_SEL-1:0]),
.fgallag( I976786b0539b07b056dad0f050eeb53f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic0ed40d42c2af78809ecb381660ef229 = (I74fdcbe9f49f7bce1f5e31d956c5883c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I976786b0539b07b056dad0f050eeb53f ;

Ic9c2f173881d25f8976d723957809f51 I96f508156d3ec21b9e796e184a8d01eb (
.fgallag_sel( I4a1b8453cb7a21745d5f74ad05653ed2[fgallag_SEL-1:0]),
.fgallag( I8e1ad4f44dcac3e770dd862413b25a4e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie03547bf9963c8a716e20e4aaef52dc7 = (I4a1b8453cb7a21745d5f74ad05653ed2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8e1ad4f44dcac3e770dd862413b25a4e ;

Ic9c2f173881d25f8976d723957809f51 I0dec86884a25e6644cb2e16860ae3f21 (
.fgallag_sel( I9c53b478b2011fac0615a152fe60d5b6[fgallag_SEL-1:0]),
.fgallag( Iaf5caa6558f0a98b91fb72db734bbec4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I26e996666f3436cfa998f34c3a05f7db = (I9c53b478b2011fac0615a152fe60d5b6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaf5caa6558f0a98b91fb72db734bbec4 ;

Ic9c2f173881d25f8976d723957809f51 Ic5b91e2b7037f76980bfdf7dff9f87e5 (
.fgallag_sel( Id75dbed8f1a5befda32c60b994681013[fgallag_SEL-1:0]),
.fgallag( I7b37d3b1b23f09c6ac46a94cf2c4ead7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idfc51f66e038c5ae625e98b615a7beaf = (Id75dbed8f1a5befda32c60b994681013[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7b37d3b1b23f09c6ac46a94cf2c4ead7 ;

Ic9c2f173881d25f8976d723957809f51 Ide56a1f91d8ee71366c2bc03c12a56a4 (
.fgallag_sel( I378a59323b74623c5524f854d6e11226[fgallag_SEL-1:0]),
.fgallag( Ief8b577d924f257ae5e1dd47009b0db2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idedf5a83a99278f57c6c9294b66b69eb = (I378a59323b74623c5524f854d6e11226[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ief8b577d924f257ae5e1dd47009b0db2 ;

Ic9c2f173881d25f8976d723957809f51 If618188514cc03de8e0cbc2e4ef78b03 (
.fgallag_sel( I080bf885464a0cc948a4450e9f7d1d26[fgallag_SEL-1:0]),
.fgallag( Ie59366fcd6132a48f3e9be1bb5b600c6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idf55d61336e413c5aa3226b3b44f27b1 = (I080bf885464a0cc948a4450e9f7d1d26[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie59366fcd6132a48f3e9be1bb5b600c6 ;

Ic9c2f173881d25f8976d723957809f51 Iec240c8670b0c2629c81fbad884f22f5 (
.fgallag_sel( If769e73adea227de1fd85c2e89d0ba08[fgallag_SEL-1:0]),
.fgallag( I273c1e28c3ed897b7d0f6b36a3a8def9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I05ce5256e568621df7129058c50e9fa6 = (If769e73adea227de1fd85c2e89d0ba08[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I273c1e28c3ed897b7d0f6b36a3a8def9 ;

Ic9c2f173881d25f8976d723957809f51 I1986a21f85b8f91030e2d6f6abff6af9 (
.fgallag_sel( Ifa6a34b83225e9d9b28b14874c4444e3[fgallag_SEL-1:0]),
.fgallag( I64b507fe58b933919d0766631985a74e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib8af108fab1636823714995f78c9d575 = (Ifa6a34b83225e9d9b28b14874c4444e3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I64b507fe58b933919d0766631985a74e ;

Ic9c2f173881d25f8976d723957809f51 Ice0ccb2d9bed9e6410714a82e945fe00 (
.fgallag_sel( I584b1d4d6fb7ee4f20ad9c96715cdf90[fgallag_SEL-1:0]),
.fgallag( I7c0376cbc3660f3d82a5da22806ef5e3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I166d54ee9aa9002c59a0aca2834632f5 = (I584b1d4d6fb7ee4f20ad9c96715cdf90[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7c0376cbc3660f3d82a5da22806ef5e3 ;

Ic9c2f173881d25f8976d723957809f51 I08f5291d3ff10a6adcb69622649b8382 (
.fgallag_sel( I265f9b91fbb62164e589dcf96818c4f5[fgallag_SEL-1:0]),
.fgallag( I3884d561185660e7e0f461b3487fdfd4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib5f971498046dd212d853ff440c553cc = (I265f9b91fbb62164e589dcf96818c4f5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3884d561185660e7e0f461b3487fdfd4 ;

Ic9c2f173881d25f8976d723957809f51 I7dccba215dc4c89caab0711114e4b3a9 (
.fgallag_sel( I3d59a47c88227734cf6fc0d6fd30db11[fgallag_SEL-1:0]),
.fgallag( I4b991f90354e3f74d105a64929a97d6f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I325d401c6a1f445dcb7a83d90d2da75e = (I3d59a47c88227734cf6fc0d6fd30db11[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4b991f90354e3f74d105a64929a97d6f ;

Ic9c2f173881d25f8976d723957809f51 Ic9d3fb480964eb59d66825df481b00bb (
.fgallag_sel( I6144b6df2c87ea0948d730343b42129f[fgallag_SEL-1:0]),
.fgallag( I9534939768f7d2532ca4e6757dfafb72 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I91eeb6252974a1f69908b7e7114b95f5 = (I6144b6df2c87ea0948d730343b42129f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9534939768f7d2532ca4e6757dfafb72 ;

Ic9c2f173881d25f8976d723957809f51 Ia51c5f316d41e78125525b5f415839d9 (
.fgallag_sel( Ia7ca7400e36ea572fba8e19bcc81ecbd[fgallag_SEL-1:0]),
.fgallag( I090228a60e5919fa88d842b1638ee296 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I898cf70b6c6b57d256490f44d257fd84 = (Ia7ca7400e36ea572fba8e19bcc81ecbd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I090228a60e5919fa88d842b1638ee296 ;

Ic9c2f173881d25f8976d723957809f51 Iccce0d7f9085d642adace115425588d4 (
.fgallag_sel( I302e61b49accf5db556b87517f2341f5[fgallag_SEL-1:0]),
.fgallag( I8994d511d611a3c1b7a8122cd3d2825e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I256f73600515ae5c410454c425b66696 = (I302e61b49accf5db556b87517f2341f5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8994d511d611a3c1b7a8122cd3d2825e ;

Ic9c2f173881d25f8976d723957809f51 I2bdfdfa3ef47aa1694a8a90b2c262b73 (
.fgallag_sel( I5d9af1abff6efe3a55c6568d936b6ec7[fgallag_SEL-1:0]),
.fgallag( I43d14ec8853bfd211aa6b887c7ebdd5a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I362d1818937fd8d777531b85e86b4145 = (I5d9af1abff6efe3a55c6568d936b6ec7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I43d14ec8853bfd211aa6b887c7ebdd5a ;

Ic9c2f173881d25f8976d723957809f51 I71602677970470ed0886e5296fb6738e (
.fgallag_sel( I8cde0aa611c476b5112edeb8f17f15bf[fgallag_SEL-1:0]),
.fgallag( Icd810cceba64ffbb087600155338911c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I21dda2280e7aa79b6abd7820829583e1 = (I8cde0aa611c476b5112edeb8f17f15bf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Icd810cceba64ffbb087600155338911c ;

Ic9c2f173881d25f8976d723957809f51 If8fc6740480a1a2c27e624016c44ba86 (
.fgallag_sel( Icaa40ec40d6d26cdf70bb5ae7d492e47[fgallag_SEL-1:0]),
.fgallag( I33ddd4cdef0a0704f204f4fdb14fd859 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I94a6499c7bd1d40e4f363a58db1aa114 = (Icaa40ec40d6d26cdf70bb5ae7d492e47[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I33ddd4cdef0a0704f204f4fdb14fd859 ;

Ic9c2f173881d25f8976d723957809f51 Ia6f3b203a8db05058dfa669cc713e0ed (
.fgallag_sel( I8346f15d822cacfeecbe5d75412cb53f[fgallag_SEL-1:0]),
.fgallag( I0c87f78f08ac77246d7b3b8604dfd700 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifb6f3d60109d87ffd54e72b3958c7e80 = (I8346f15d822cacfeecbe5d75412cb53f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0c87f78f08ac77246d7b3b8604dfd700 ;

Ic9c2f173881d25f8976d723957809f51 I0f9982dc85082ca9eb67b035886ff0df (
.fgallag_sel( I5ee364aab320ab40c0f65feda6f53b18[fgallag_SEL-1:0]),
.fgallag( I54745c58c61eba829e4717cd842d519d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia3fca25225f6cd049ec92b44cdb57049 = (I5ee364aab320ab40c0f65feda6f53b18[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I54745c58c61eba829e4717cd842d519d ;

Ic9c2f173881d25f8976d723957809f51 I2c9948a993cc075d0b695750c6033bbb (
.fgallag_sel( I1f0ecba054900f96cd7100741191c5f4[fgallag_SEL-1:0]),
.fgallag( I9e278d7b6cccaa39163d0867427709ed ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iefa9788b8791b23ea0ca3d756d7e4019 = (I1f0ecba054900f96cd7100741191c5f4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9e278d7b6cccaa39163d0867427709ed ;

Ic9c2f173881d25f8976d723957809f51 I1fa5a07fde17cf8ad445bd8c3a7f45ba (
.fgallag_sel( I4faf2caf62966416118a54015908c889[fgallag_SEL-1:0]),
.fgallag( I3e5d8af6fed6b47aebf2eef7010afa8b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2b790f210029547ce774150b5390eb12 = (I4faf2caf62966416118a54015908c889[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3e5d8af6fed6b47aebf2eef7010afa8b ;

Ic9c2f173881d25f8976d723957809f51 Iccf07866aa6c7c266464f3b72ee72fcc (
.fgallag_sel( Idd0329980a36f87859150530ab44b52d[fgallag_SEL-1:0]),
.fgallag( Ie96538fd32c8f8d7a3144012d10b29a5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5c474a60ee2779b8f1477d07f4ca88d1 = (Idd0329980a36f87859150530ab44b52d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie96538fd32c8f8d7a3144012d10b29a5 ;

Ic9c2f173881d25f8976d723957809f51 I1ca6e00c5f6a111fcaf071628d0ac6d9 (
.fgallag_sel( Ie66bc10dde27f08813d4d347fd7cf6ce[fgallag_SEL-1:0]),
.fgallag( I050a226112c903de442358e2d5be8274 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie542464c6c79a43b078a8314c4def3b6 = (Ie66bc10dde27f08813d4d347fd7cf6ce[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I050a226112c903de442358e2d5be8274 ;

Ic9c2f173881d25f8976d723957809f51 I524f2621f8c0ea24dc195e5c586bb5ab (
.fgallag_sel( Ie1d8b3ea7c6603cebf2f9adb776910b7[fgallag_SEL-1:0]),
.fgallag( I4df410c6a7eea67fd73cc33c791e7aa0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0ae4560405030e9485f14f6eca025625 = (Ie1d8b3ea7c6603cebf2f9adb776910b7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4df410c6a7eea67fd73cc33c791e7aa0 ;

Ic9c2f173881d25f8976d723957809f51 I66030ce1b7c5d2bc3b06979194c99bd2 (
.fgallag_sel( Ia37488e9a50cf5cc08de74ade676db96[fgallag_SEL-1:0]),
.fgallag( Id7e318f124e0534c8e0538f99616ed01 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic14dfb6df2b9a62e5c9471684c0cb07f = (Ia37488e9a50cf5cc08de74ade676db96[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id7e318f124e0534c8e0538f99616ed01 ;

Ic9c2f173881d25f8976d723957809f51 I46bc851291db247c4259decfb7234484 (
.fgallag_sel( I08aa45211cab01d567cd5eb172fd2f0c[fgallag_SEL-1:0]),
.fgallag( I66ba7e48a07f5fdfe16d23b0dc243514 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia744719b1036a2236173a80ce326bb7d = (I08aa45211cab01d567cd5eb172fd2f0c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I66ba7e48a07f5fdfe16d23b0dc243514 ;

Ic9c2f173881d25f8976d723957809f51 I561255fa79e05d817e386ebe4e043d44 (
.fgallag_sel( If4ff0c63ec1deb46412858e496451a01[fgallag_SEL-1:0]),
.fgallag( I62e6e8be411f12cd5c4d63f1825521f3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic3f0e0640b27dd1a3bd39f6b9507c7fe = (If4ff0c63ec1deb46412858e496451a01[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I62e6e8be411f12cd5c4d63f1825521f3 ;

Ic9c2f173881d25f8976d723957809f51 Icdb8b0869a3ce682ad2680465f8695c1 (
.fgallag_sel( Ife7bfd15fc4c392b5d2288d9a4e879b3[fgallag_SEL-1:0]),
.fgallag( I2f94d5aad80c081124e3efa3804af183 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I82fa0db281b140ed781dcf5c53625117 = (Ife7bfd15fc4c392b5d2288d9a4e879b3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2f94d5aad80c081124e3efa3804af183 ;

Ic9c2f173881d25f8976d723957809f51 I00624bef8433ebf32bbd08743e7187e5 (
.fgallag_sel( I24ac26debafd03c7333d174e8725afd6[fgallag_SEL-1:0]),
.fgallag( I7a91b23716bf81bea4956eafb467c96a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5dfa454e544e731a6254e73c97d79e06 = (I24ac26debafd03c7333d174e8725afd6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7a91b23716bf81bea4956eafb467c96a ;

Ic9c2f173881d25f8976d723957809f51 I8c6c53466fc7de071f4c0fd02dbd4ff7 (
.fgallag_sel( I99d80ad68e2563d0f78a0e3bb82c5328[fgallag_SEL-1:0]),
.fgallag( I17572136bb435e84505c016523a6ec88 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3a57ff68cdc9b93c07bc79f8cea77473 = (I99d80ad68e2563d0f78a0e3bb82c5328[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I17572136bb435e84505c016523a6ec88 ;

Ic9c2f173881d25f8976d723957809f51 I89202989e60389422fb0a22d1f054d41 (
.fgallag_sel( I9943733ef305983c629565c881054bbf[fgallag_SEL-1:0]),
.fgallag( I9b0ac56afa21022e8bc69f5d20d17b66 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2f363d2944c634905ef5ec14c9cedf52 = (I9943733ef305983c629565c881054bbf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9b0ac56afa21022e8bc69f5d20d17b66 ;

Ic9c2f173881d25f8976d723957809f51 Ie35bcd6320f45ba64ea820c450920a57 (
.fgallag_sel( I7cb4420bc55c03a6500f5228d31fe43c[fgallag_SEL-1:0]),
.fgallag( Id9468cba18d4c67a84cb2b16d2cf495e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id15ed601c43171647305818c6f30ace5 = (I7cb4420bc55c03a6500f5228d31fe43c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id9468cba18d4c67a84cb2b16d2cf495e ;

Ic9c2f173881d25f8976d723957809f51 Ib305e5243db3c2c59808dc263c0a61f4 (
.fgallag_sel( Ic4d19dec464359c0a9fa75148fe90c73[fgallag_SEL-1:0]),
.fgallag( I2bda0265c40a5cedc359dee75fb15b4c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I75bed085cf80c0672fb41df1d6fc4545 = (Ic4d19dec464359c0a9fa75148fe90c73[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2bda0265c40a5cedc359dee75fb15b4c ;

Ic9c2f173881d25f8976d723957809f51 I4eff3bf39b3c3b08692cbde60e16c227 (
.fgallag_sel( I44993416e1d22613dbd78402c37a934d[fgallag_SEL-1:0]),
.fgallag( I318ebdf91ab8e83b80a880395879fc77 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib7f95eeae4f4565133ae98a0538e56c3 = (I44993416e1d22613dbd78402c37a934d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I318ebdf91ab8e83b80a880395879fc77 ;

Ic9c2f173881d25f8976d723957809f51 I72499f0beafbc997de05a24a7ca88d18 (
.fgallag_sel( Ibc9b94a9dea471805cb442ac6904bc97[fgallag_SEL-1:0]),
.fgallag( I8ac8dbc25a20c0c27e09240a5cd1bfd2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5a7c45c0b4ce4206080f2b50cb0a169f = (Ibc9b94a9dea471805cb442ac6904bc97[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8ac8dbc25a20c0c27e09240a5cd1bfd2 ;

Ic9c2f173881d25f8976d723957809f51 I7543e09c423bb7b6e59e4dc911b46490 (
.fgallag_sel( I917d9f9b144d3bffafc77bddae7fba6b[fgallag_SEL-1:0]),
.fgallag( Id8c4e5d6318622bd8ec2974684f542b6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I27cba499cffd339eddcdb4e2c846ee69 = (I917d9f9b144d3bffafc77bddae7fba6b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id8c4e5d6318622bd8ec2974684f542b6 ;

Ic9c2f173881d25f8976d723957809f51 Iccd2411b4a46915e8909fabc724e0b73 (
.fgallag_sel( Ibc91c6c3d56bb8a14e22909c43ffec51[fgallag_SEL-1:0]),
.fgallag( I8df19e0871c18890419c593410596b59 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifafce4fed1394ac5fa8849145960f2b5 = (Ibc91c6c3d56bb8a14e22909c43ffec51[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8df19e0871c18890419c593410596b59 ;

Ic9c2f173881d25f8976d723957809f51 Icdf677f62d44cf55263e2c5554bfb620 (
.fgallag_sel( If7c2d3eddd96b47b6c2aea8b27c8c7f4[fgallag_SEL-1:0]),
.fgallag( Ifb977d4c5bac50b9d7f2f814a500f0f2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1d6de59e71e329f79055285b3a50c2b4 = (If7c2d3eddd96b47b6c2aea8b27c8c7f4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifb977d4c5bac50b9d7f2f814a500f0f2 ;

Ic9c2f173881d25f8976d723957809f51 Ia2ebe09ffca58a7fd6f23bcfe29f94cb (
.fgallag_sel( I4df093ed94d26b058e97db550e347e3c[fgallag_SEL-1:0]),
.fgallag( Id9a1f5bd846dc7d093ed9392722317be ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9265fbbb34a66f13193ea1220ecb0589 = (I4df093ed94d26b058e97db550e347e3c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id9a1f5bd846dc7d093ed9392722317be ;

Ic9c2f173881d25f8976d723957809f51 I2ec614edfd0e3053872fd21859e74d57 (
.fgallag_sel( Ie90303b0326bee4ab203a8cf1e643da9[fgallag_SEL-1:0]),
.fgallag( Ic886ecf946cd5c297012444cb34980ab ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifcc01d5d37df8c68972086c44575e8d6 = (Ie90303b0326bee4ab203a8cf1e643da9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic886ecf946cd5c297012444cb34980ab ;

Ic9c2f173881d25f8976d723957809f51 If1125f76f5373be58c5eb978f3ce270e (
.fgallag_sel( I19030d352fd059156ee42c66f9270beb[fgallag_SEL-1:0]),
.fgallag( I37085a233f195dce1a76d05b0157fcac ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I57c25f5b2fecd18092653842e49e8d11 = (I19030d352fd059156ee42c66f9270beb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I37085a233f195dce1a76d05b0157fcac ;

Ic9c2f173881d25f8976d723957809f51 Ifa6560f13b8190ecf16994ebed29b9b1 (
.fgallag_sel( I36767a902c53a384128ae1443cf88963[fgallag_SEL-1:0]),
.fgallag( Ia2812d1ba8ca6831a2f059eb23384b38 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4b70004412f2ef37ac00fc19592b1f30 = (I36767a902c53a384128ae1443cf88963[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia2812d1ba8ca6831a2f059eb23384b38 ;

Ic9c2f173881d25f8976d723957809f51 I22fc3f82c4bda5fffa1c7615782288a1 (
.fgallag_sel( I868dffa3f07407f7996bb5bc596939b7[fgallag_SEL-1:0]),
.fgallag( Id176f2681568337762559e78cde29ba6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib952f8ef85514b1832324867adc72ce0 = (I868dffa3f07407f7996bb5bc596939b7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id176f2681568337762559e78cde29ba6 ;

Ic9c2f173881d25f8976d723957809f51 I5647a63be5649f1ec1f4ce44cb6aa177 (
.fgallag_sel( I7d928be164d0dce8b1322ff230c053e9[fgallag_SEL-1:0]),
.fgallag( Ia0c4e9942a4b08f69c2a027a712c9e39 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I08494381ebeda641f05b917fa31910a8 = (I7d928be164d0dce8b1322ff230c053e9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia0c4e9942a4b08f69c2a027a712c9e39 ;

Ic9c2f173881d25f8976d723957809f51 I24cccd71b9fc7f505ccb3e9caa249f7a (
.fgallag_sel( I98be4971a8a9a08abb3ebe474d7f0c6d[fgallag_SEL-1:0]),
.fgallag( I2da299005fed6f2b710e25acd48ebe91 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3f0568074c465ac281150bb70bbd76ec = (I98be4971a8a9a08abb3ebe474d7f0c6d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2da299005fed6f2b710e25acd48ebe91 ;

Ic9c2f173881d25f8976d723957809f51 I99a9fac6551fa4e7b0a0266eeb103062 (
.fgallag_sel( I779e70dea33201e9237f29681ffd5e27[fgallag_SEL-1:0]),
.fgallag( Ia1038e3b807e16a30f6f4564509ddd30 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib6b79505990d6499127f78e3186cc2a8 = (I779e70dea33201e9237f29681ffd5e27[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia1038e3b807e16a30f6f4564509ddd30 ;

Ic9c2f173881d25f8976d723957809f51 I945ffb47460675a3ee6a01a66b65e34c (
.fgallag_sel( Ie2262914042172ab7e08599278f36af5[fgallag_SEL-1:0]),
.fgallag( I25d94516522c19c0e53b5f52f4480216 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5404c19d5b4c44dddcca70138fbe79de = (Ie2262914042172ab7e08599278f36af5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I25d94516522c19c0e53b5f52f4480216 ;

Ic9c2f173881d25f8976d723957809f51 Ibff09d656542ae107d7ec4ddf86f4158 (
.fgallag_sel( I4001323da8f7956cdd480ac2d56df929[fgallag_SEL-1:0]),
.fgallag( I4b96be53e3d059113bb74b27ffe30179 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7265ecc942bf501ad034704f517d4e8d = (I4001323da8f7956cdd480ac2d56df929[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4b96be53e3d059113bb74b27ffe30179 ;

Ic9c2f173881d25f8976d723957809f51 I141551a66f1b8c9b3f04ca72803b31dc (
.fgallag_sel( Ib1cd6731034887a0a55e405c9db3e8de[fgallag_SEL-1:0]),
.fgallag( Ic091d8daff9f609c53cb191ed6b6ddeb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1c114e8dfd37b1d182028679b3974a1b = (Ib1cd6731034887a0a55e405c9db3e8de[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic091d8daff9f609c53cb191ed6b6ddeb ;

Ic9c2f173881d25f8976d723957809f51 I2810971df22b92df23514fa2fa03afd4 (
.fgallag_sel( I51aa496e8c03944c28a908102514e6f8[fgallag_SEL-1:0]),
.fgallag( I2468caeaf9733c8bc6a485542b6b263f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9fa799fd606c85184ce84138a90f03e1 = (I51aa496e8c03944c28a908102514e6f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2468caeaf9733c8bc6a485542b6b263f ;

Ic9c2f173881d25f8976d723957809f51 Ic9867e497014c45ab4b33ef05eaf5534 (
.fgallag_sel( I6415f3996318472532e161510ccc8ca3[fgallag_SEL-1:0]),
.fgallag( I6611d1fa58dd253fe6344a41584d7e22 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id8b3ba6e7ffd04674b2ae10b928f26f0 = (I6415f3996318472532e161510ccc8ca3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6611d1fa58dd253fe6344a41584d7e22 ;

Ic9c2f173881d25f8976d723957809f51 Ibeac37239c6549d44f5614d459ad2a5c (
.fgallag_sel( Ia11b671b59240988737979328c472812[fgallag_SEL-1:0]),
.fgallag( I8afb33eced17e8675a8e2bd90d16030b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id4cc4e9883ae7b27bed350ba292d9349 = (Ia11b671b59240988737979328c472812[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8afb33eced17e8675a8e2bd90d16030b ;

Ic9c2f173881d25f8976d723957809f51 I9ec0aa74cc34a9090bbce22e28502dfd (
.fgallag_sel( Id4fabe0165a117a402dc14f2f3ec626a[fgallag_SEL-1:0]),
.fgallag( Idac55755226133905d3250273b1eccb8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5c3099cb6fc046e62863a69945ae3e04 = (Id4fabe0165a117a402dc14f2f3ec626a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idac55755226133905d3250273b1eccb8 ;

Ic9c2f173881d25f8976d723957809f51 Ic2152f424753e4aa2ea051ff9d6121bb (
.fgallag_sel( I57238f501ab7278b308d76211ced8cf7[fgallag_SEL-1:0]),
.fgallag( I4cd564459b8d65976195b2994e7d44f2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If48b274e1e1809931eb2be69a565a443 = (I57238f501ab7278b308d76211ced8cf7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4cd564459b8d65976195b2994e7d44f2 ;

Ic9c2f173881d25f8976d723957809f51 Ica6370f606cf528e491ebf370aa5ea49 (
.fgallag_sel( I9b257f8556ca4e5402637f01081b78e1[fgallag_SEL-1:0]),
.fgallag( I2280162ee1c08ccc9f0c17d1ca0e3628 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1667cbf3caf9a10527531b6aa69df847 = (I9b257f8556ca4e5402637f01081b78e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2280162ee1c08ccc9f0c17d1ca0e3628 ;

Ic9c2f173881d25f8976d723957809f51 I740c13219d137b936824f7cc7538a973 (
.fgallag_sel( I2e093412a9fa3972cea01664389d8c27[fgallag_SEL-1:0]),
.fgallag( I28b3ba64175358f277427fd790a9228b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I80ddcee29ed7af07148977eddab4bccd = (I2e093412a9fa3972cea01664389d8c27[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I28b3ba64175358f277427fd790a9228b ;

Ic9c2f173881d25f8976d723957809f51 Ia005d9743c601eb3653c6b092400bacc (
.fgallag_sel( I17907fd8c6975c8c642535ff929221a6[fgallag_SEL-1:0]),
.fgallag( I6c03138440f9bd0cb2cfe12abf619c10 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I32ab257af6a54e78706c6d83b579bcd6 = (I17907fd8c6975c8c642535ff929221a6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6c03138440f9bd0cb2cfe12abf619c10 ;

Ic9c2f173881d25f8976d723957809f51 I2a2b7b0432b44bae28ac48173f7b485a (
.fgallag_sel( I3c6577b04ad56d864bbaa2c048323c11[fgallag_SEL-1:0]),
.fgallag( Ib3709eb9dfc3a594d38ea5a0ef0cd444 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I907f4db1352049380285f358cac2b439 = (I3c6577b04ad56d864bbaa2c048323c11[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib3709eb9dfc3a594d38ea5a0ef0cd444 ;

Ic9c2f173881d25f8976d723957809f51 I518f47a19bc399a2420c647aff95f638 (
.fgallag_sel( I6f0c341c05eaa8f35bbce4521f6e8f94[fgallag_SEL-1:0]),
.fgallag( I44cf5ba18d7d029df13f446f09191b2c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I22cd5fb22f122d99e37e6c1ca2666301 = (I6f0c341c05eaa8f35bbce4521f6e8f94[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I44cf5ba18d7d029df13f446f09191b2c ;

Ic9c2f173881d25f8976d723957809f51 I38ca8a80bf2eb73aef3971fc6aeec316 (
.fgallag_sel( Ib72ba950ecf9ae2668374f6633a67ca7[fgallag_SEL-1:0]),
.fgallag( I6aa1e5acf0c2b01c94438bd1cff484c6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I892abe227878c5232de3ccd90e8c13e5 = (Ib72ba950ecf9ae2668374f6633a67ca7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6aa1e5acf0c2b01c94438bd1cff484c6 ;

Ic9c2f173881d25f8976d723957809f51 If4eae9d96138b09b1b3ba3c2968ea039 (
.fgallag_sel( I3d7c72d725f4563bb562e2992093cb02[fgallag_SEL-1:0]),
.fgallag( Ia23629f3881e4119c36576f7da58ceaa ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If5086f7447696a697be414fe50ad91fd = (I3d7c72d725f4563bb562e2992093cb02[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia23629f3881e4119c36576f7da58ceaa ;

Ic9c2f173881d25f8976d723957809f51 Ic5fced29c8c9b7e5f06b65fab1f16af0 (
.fgallag_sel( I813c881ac61a59041be3be78f6a466c8[fgallag_SEL-1:0]),
.fgallag( I2f12d1fa0b815564cefafc28ceb3de82 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9dc20c15b19d9351497997c81511c744 = (I813c881ac61a59041be3be78f6a466c8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2f12d1fa0b815564cefafc28ceb3de82 ;

Ic9c2f173881d25f8976d723957809f51 I3cb5722b97ecd4f57fa0a8fdf3e04b28 (
.fgallag_sel( I866510e7dc721fa5aac312bc5ab5ba0a[fgallag_SEL-1:0]),
.fgallag( Ib09ac099bcf61b09922b353403b29987 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I254c64de80d2a159aa0b3f3170042079 = (I866510e7dc721fa5aac312bc5ab5ba0a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib09ac099bcf61b09922b353403b29987 ;

Ic9c2f173881d25f8976d723957809f51 I20bfdcf809dc96ac5a46325031429066 (
.fgallag_sel( Ib4432359f97849dff6ad3e0f044157bd[fgallag_SEL-1:0]),
.fgallag( I3c2b6da8e286d0a7b628ba1071f29424 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4dae38e87f09d78c748974da00f274f8 = (Ib4432359f97849dff6ad3e0f044157bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3c2b6da8e286d0a7b628ba1071f29424 ;

Ic9c2f173881d25f8976d723957809f51 I9e99f67736c399017f0f71e2defb96ab (
.fgallag_sel( Ic86aa6eb1b4dcc2520309089b43292e6[fgallag_SEL-1:0]),
.fgallag( I550630b507ceec38b960ab2a86a57f1a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic8edf24599f1eee2af3576dfb2a6829a = (Ic86aa6eb1b4dcc2520309089b43292e6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I550630b507ceec38b960ab2a86a57f1a ;

Ic9c2f173881d25f8976d723957809f51 Ibfa7d030ba9a5dd5aa12a990175f3b1c (
.fgallag_sel( I0731115afe5c15bcf131f7ef4f05802b[fgallag_SEL-1:0]),
.fgallag( I795c1c91cb6b7870b7efb07d67085be1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I144ca4c629cc3134a991414038cfc9cf = (I0731115afe5c15bcf131f7ef4f05802b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I795c1c91cb6b7870b7efb07d67085be1 ;

Ic9c2f173881d25f8976d723957809f51 I0afa41900d31951d6b42c44b1e9759cb (
.fgallag_sel( Ib080b8fd34385aa7986dace4afd95267[fgallag_SEL-1:0]),
.fgallag( I531b70d12349f3bc67e6a3ec53368d97 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I379ed527c944420bb59be58b85ab4704 = (Ib080b8fd34385aa7986dace4afd95267[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I531b70d12349f3bc67e6a3ec53368d97 ;

Ic9c2f173881d25f8976d723957809f51 I32f32c938b26f4d567d9a4393a8ffbfe (
.fgallag_sel( I134890b77451d0b78afc7402a6a28048[fgallag_SEL-1:0]),
.fgallag( Id8a109043bc922b718c203bd5d60a999 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id37ddd7be0621f84793d1600ce915236 = (I134890b77451d0b78afc7402a6a28048[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id8a109043bc922b718c203bd5d60a999 ;

Ic9c2f173881d25f8976d723957809f51 I8182b58ba5cc359d93cf1f1568d2b9ad (
.fgallag_sel( I956da75f13433c1dd7a3cbd3b78922c1[fgallag_SEL-1:0]),
.fgallag( Ic126109499ee1dc2787ab05b404e7ae2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I20bbdbbee46a2be5c6caa56786345e8b = (I956da75f13433c1dd7a3cbd3b78922c1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic126109499ee1dc2787ab05b404e7ae2 ;

Ic9c2f173881d25f8976d723957809f51 I22d0d1a5ba4eb56b3a2af8a732dde64c (
.fgallag_sel( I440b26c9f1b9ccf70f97c9d5f732d38e[fgallag_SEL-1:0]),
.fgallag( I1cd8ba53b876e2436901749e355f354b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I02199c9dc39a2c8be49a1c96aa89de15 = (I440b26c9f1b9ccf70f97c9d5f732d38e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1cd8ba53b876e2436901749e355f354b ;

Ic9c2f173881d25f8976d723957809f51 Ie233e3a0a524d9df92af21058db6aa3e (
.fgallag_sel( I5e3a441faca44bffc4368d96d8fb0bfd[fgallag_SEL-1:0]),
.fgallag( I4e8ff51a6f70f8ca6a17a1dea8caf0a9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I17b1742efeadf5df716128d6603ebe99 = (I5e3a441faca44bffc4368d96d8fb0bfd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4e8ff51a6f70f8ca6a17a1dea8caf0a9 ;

Ic9c2f173881d25f8976d723957809f51 I31ad0e243f034e0b06c9f82860683341 (
.fgallag_sel( I21d7ba25247a87a1a9c245d0d1f553b0[fgallag_SEL-1:0]),
.fgallag( Ic1a27480c9acc1684f3fed116d74cb5f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I68da2c2a43373cf8145e6f7072bb5ca9 = (I21d7ba25247a87a1a9c245d0d1f553b0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic1a27480c9acc1684f3fed116d74cb5f ;

Ic9c2f173881d25f8976d723957809f51 I8d076b70cbf2db7913f0ad5f32d38c50 (
.fgallag_sel( I55aafa8162cfc4fccfae68cf78cd1c2b[fgallag_SEL-1:0]),
.fgallag( I0df7a888610865486aa1aaa2703dd041 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I27f3ef61a2ffbd4154a7b683aacd4844 = (I55aafa8162cfc4fccfae68cf78cd1c2b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0df7a888610865486aa1aaa2703dd041 ;

Ic9c2f173881d25f8976d723957809f51 Id9fe97a4843e48be6074128d5803436e (
.fgallag_sel( Ib99c25f0d8d6493cac4d5c816884c704[fgallag_SEL-1:0]),
.fgallag( If6448c72403a3d0bd904beac87f8aa96 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0726f4d2f2b1d495b1b439f998193435 = (Ib99c25f0d8d6493cac4d5c816884c704[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If6448c72403a3d0bd904beac87f8aa96 ;

Ic9c2f173881d25f8976d723957809f51 I02c20f5c3680c62e4baaf109879e5e34 (
.fgallag_sel( Iee7c9f0a0e8ca127efee008b4874edbd[fgallag_SEL-1:0]),
.fgallag( Iecf45496b391208d62e88544b5d2ca49 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I05e3c3e8567ed11012cf9f9d7ecb629a = (Iee7c9f0a0e8ca127efee008b4874edbd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iecf45496b391208d62e88544b5d2ca49 ;

Ic9c2f173881d25f8976d723957809f51 I8318346849d58d493b8d4723ac596692 (
.fgallag_sel( I17b4a3baae65161387f472037ffc6fc4[fgallag_SEL-1:0]),
.fgallag( Ib0fd0a839c85f3da5ae7b221f6e623d6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I210ade98fc479cdb069e2b028f1920d4 = (I17b4a3baae65161387f472037ffc6fc4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib0fd0a839c85f3da5ae7b221f6e623d6 ;

Ic9c2f173881d25f8976d723957809f51 Ib05f7f62fe4ab3221059b72198e1d569 (
.fgallag_sel( Ie7b7b202a968fe73f6b1e02a044414c5[fgallag_SEL-1:0]),
.fgallag( Ie045750c9289c899860823f90a306f3c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic89a704c9de69cff5b09d1b3bb220fe8 = (Ie7b7b202a968fe73f6b1e02a044414c5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie045750c9289c899860823f90a306f3c ;

Ic9c2f173881d25f8976d723957809f51 Id72885e0e75e2275156582e3126be1d1 (
.fgallag_sel( I479ab5c0e483c36267d8248340006666[fgallag_SEL-1:0]),
.fgallag( I1627b19e0ca42f9c264b626809fb37b7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic8ba8abf8a87610d08fb5a8174639f99 = (I479ab5c0e483c36267d8248340006666[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1627b19e0ca42f9c264b626809fb37b7 ;

Ic9c2f173881d25f8976d723957809f51 Ideb266655a1ec6b7bb94536f8d42cc8d (
.fgallag_sel( I777bfe165e25d7fde4fc950f23db7b84[fgallag_SEL-1:0]),
.fgallag( Ic9593f3fe23f258c2ab4ddcadaa8ca4c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9c0a1bb49be6604f75611b92d937c124 = (I777bfe165e25d7fde4fc950f23db7b84[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic9593f3fe23f258c2ab4ddcadaa8ca4c ;

Ic9c2f173881d25f8976d723957809f51 Id76d9386034980aa7086d38ceb827cf4 (
.fgallag_sel( I146d505a34ddb8d65e0a1769f623a7fd[fgallag_SEL-1:0]),
.fgallag( Idc0085a6595a7de7e2bc87c789b7d935 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iff70fe838ee16e8e35b1034135555acc = (I146d505a34ddb8d65e0a1769f623a7fd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idc0085a6595a7de7e2bc87c789b7d935 ;

Ic9c2f173881d25f8976d723957809f51 Ie08b9024aa7d1aa566173671f48bc6ab (
.fgallag_sel( Ia85239bddc04bf50bcf037ed2f76d7ac[fgallag_SEL-1:0]),
.fgallag( Id029b4c310acea870263d3715689e729 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibb4daaccffcf82b4cb4c431923c71f3f = (Ia85239bddc04bf50bcf037ed2f76d7ac[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id029b4c310acea870263d3715689e729 ;

Ic9c2f173881d25f8976d723957809f51 I526e69458c7eff77bc4451817cc57657 (
.fgallag_sel( Ia7306bacf3c2b180d3261a5c1f0f4a30[fgallag_SEL-1:0]),
.fgallag( Iec123ddb8d1e623d03d85a667c97ef31 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9c1fd2b57c1756bf67bc8cf5ed4a1912 = (Ia7306bacf3c2b180d3261a5c1f0f4a30[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iec123ddb8d1e623d03d85a667c97ef31 ;

Ic9c2f173881d25f8976d723957809f51 Ia0d4ae41c544627fb9766d80da5424a7 (
.fgallag_sel( I2018147b86e47af5842c4f29d047d157[fgallag_SEL-1:0]),
.fgallag( I89f0b0713e165a454e187fa51e89c642 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I71d437815bcfb755e16fc442431b6f68 = (I2018147b86e47af5842c4f29d047d157[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I89f0b0713e165a454e187fa51e89c642 ;

Ic9c2f173881d25f8976d723957809f51 I6ac3d38fc5fc63607a63c4c30b99e32c (
.fgallag_sel( Id17a85459845f8a8be694c4bf1fc29c9[fgallag_SEL-1:0]),
.fgallag( Id812cf3919ed50a5e3897d129eeb4b8d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4e3e1eb8ea6dfb08ea2634a9bab8319b = (Id17a85459845f8a8be694c4bf1fc29c9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id812cf3919ed50a5e3897d129eeb4b8d ;

Ic9c2f173881d25f8976d723957809f51 I306564b8b1e65d8a373ea722945acdf6 (
.fgallag_sel( Ic012b15584d9d25af38f83d0526503da[fgallag_SEL-1:0]),
.fgallag( I2d65b5115be2a22ed1e29426be3f0d15 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1fa2749e15c3bd7253a023eb01140cc7 = (Ic012b15584d9d25af38f83d0526503da[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2d65b5115be2a22ed1e29426be3f0d15 ;

Ic9c2f173881d25f8976d723957809f51 Icb614058c4c965e827bce2542b2285ef (
.fgallag_sel( I7f09bd4a45143a036ce04af11b9927f9[fgallag_SEL-1:0]),
.fgallag( I47c8671569e2c5c2a21f27aff2d1f4b8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie19e8502010d0c178f9f2da8df3fa63d = (I7f09bd4a45143a036ce04af11b9927f9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I47c8671569e2c5c2a21f27aff2d1f4b8 ;

Ic9c2f173881d25f8976d723957809f51 I1ff45c618d3a04edd62c7a6351300ec1 (
.fgallag_sel( Ica32f94af6e6f3eaf2b724a2173fa463[fgallag_SEL-1:0]),
.fgallag( Iaf2144dab2167cd2629067e40bea3053 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia512ada6f00f86ff495ae12ead6607d3 = (Ica32f94af6e6f3eaf2b724a2173fa463[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaf2144dab2167cd2629067e40bea3053 ;

Ic9c2f173881d25f8976d723957809f51 Iad1c0882ca7d98fc779c6982c5f588fd (
.fgallag_sel( Ib750bb83ddfbbad2a2be8d1c8392b4ff[fgallag_SEL-1:0]),
.fgallag( I4c2b80e4bbbd4c5e8d0da28c5d0f681e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If7b2398d3426250d73917539ff743c8a = (Ib750bb83ddfbbad2a2be8d1c8392b4ff[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4c2b80e4bbbd4c5e8d0da28c5d0f681e ;

Ic9c2f173881d25f8976d723957809f51 I9e99d12ae2805e75c8b4ff0627306bee (
.fgallag_sel( I3906ece39480f96020717c6243e8ba4c[fgallag_SEL-1:0]),
.fgallag( I6300fbbd385ad9280c751076bc68d70c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6446a839157f78880fc3fc7d8c378c78 = (I3906ece39480f96020717c6243e8ba4c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6300fbbd385ad9280c751076bc68d70c ;

Ic9c2f173881d25f8976d723957809f51 I82579bd8a2860f3e3c19c4306b285c62 (
.fgallag_sel( Ie68ce21ade07fa53c30ebf27216b03f9[fgallag_SEL-1:0]),
.fgallag( Iea078843b3c5139a395997c54462850a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I53504e8899a821cebe69ed590a3fd7fc = (Ie68ce21ade07fa53c30ebf27216b03f9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iea078843b3c5139a395997c54462850a ;

Ic9c2f173881d25f8976d723957809f51 Ie375b66e4d5059edf550c2c136461bbd (
.fgallag_sel( I6cc6fa167c0d2b4b62ddbeecea175ed2[fgallag_SEL-1:0]),
.fgallag( I654debf65019f2748e631a051f3b17ca ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If7d5fe39b147f24303884de3a30d669d = (I6cc6fa167c0d2b4b62ddbeecea175ed2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I654debf65019f2748e631a051f3b17ca ;

Ic9c2f173881d25f8976d723957809f51 I534dfe4fa3ed598e76b4a37591a02c89 (
.fgallag_sel( Ibddf3468ae7c27d5a4b1388e524aa9c2[fgallag_SEL-1:0]),
.fgallag( I1e88b57c19a1ddfc1c1f0e168b60f814 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I24c005d076b3c887d45d1285a4fe1bc5 = (Ibddf3468ae7c27d5a4b1388e524aa9c2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1e88b57c19a1ddfc1c1f0e168b60f814 ;

Ic9c2f173881d25f8976d723957809f51 Ic3a6d3d92f2849aa7be63e7124e564f8 (
.fgallag_sel( Iadcb2b3acaac2e1bb505c65d3cbe4235[fgallag_SEL-1:0]),
.fgallag( Ibaf7ab7333434b0d7e76e436ee40a406 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I18e00688f19c522b305d223ead684fb7 = (Iadcb2b3acaac2e1bb505c65d3cbe4235[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibaf7ab7333434b0d7e76e436ee40a406 ;

Ic9c2f173881d25f8976d723957809f51 Ife78eed3f26b5ddd17a091c65891ad27 (
.fgallag_sel( I37cd96b8b0a4939d9a70098fd8bcf452[fgallag_SEL-1:0]),
.fgallag( I1af14572832bd6d6b5890b8340b79ec7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0258ec63762460afb41bcd6e8869ec69 = (I37cd96b8b0a4939d9a70098fd8bcf452[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1af14572832bd6d6b5890b8340b79ec7 ;

Ic9c2f173881d25f8976d723957809f51 I378b470c0406630a49e2db2d2d1261a7 (
.fgallag_sel( Ib34b169dcc76daee2d1aa2b2a7513af3[fgallag_SEL-1:0]),
.fgallag( I652d3ed935b39f8fda8d84296456d633 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id1280129b20bd6389618695aec9efeed = (Ib34b169dcc76daee2d1aa2b2a7513af3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I652d3ed935b39f8fda8d84296456d633 ;

Ic9c2f173881d25f8976d723957809f51 Iccc5298adfb3a7a1dc1381154b29111d (
.fgallag_sel( If36fc316d6ec7c7e09eae77807b37099[fgallag_SEL-1:0]),
.fgallag( I5e33cad360aae934f418852541f5f2bd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I907fd3abdcadda1cd7149c7cf01e5751 = (If36fc316d6ec7c7e09eae77807b37099[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5e33cad360aae934f418852541f5f2bd ;

Ic9c2f173881d25f8976d723957809f51 I9f2a0d53e12f9225ac0b42d6444ec936 (
.fgallag_sel( Ifd214c332218ac5c0fe5aded4b952711[fgallag_SEL-1:0]),
.fgallag( If950e448e3cba7cc9aa7aff7718775f7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I73f044469c4dbcd5a98c0f83d6d043c4 = (Ifd214c332218ac5c0fe5aded4b952711[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If950e448e3cba7cc9aa7aff7718775f7 ;

Ic9c2f173881d25f8976d723957809f51 Ib270c26ef164be344d26ad66a2ed11dd (
.fgallag_sel( Idcd0fc8f86e2b6f03606b818b8346e5a[fgallag_SEL-1:0]),
.fgallag( I9adf8836419a1c85b146e5e36de68af5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2934a8783b90254606bcd933c629577f = (Idcd0fc8f86e2b6f03606b818b8346e5a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9adf8836419a1c85b146e5e36de68af5 ;

Ic9c2f173881d25f8976d723957809f51 Ib85b64da247f24dbae43b98c3af3d0a6 (
.fgallag_sel( If486aa8ac2cfb46f936714812cc760df[fgallag_SEL-1:0]),
.fgallag( I0f2bcdf124dff4219fd1a35ed1db7937 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id26b2a9c13424769e1627b1549159a7e = (If486aa8ac2cfb46f936714812cc760df[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0f2bcdf124dff4219fd1a35ed1db7937 ;

Ic9c2f173881d25f8976d723957809f51 I7e09ed0224f9736e7e62b78976ad026a (
.fgallag_sel( I2d8e5b5fdbda7d599423c38aaace6658[fgallag_SEL-1:0]),
.fgallag( Iae82e5de28b12f962bd7c5e221317ac2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2115e45deea528402794afadd17d9fe7 = (I2d8e5b5fdbda7d599423c38aaace6658[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iae82e5de28b12f962bd7c5e221317ac2 ;

Ic9c2f173881d25f8976d723957809f51 I3d1c29904f40ae7a959a632fad15257f (
.fgallag_sel( I6d0878fb7ec75c0a26be4dbba62f80dc[fgallag_SEL-1:0]),
.fgallag( Ia7b3cb9de8e18f41561c2a46dda8696a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I978020f8aaeb98cc1cea9360ec06da22 = (I6d0878fb7ec75c0a26be4dbba62f80dc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia7b3cb9de8e18f41561c2a46dda8696a ;

Ic9c2f173881d25f8976d723957809f51 I446fca9581378e7f0fedf6968b4d0776 (
.fgallag_sel( I16a16ff0e8a6685a09803634da429fd2[fgallag_SEL-1:0]),
.fgallag( Id0119672c8b017bce6fdba53d4dccf8b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icded30641e4770e30ee34bbf8d2a5721 = (I16a16ff0e8a6685a09803634da429fd2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id0119672c8b017bce6fdba53d4dccf8b ;

Ic9c2f173881d25f8976d723957809f51 I70165c87f1188ef18a62326c52b4590c (
.fgallag_sel( Idb211abaa54ac26e7379c64a63f7d07c[fgallag_SEL-1:0]),
.fgallag( I4aaef2f654ba03b1dc05719c81d5da69 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I02e3cbacce4e97e3088360f0acccee44 = (Idb211abaa54ac26e7379c64a63f7d07c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4aaef2f654ba03b1dc05719c81d5da69 ;

Ic9c2f173881d25f8976d723957809f51 Ia42b8bbe94d46d99af358f9ef4ab8516 (
.fgallag_sel( I351205eb71acb31b59d2b4470f0ba28c[fgallag_SEL-1:0]),
.fgallag( Ia6355e548635a4107a11c7952aa8b3d9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icbdf81888af42710561aec48ce84e3cb = (I351205eb71acb31b59d2b4470f0ba28c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia6355e548635a4107a11c7952aa8b3d9 ;

Ic9c2f173881d25f8976d723957809f51 Ibfa9b3c5fd70271b1ac615ecd37195c3 (
.fgallag_sel( If5660c495bf7690252783d888d1ad6e8[fgallag_SEL-1:0]),
.fgallag( I0bd950eee6abde9d1eaaabbe902fff5d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iea3ce04a4b8cc466e892aab886e63744 = (If5660c495bf7690252783d888d1ad6e8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0bd950eee6abde9d1eaaabbe902fff5d ;

Ic9c2f173881d25f8976d723957809f51 I33cb9d977791fd79db2890e62669c2e2 (
.fgallag_sel( I3a5229cb8e44a15560b5c7bef96e65cc[fgallag_SEL-1:0]),
.fgallag( I93caf487f67a2adce04a7b2cd7fff358 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3ca9464d884ccc7e2f396a74baea5bb9 = (I3a5229cb8e44a15560b5c7bef96e65cc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I93caf487f67a2adce04a7b2cd7fff358 ;

Ic9c2f173881d25f8976d723957809f51 I89c1f5b3ea8c41c0b55cff773f1d7df8 (
.fgallag_sel( I889b9b0828e97fe44d8366c5ef71a8f2[fgallag_SEL-1:0]),
.fgallag( If68a9cc5609ea7d87062bad2ebddb1a8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7b8d02aa08cde64a409f3766f940233c = (I889b9b0828e97fe44d8366c5ef71a8f2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If68a9cc5609ea7d87062bad2ebddb1a8 ;

Ic9c2f173881d25f8976d723957809f51 Iafa2fdf3f9d1c03f5e7003cb0ca1db29 (
.fgallag_sel( Ie23062e00e39ead706f5b6ead233747d[fgallag_SEL-1:0]),
.fgallag( If201a7afedfd1c329b55048e6bbad629 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I86ad427fe92cd4346b32ecf3c99c93c7 = (Ie23062e00e39ead706f5b6ead233747d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If201a7afedfd1c329b55048e6bbad629 ;

Ic9c2f173881d25f8976d723957809f51 I5fad54f1dbf719b0678522dafb06f695 (
.fgallag_sel( I8a2589544c75ecfdc31d28912c639695[fgallag_SEL-1:0]),
.fgallag( I1f8936599ead5ce1cd85132e382533f1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6667614b2fe12d6f63ac7737bf069b42 = (I8a2589544c75ecfdc31d28912c639695[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1f8936599ead5ce1cd85132e382533f1 ;

Ic9c2f173881d25f8976d723957809f51 I9f97bb7c91636a169ae44e096456b16f (
.fgallag_sel( I5c21c59147e9c3a74c7cbbb6f2a23919[fgallag_SEL-1:0]),
.fgallag( I37eb148270af62adba8341c83411f9f2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I909cbd582f015b4eabefd660b2039ccc = (I5c21c59147e9c3a74c7cbbb6f2a23919[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I37eb148270af62adba8341c83411f9f2 ;

Ic9c2f173881d25f8976d723957809f51 I39f0eeccfcc0cf5a0723e04bb90844ad (
.fgallag_sel( Idacd78e24408e432abbbfb0c447fdde5[fgallag_SEL-1:0]),
.fgallag( Ie4729048b95fede1806dbd006de01338 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie3433004b0ea3bba81f0b7502c69c821 = (Idacd78e24408e432abbbfb0c447fdde5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie4729048b95fede1806dbd006de01338 ;

Ic9c2f173881d25f8976d723957809f51 Ibf3028258671c7e2f825d8dc5daa69ed (
.fgallag_sel( I0e8b171fe5080485a7f4fef83f1f1528[fgallag_SEL-1:0]),
.fgallag( I02330d212434a6e8c303db2c3d36a3e5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If548fc27869a7e48fedc89bd5c8037f0 = (I0e8b171fe5080485a7f4fef83f1f1528[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I02330d212434a6e8c303db2c3d36a3e5 ;

Ic9c2f173881d25f8976d723957809f51 I6d370ac445a6f109441d51743bbdb8f0 (
.fgallag_sel( Ib22c2bd76e6c29cc2f1440885bf24b7b[fgallag_SEL-1:0]),
.fgallag( Id89498cf205e0cdef4886afd878c48f6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7cc21b5c21f6bc0603c3d57c86feeb00 = (Ib22c2bd76e6c29cc2f1440885bf24b7b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id89498cf205e0cdef4886afd878c48f6 ;

Ic9c2f173881d25f8976d723957809f51 I9d3521ed906da986e321765d554a4d35 (
.fgallag_sel( I149559fccd9def4ec1ead1fdcff3c7fd[fgallag_SEL-1:0]),
.fgallag( I547ae5055196f12eeeb36d69c325b84d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9ce2b40cd4433999690bb6e5c368e9b8 = (I149559fccd9def4ec1ead1fdcff3c7fd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I547ae5055196f12eeeb36d69c325b84d ;

Ic9c2f173881d25f8976d723957809f51 I2c3d4dd3b336fccec3a1143e69ed78a5 (
.fgallag_sel( Icfa8fed3239748abca27a5fc17de79c0[fgallag_SEL-1:0]),
.fgallag( I4871ccbe2f182791243b7bdcc9b8e286 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie102c1592ae8606ab75b1f7101b44918 = (Icfa8fed3239748abca27a5fc17de79c0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4871ccbe2f182791243b7bdcc9b8e286 ;

Ic9c2f173881d25f8976d723957809f51 I276d54ab3676216a75f18526621e872d (
.fgallag_sel( I2ff115fa483f080d93bada49a9566b33[fgallag_SEL-1:0]),
.fgallag( I12fd829f22ba908180290432320a3660 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I23ef94c5c29e674714d4ea1ad2d3f0e8 = (I2ff115fa483f080d93bada49a9566b33[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I12fd829f22ba908180290432320a3660 ;

Ic9c2f173881d25f8976d723957809f51 Ic16e68414dbff48be77bb1b20c7e2138 (
.fgallag_sel( Ibee4f3cd2f516c29ab68e07a640ab65e[fgallag_SEL-1:0]),
.fgallag( I8f967710d03870e026564db0df46d146 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I990c1f1dbce95ae4dfc62588c9cc9e1f = (Ibee4f3cd2f516c29ab68e07a640ab65e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8f967710d03870e026564db0df46d146 ;

Ic9c2f173881d25f8976d723957809f51 I273104989bbc820b2b3dcd69886916bd (
.fgallag_sel( Ie495ab560f59ad038992c573de7d2f5b[fgallag_SEL-1:0]),
.fgallag( Ia347d80a70a49605c51d19bc2e696aef ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9d2e71f9a6d7eb4221978fef3c10d678 = (Ie495ab560f59ad038992c573de7d2f5b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia347d80a70a49605c51d19bc2e696aef ;

Ic9c2f173881d25f8976d723957809f51 I32a985892267ffdfd05d1642a543c8bc (
.fgallag_sel( Ibd812def78c3a9c02f9ba45cc0413711[fgallag_SEL-1:0]),
.fgallag( I730db85d3d11d8327c6d48b8b87a00a4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I34754a80000aa92f8a7e4997b91f6d07 = (Ibd812def78c3a9c02f9ba45cc0413711[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I730db85d3d11d8327c6d48b8b87a00a4 ;

Ic9c2f173881d25f8976d723957809f51 If6925d633ff1419f91f29fc5972458ec (
.fgallag_sel( I98166634dc80201b0cefb01d9559c228[fgallag_SEL-1:0]),
.fgallag( I5c6a3ec08cb17d6646bb3e63411a9698 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I055273589d8d967bd5e255808051a101 = (I98166634dc80201b0cefb01d9559c228[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5c6a3ec08cb17d6646bb3e63411a9698 ;

Ic9c2f173881d25f8976d723957809f51 I588cddf91a30b19ecdd088ca9e3f3c96 (
.fgallag_sel( Ic2f03a980b5f0b042853ca746abab22b[fgallag_SEL-1:0]),
.fgallag( I7b5baeec7b11eca457dcd9d2b2b64ac5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5142a2511a55a7ad420618d874b0dddd = (Ic2f03a980b5f0b042853ca746abab22b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7b5baeec7b11eca457dcd9d2b2b64ac5 ;

Ic9c2f173881d25f8976d723957809f51 I9a48d8c36c68b02180ca67a4e5ef01bf (
.fgallag_sel( I2807a88097d2683ebdb9e0e785e3af02[fgallag_SEL-1:0]),
.fgallag( Ic4c7a9d491c560d7b6c410d8216f59bf ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5e008272bf3a470d74ca6b5cf39bf28f = (I2807a88097d2683ebdb9e0e785e3af02[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic4c7a9d491c560d7b6c410d8216f59bf ;

Ic9c2f173881d25f8976d723957809f51 Ie2edd957842af319f726eea427aa8276 (
.fgallag_sel( I8bebbb3a676c8506af0768516abcd740[fgallag_SEL-1:0]),
.fgallag( I2151735079b41a7f8cbfe2b93f1b7470 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5c31bbaf08a6e8971f585cdae36384f5 = (I8bebbb3a676c8506af0768516abcd740[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2151735079b41a7f8cbfe2b93f1b7470 ;

Ic9c2f173881d25f8976d723957809f51 Ic4e86616964de49adb76c9081d3b0c0e (
.fgallag_sel( I31d380f34691c9fe9022035f233b77e2[fgallag_SEL-1:0]),
.fgallag( Ia69e34af60619fa04e8478e2d04768bb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I509af9c5f9d6bf3be233847dbd05e3fa = (I31d380f34691c9fe9022035f233b77e2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia69e34af60619fa04e8478e2d04768bb ;

Ic9c2f173881d25f8976d723957809f51 I4e8ae43a78e1ba9503506aa4f3441f4b (
.fgallag_sel( I1ffb5675c98ab5b3c62b24eb23441473[fgallag_SEL-1:0]),
.fgallag( I7f9984597d0e7bcda92f13fbb8805687 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3182472e08e707cbc36d60ba54613129 = (I1ffb5675c98ab5b3c62b24eb23441473[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7f9984597d0e7bcda92f13fbb8805687 ;

Ic9c2f173881d25f8976d723957809f51 I903eb140aabe11913ecc9463f6183e6d (
.fgallag_sel( If56424546ec4f3445853538207ea864e[fgallag_SEL-1:0]),
.fgallag( I342ef25fefdb6a326dac80d76052bbd9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If2455c2d04521a8d8c59965759eb328b = (If56424546ec4f3445853538207ea864e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I342ef25fefdb6a326dac80d76052bbd9 ;

Ic9c2f173881d25f8976d723957809f51 I4e872c070f9ee144d84a53fcad006e2e (
.fgallag_sel( I31a49be4a34d9bac2e0d815097439772[fgallag_SEL-1:0]),
.fgallag( Id1414254ab35ee805c4010432eb24243 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib759c72355cd6e146edb26ad106a0418 = (I31a49be4a34d9bac2e0d815097439772[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id1414254ab35ee805c4010432eb24243 ;

Ic9c2f173881d25f8976d723957809f51 I2afbd832bb84a19568aa5a3bdaff5cae (
.fgallag_sel( I6b96a2498078953e87de223aa2236d50[fgallag_SEL-1:0]),
.fgallag( I8db7cc6cb4bf55131bee6b00e76baf46 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6826c8a05953c4df79e31a19adfa2693 = (I6b96a2498078953e87de223aa2236d50[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8db7cc6cb4bf55131bee6b00e76baf46 ;

Ic9c2f173881d25f8976d723957809f51 I46c8a60fb5804c089a8a91dbc788f21c (
.fgallag_sel( I79bf36e298a85a42c7432f877055f0b4[fgallag_SEL-1:0]),
.fgallag( I355aec2468fa96e2f32c8c324c48c5f5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I56122ba51d99f9ca67828649860d409e = (I79bf36e298a85a42c7432f877055f0b4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I355aec2468fa96e2f32c8c324c48c5f5 ;

Ic9c2f173881d25f8976d723957809f51 I6ae7f1a86df8dd91a6a06f5173b57d1c (
.fgallag_sel( I90c070b9bde5da05e8a5d25d2de3ba6b[fgallag_SEL-1:0]),
.fgallag( Ic45ea6e09fd20a2285b7e6e2507910f4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1bcda37ae1a26452a3443142fbee54f9 = (I90c070b9bde5da05e8a5d25d2de3ba6b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic45ea6e09fd20a2285b7e6e2507910f4 ;

Ic9c2f173881d25f8976d723957809f51 I6d8a1165a1b88a9a35f625e8e644be1f (
.fgallag_sel( I28d0e4e6d772dd58d845d91952ada300[fgallag_SEL-1:0]),
.fgallag( I288b192ad6d04370df8084511c7f44ce ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3f7dda67dc14fdf45bfb9c4e01dd7f38 = (I28d0e4e6d772dd58d845d91952ada300[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I288b192ad6d04370df8084511c7f44ce ;

Ic9c2f173881d25f8976d723957809f51 I5c611a471a62b31bb9b6ea6c2284d526 (
.fgallag_sel( I7232b4e277acc6f1acefcb606ca24508[fgallag_SEL-1:0]),
.fgallag( I4d589e9479ee494636d90a910e530863 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6fd4da8e1e3cb360964d6e425d174465 = (I7232b4e277acc6f1acefcb606ca24508[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4d589e9479ee494636d90a910e530863 ;

Ic9c2f173881d25f8976d723957809f51 Idcba369fe9af4b0c4331e464da884c6d (
.fgallag_sel( I32da124c433c55f692ffa4734d0dc8fc[fgallag_SEL-1:0]),
.fgallag( Ib8fcb6e6569d34c67145861431ad5334 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5f7baab0fcf12df1e886e17375732c04 = (I32da124c433c55f692ffa4734d0dc8fc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib8fcb6e6569d34c67145861431ad5334 ;

Ic9c2f173881d25f8976d723957809f51 I2699611aa477270ee42894b065336c12 (
.fgallag_sel( I56e487db14eeb8d93f494d2f11b57a49[fgallag_SEL-1:0]),
.fgallag( I5405b3c646988338f12191bb8cb02205 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I87303a5c7e205b0b1b196ae97a0c994f = (I56e487db14eeb8d93f494d2f11b57a49[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5405b3c646988338f12191bb8cb02205 ;

Ic9c2f173881d25f8976d723957809f51 I73b0f431362e5dcf8e2affa740e48b80 (
.fgallag_sel( I94d3c02bd5b8e84926d4b3c2f56efeac[fgallag_SEL-1:0]),
.fgallag( I371946ff4a809b62ceed2334a9656787 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5ebd9eab33e2e8cd6b2f7c1f3bd2e39f = (I94d3c02bd5b8e84926d4b3c2f56efeac[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I371946ff4a809b62ceed2334a9656787 ;

Ic9c2f173881d25f8976d723957809f51 I63e0a4fa13588981cc131d37156dcac3 (
.fgallag_sel( I0c35b2e9176f9a06e26ca67d036411b4[fgallag_SEL-1:0]),
.fgallag( I6d5be8ddd471c1ddf781949169bd9807 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7f4bd63152869ed52c49aa41eea5ea1e = (I0c35b2e9176f9a06e26ca67d036411b4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6d5be8ddd471c1ddf781949169bd9807 ;

Ic9c2f173881d25f8976d723957809f51 I42a5fbf7dbf99f1f636c13cb623e77f5 (
.fgallag_sel( Ia6ee7b70d0b7fe7c346760b1784e50b9[fgallag_SEL-1:0]),
.fgallag( I499f6bbf3456d23378ff02b6f65a5ae4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id243e47daf8a5e75fe52a828af95b5aa = (Ia6ee7b70d0b7fe7c346760b1784e50b9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I499f6bbf3456d23378ff02b6f65a5ae4 ;

Ic9c2f173881d25f8976d723957809f51 I159448573c2ef7f74c065c3594229e62 (
.fgallag_sel( I7ce57c278c683ad045526e49bcc47412[fgallag_SEL-1:0]),
.fgallag( I0c81821914371a777679053e2aa5a55e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I62bd2c30206c591bcb87f31543bda72e = (I7ce57c278c683ad045526e49bcc47412[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0c81821914371a777679053e2aa5a55e ;

Ic9c2f173881d25f8976d723957809f51 I483a97fdbd014be94ce553768bd54ff7 (
.fgallag_sel( Ie3d3e681cac0bb919946ac27057409e2[fgallag_SEL-1:0]),
.fgallag( Ief591e9d4759a4b1059574bb624e4ce6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic1238f5f1f2011fa1869cdb2f50e6a30 = (Ie3d3e681cac0bb919946ac27057409e2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ief591e9d4759a4b1059574bb624e4ce6 ;

Ic9c2f173881d25f8976d723957809f51 I041c8cc1fb58a5a3beec7cb7c67c3deb (
.fgallag_sel( I8ea0a8cdd6506c982ad75f23136bcebe[fgallag_SEL-1:0]),
.fgallag( Ie40648c85ed87c979a54dfc1f85d1cc8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7f2885836616ac775eb9406e8f5d5214 = (I8ea0a8cdd6506c982ad75f23136bcebe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie40648c85ed87c979a54dfc1f85d1cc8 ;

Ic9c2f173881d25f8976d723957809f51 I40e446d0a9e67baf02d83de201d99ab5 (
.fgallag_sel( Ic812f8bc775c5ee6a83e2b9aeb22b2a4[fgallag_SEL-1:0]),
.fgallag( I36956634f94d6053aa455b29bc0b7a0f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If1608747d211db3fdf51ecf7464c494c = (Ic812f8bc775c5ee6a83e2b9aeb22b2a4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I36956634f94d6053aa455b29bc0b7a0f ;

Ic9c2f173881d25f8976d723957809f51 I649f099d2f0d4fef8672ff7f4af29f34 (
.fgallag_sel( I0f0adf7fe957b9a68772bd8a1bc163d4[fgallag_SEL-1:0]),
.fgallag( I05a652e83a9b8c2c38de64de6a70f8bc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iccd84e19d39b19bec98dad532ea5b3ce = (I0f0adf7fe957b9a68772bd8a1bc163d4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I05a652e83a9b8c2c38de64de6a70f8bc ;

Ic9c2f173881d25f8976d723957809f51 Ia29511dffc38f7ccb2c9f2b3f7c4976b (
.fgallag_sel( If09562f8d82bc1dea7c38ed51523a889[fgallag_SEL-1:0]),
.fgallag( Iaefa87388884b85eed690e9917bc9d5b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idf7e508a586310bf4ca23c84f8240691 = (If09562f8d82bc1dea7c38ed51523a889[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaefa87388884b85eed690e9917bc9d5b ;

Ic9c2f173881d25f8976d723957809f51 I9b31fd53fc97ebaa28e18dfbf651d9ff (
.fgallag_sel( Ib0fd21d66cd89c4e5c95fbc9c7680b62[fgallag_SEL-1:0]),
.fgallag( I98836c38732b8da439946aa5fcbbd963 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic8ef3162d3d0c57faf5dd1bddef1622a = (Ib0fd21d66cd89c4e5c95fbc9c7680b62[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I98836c38732b8da439946aa5fcbbd963 ;

Ic9c2f173881d25f8976d723957809f51 I5bd1dce1a542ea17b51cff8432d5eb13 (
.fgallag_sel( I5a2b2bfadc638fe3fdc31136a8f09a8d[fgallag_SEL-1:0]),
.fgallag( I8ff116e234a1007cc47989f3fdcf88d6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I68115420b3b9b8ca8ca584c260e924ec = (I5a2b2bfadc638fe3fdc31136a8f09a8d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8ff116e234a1007cc47989f3fdcf88d6 ;

Ic9c2f173881d25f8976d723957809f51 Ib7d1dc61f7e873beba51137590ea2d6d (
.fgallag_sel( Ica914d8c556285d6b90b35747065a6e5[fgallag_SEL-1:0]),
.fgallag( I53dfee31709f8eca30897d6bf1618418 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5bac906cb51bae905ea33717fe015201 = (Ica914d8c556285d6b90b35747065a6e5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I53dfee31709f8eca30897d6bf1618418 ;

Ic9c2f173881d25f8976d723957809f51 Ib62fdbcf78f57e89352048407087c4d9 (
.fgallag_sel( I00c5d739bccb0ab6d05da70fe51aafea[fgallag_SEL-1:0]),
.fgallag( I3ac389b6b81baf93095cc3e9e9c3d8ef ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9f261cb4883275f5f9187a1a6e8fee08 = (I00c5d739bccb0ab6d05da70fe51aafea[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3ac389b6b81baf93095cc3e9e9c3d8ef ;

Ic9c2f173881d25f8976d723957809f51 I76810b99ccf11161d098661f993816bb (
.fgallag_sel( I18e448761bc014ce490b766183350312[fgallag_SEL-1:0]),
.fgallag( Ief52e91e9170809b980aa881bf76957a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iecfe32305d22e6d91c3f7d4af2ad9d2f = (I18e448761bc014ce490b766183350312[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ief52e91e9170809b980aa881bf76957a ;

Ic9c2f173881d25f8976d723957809f51 If7ef49486039067dc7c000014592376a (
.fgallag_sel( I1b5920f488e9469bd416a6af3072a30b[fgallag_SEL-1:0]),
.fgallag( Iebf813928bcad8ee3b6911057c59752b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib30aa869fd577fb3315608a85947dc7d = (I1b5920f488e9469bd416a6af3072a30b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iebf813928bcad8ee3b6911057c59752b ;

Ic9c2f173881d25f8976d723957809f51 I20936cbcf6ff7fcaebc35bb1bddff027 (
.fgallag_sel( I70b41ffed4b6d88ddff219c567b8e968[fgallag_SEL-1:0]),
.fgallag( I57ae0d331753595cd56d45a28cd5c790 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I82209dd60aeaffa4b05b38230c27147b = (I70b41ffed4b6d88ddff219c567b8e968[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I57ae0d331753595cd56d45a28cd5c790 ;

Ic9c2f173881d25f8976d723957809f51 Id0f11df9edf86d7390939518bf0727e8 (
.fgallag_sel( I935e083b4561da7d015e98ca7f02854e[fgallag_SEL-1:0]),
.fgallag( Ibd173152b9400b4c8011451d68b07e4c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifa110a9cdb359c2b0567d25d4dba725a = (I935e083b4561da7d015e98ca7f02854e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibd173152b9400b4c8011451d68b07e4c ;

Ic9c2f173881d25f8976d723957809f51 I63789eadd367958852651d2257ad9658 (
.fgallag_sel( Iaca9ef263bf220d786242b88c994fd21[fgallag_SEL-1:0]),
.fgallag( Idc21b018b7b6f2e0bc627e8968e06eda ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1451eec261d2367ec6e7b2d50a20679a = (Iaca9ef263bf220d786242b88c994fd21[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idc21b018b7b6f2e0bc627e8968e06eda ;

Ic9c2f173881d25f8976d723957809f51 I8e6886fc4de36e40170208325c87af29 (
.fgallag_sel( I92169291959eb33452b79bfd32618cbc[fgallag_SEL-1:0]),
.fgallag( I783423950d0e0229826b2249f5cfdf5c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id8f178b6565e3a57c5370aaad14f0639 = (I92169291959eb33452b79bfd32618cbc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I783423950d0e0229826b2249f5cfdf5c ;

Ic9c2f173881d25f8976d723957809f51 I6cb0d3275b8f070d5e9f9a6c5efb5949 (
.fgallag_sel( I126dabc3ebb9c4157adf62b57f217bd0[fgallag_SEL-1:0]),
.fgallag( I6b8fc6d29fb4549e3f191f913bccff9e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I67fb672706bbd331c27ab1eb386c24b5 = (I126dabc3ebb9c4157adf62b57f217bd0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6b8fc6d29fb4549e3f191f913bccff9e ;

Ic9c2f173881d25f8976d723957809f51 Ide4d16fa7756e3cd6cc862d5dff2bd1d (
.fgallag_sel( If4433b1ef2eb963cd301946958b69884[fgallag_SEL-1:0]),
.fgallag( Idc98380b110c22495027a7cdb6f2029d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I112661c3273bde5c91b800dd8ddb08a9 = (If4433b1ef2eb963cd301946958b69884[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idc98380b110c22495027a7cdb6f2029d ;

Ic9c2f173881d25f8976d723957809f51 I4fa55c0c4074f9fea3e89a7229a5ddb9 (
.fgallag_sel( I67ac5b9b794787b3c4738c3366689871[fgallag_SEL-1:0]),
.fgallag( Ieb72df81e325eda4d80a237454fa9dbd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia4979ed96ea3e7332635e1f1a14d9ed4 = (I67ac5b9b794787b3c4738c3366689871[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ieb72df81e325eda4d80a237454fa9dbd ;

Ic9c2f173881d25f8976d723957809f51 I7f8b57a08c667de76fa25d130bc033ee (
.fgallag_sel( I4f022d70078c412bdbef158f750d3da3[fgallag_SEL-1:0]),
.fgallag( If70e7ed8d4989cd75d37af1dc5d185ed ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I11a094c5fa993419d19f6361157d6ad0 = (I4f022d70078c412bdbef158f750d3da3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If70e7ed8d4989cd75d37af1dc5d185ed ;

Ic9c2f173881d25f8976d723957809f51 I1ad8c2bf20ecbc22512a759064b9716a (
.fgallag_sel( I6be6165385f6a77aeedb88f2baaa9cab[fgallag_SEL-1:0]),
.fgallag( Ifc99661bc592c2c43bae53db10c8d472 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I38007605c51aa852477e1901bdd292f0 = (I6be6165385f6a77aeedb88f2baaa9cab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifc99661bc592c2c43bae53db10c8d472 ;

Ic9c2f173881d25f8976d723957809f51 I39d05df6a4049f5e323b02a271664101 (
.fgallag_sel( Id1f7fe91547e158e1d39edffb1421ff3[fgallag_SEL-1:0]),
.fgallag( Ic8860cc8d323e5a4c68233109ed70512 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icae30bad38ea69b85fa826ad52e25a51 = (Id1f7fe91547e158e1d39edffb1421ff3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic8860cc8d323e5a4c68233109ed70512 ;

Ic9c2f173881d25f8976d723957809f51 I62efe997ac7a7540c103bb4980497d75 (
.fgallag_sel( I7a51924134902612db53941390891245[fgallag_SEL-1:0]),
.fgallag( I439288f09536ca87fa0feb5f6436716e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1afd8ef52cb1eef06769b7a27c95fa03 = (I7a51924134902612db53941390891245[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I439288f09536ca87fa0feb5f6436716e ;

Ic9c2f173881d25f8976d723957809f51 I72b39192af0e0999a9bb399c090b0fd3 (
.fgallag_sel( I45128b9e29dd2fdd94a78fc5ffdff2b1[fgallag_SEL-1:0]),
.fgallag( I66c4beb8fe2d9f363c8e153a12f216ca ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9c5442889b71c19de290cf33fa393bd9 = (I45128b9e29dd2fdd94a78fc5ffdff2b1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I66c4beb8fe2d9f363c8e153a12f216ca ;

Ic9c2f173881d25f8976d723957809f51 Ic57dfea6981ce6ea93c14ac1b01035e1 (
.fgallag_sel( I7f1082408c8ebb5be18e8f71ff9510e5[fgallag_SEL-1:0]),
.fgallag( Ib2a96d55b1f7bf9b89286de32e59fad3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I772891870fc29b32eeed162f198217e9 = (I7f1082408c8ebb5be18e8f71ff9510e5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib2a96d55b1f7bf9b89286de32e59fad3 ;

Ic9c2f173881d25f8976d723957809f51 I9ed6dc4b8751eec9918743e59e64009d (
.fgallag_sel( I655ebf19c2f4b3dde716668f9ce12e59[fgallag_SEL-1:0]),
.fgallag( I3028dabd706c9e5768eac56c66463955 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If4167812b028552487002b44bdae0caa = (I655ebf19c2f4b3dde716668f9ce12e59[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3028dabd706c9e5768eac56c66463955 ;

Ic9c2f173881d25f8976d723957809f51 I391f2aecfea088a35d1fefd024186f4b (
.fgallag_sel( Ibc9d493a507122d92af42d858cdc4c61[fgallag_SEL-1:0]),
.fgallag( I265f3da3571d2ddb786b98ba3959823b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4d470ec03c4967c49989f59671d735bc = (Ibc9d493a507122d92af42d858cdc4c61[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I265f3da3571d2ddb786b98ba3959823b ;

Ic9c2f173881d25f8976d723957809f51 I2728235aa9921a96c20fd4e2e87f02b6 (
.fgallag_sel( Ib3d3103e5ee4feb160a97c7e26f7102b[fgallag_SEL-1:0]),
.fgallag( If8d81c152d863660081339144b37a052 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia28efddccf0f15c926e3901002bf6c9f = (Ib3d3103e5ee4feb160a97c7e26f7102b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If8d81c152d863660081339144b37a052 ;

Ic9c2f173881d25f8976d723957809f51 Ib919e1934f67b036adc5c17d4648206e (
.fgallag_sel( I6cc56b119e72175df3b7ce64dc3d9305[fgallag_SEL-1:0]),
.fgallag( Ie9cba6422546d378655d0ef98ef974fb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1f3c6900aaf35b7e0cf71c04d917cb71 = (I6cc56b119e72175df3b7ce64dc3d9305[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie9cba6422546d378655d0ef98ef974fb ;

Ic9c2f173881d25f8976d723957809f51 I06dfc780ca37944c5585f705b4e42e60 (
.fgallag_sel( I57cf4a9378f1cdd94a1a5608dc57e05f[fgallag_SEL-1:0]),
.fgallag( Iaddf6de71a6329eb536f54e3d18d43d6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8788a098d0d9b94af7b93f6b5ef0cce2 = (I57cf4a9378f1cdd94a1a5608dc57e05f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaddf6de71a6329eb536f54e3d18d43d6 ;

Ic9c2f173881d25f8976d723957809f51 I333b776f6b7b89789cb90ff23a76dab2 (
.fgallag_sel( I4160ab1aa18e8151c0a5c23b9edeb907[fgallag_SEL-1:0]),
.fgallag( I280ed7bf157554fcad915f0e7fa12653 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I46a61c4cc712f8ffcf45f93d11f0e146 = (I4160ab1aa18e8151c0a5c23b9edeb907[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I280ed7bf157554fcad915f0e7fa12653 ;

Ic9c2f173881d25f8976d723957809f51 Ia26c828a625dd02473c0b5c5b75efe22 (
.fgallag_sel( Ia1f183f2d904d006e46399424e06c614[fgallag_SEL-1:0]),
.fgallag( I0ca797b233dcdac8e390e1e41d99b196 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2a826f08bf1fc30c125cdb9a93bea1b3 = (Ia1f183f2d904d006e46399424e06c614[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0ca797b233dcdac8e390e1e41d99b196 ;

Ic9c2f173881d25f8976d723957809f51 I38b714eacc0ad5b277bbe128c15c305a (
.fgallag_sel( If979702738671323995e56108bc9376c[fgallag_SEL-1:0]),
.fgallag( I150792edd72cc07cf8242d787cb52056 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2614ad9be5eee336ad67441c050bd366 = (If979702738671323995e56108bc9376c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I150792edd72cc07cf8242d787cb52056 ;

Ic9c2f173881d25f8976d723957809f51 Iacf9b429789d62f032ee3824d98b8996 (
.fgallag_sel( Ibc96fe0a6bf1f95036f97c7d44fab575[fgallag_SEL-1:0]),
.fgallag( I186c13747ff5a1ee6e562ad9e5faabd9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iecd35290f27c4375873e964f2db90ba9 = (Ibc96fe0a6bf1f95036f97c7d44fab575[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I186c13747ff5a1ee6e562ad9e5faabd9 ;

Ic9c2f173881d25f8976d723957809f51 I1d28d6c4e0497062cb8b9c192d2e59f0 (
.fgallag_sel( I755a38220a693ba43701d30e7e9508ad[fgallag_SEL-1:0]),
.fgallag( I6fb8240f8c68b71cafe4c2c43ac7db33 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9b90edd08194934b456cf88beedf8785 = (I755a38220a693ba43701d30e7e9508ad[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6fb8240f8c68b71cafe4c2c43ac7db33 ;

Ic9c2f173881d25f8976d723957809f51 I60f47f35433f3a6ffd49f5a5331f2db0 (
.fgallag_sel( I896fb82baa9647a14f4b5b1ecfa70a15[fgallag_SEL-1:0]),
.fgallag( I166f5cab59c2a66117f2287d2b11c096 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7db63c5bb5e53cbc83051b5c80c1a19c = (I896fb82baa9647a14f4b5b1ecfa70a15[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I166f5cab59c2a66117f2287d2b11c096 ;

Ic9c2f173881d25f8976d723957809f51 I94345193b88849094fbe9131a1167b97 (
.fgallag_sel( I23d1c973d7a2048353fbb68e4a294c08[fgallag_SEL-1:0]),
.fgallag( Ie896986a747c1cd8ccad7117125c6e0d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iaec5353d68ad9092c0fb74683f876213 = (I23d1c973d7a2048353fbb68e4a294c08[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie896986a747c1cd8ccad7117125c6e0d ;

Ic9c2f173881d25f8976d723957809f51 I3192037148141092fc87106df110e609 (
.fgallag_sel( If9fd1e08af14f2fd4ca363383f48580a[fgallag_SEL-1:0]),
.fgallag( I0c829f14ef188ff7ae1417e28903f2b3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iec7f88e1ed763c1f55c90b39870875c2 = (If9fd1e08af14f2fd4ca363383f48580a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0c829f14ef188ff7ae1417e28903f2b3 ;

Ic9c2f173881d25f8976d723957809f51 Idf341b16ab8af615889226e66bd461a2 (
.fgallag_sel( I8f3782f78d88a5c3bc93709564999b30[fgallag_SEL-1:0]),
.fgallag( I3591d4f320f8401ef8ad8f92d2d89bf6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I32f96b4803590ac0f86d2178cac9e4a8 = (I8f3782f78d88a5c3bc93709564999b30[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3591d4f320f8401ef8ad8f92d2d89bf6 ;

Ic9c2f173881d25f8976d723957809f51 Ic734a34cce503a71197ab291a31584c5 (
.fgallag_sel( I986d61d79ce31f4677f3293339db6ad2[fgallag_SEL-1:0]),
.fgallag( I3816895f23a1381e42aaeb64dd158fda ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idc0fc3de3b05c5beebbf24649662f02e = (I986d61d79ce31f4677f3293339db6ad2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3816895f23a1381e42aaeb64dd158fda ;

Ic9c2f173881d25f8976d723957809f51 I27b47ef81e78b671d50489ee2e212fef (
.fgallag_sel( Ica4d93d9fad21316002008ade5106a9d[fgallag_SEL-1:0]),
.fgallag( Ic9c34a36b2fde9649064680904ec9150 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9d54e626fd0b2e435b117ae6b5d5e194 = (Ica4d93d9fad21316002008ade5106a9d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic9c34a36b2fde9649064680904ec9150 ;

Ic9c2f173881d25f8976d723957809f51 Ide7cb1f73ed9279ba76e40e20d02bf22 (
.fgallag_sel( If77592d5d8bed32477fd690341e543d0[fgallag_SEL-1:0]),
.fgallag( If7eb75eccc5a6384c80d99b64d534fca ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id5cff86905cde551a008a19305e87f94 = (If77592d5d8bed32477fd690341e543d0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If7eb75eccc5a6384c80d99b64d534fca ;

Ic9c2f173881d25f8976d723957809f51 I235283180965f1578ee34e7b470c9119 (
.fgallag_sel( I25b70c6b830cbfe1b41d8f289c751924[fgallag_SEL-1:0]),
.fgallag( Ib788a897a1d1b86b2c16caade11846ee ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3837a2e882da18f37f074b51cf5cbf85 = (I25b70c6b830cbfe1b41d8f289c751924[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib788a897a1d1b86b2c16caade11846ee ;

Ic9c2f173881d25f8976d723957809f51 I5b8c6c6889332682e4d0f848557437d2 (
.fgallag_sel( I2a5d65eeffa18dd9af9fe36463dafd7c[fgallag_SEL-1:0]),
.fgallag( I6a5fec9dad124f6d8c5574bcc2643ede ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib584dc3e5dd346562062794c0f1c5f9e = (I2a5d65eeffa18dd9af9fe36463dafd7c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6a5fec9dad124f6d8c5574bcc2643ede ;

Ic9c2f173881d25f8976d723957809f51 I0f2f2f2cbbb641fd8e40e0ccf385240b (
.fgallag_sel( Ibafa6e10bd4edf5d224fdeb2f9adbf98[fgallag_SEL-1:0]),
.fgallag( I3936f324b08bea1bc5f8bcd12437b161 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I20ac1027f7da12ad62120cd3b0603c7e = (Ibafa6e10bd4edf5d224fdeb2f9adbf98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3936f324b08bea1bc5f8bcd12437b161 ;

Ic9c2f173881d25f8976d723957809f51 I73f2afb2fa48cc332d4085e951661bb7 (
.fgallag_sel( Ifc25402bd879bc5c43b4945b60cd4540[fgallag_SEL-1:0]),
.fgallag( I1a59337d4da3e3ad1a738a9c3b56ef8c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8adacef11a4f33ff1ccea285fd1a8b74 = (Ifc25402bd879bc5c43b4945b60cd4540[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1a59337d4da3e3ad1a738a9c3b56ef8c ;

Ic9c2f173881d25f8976d723957809f51 Ida379f416970ea6b6c2f09c345080aa9 (
.fgallag_sel( Iec48da6882325d8a33e0e0e845eb18a0[fgallag_SEL-1:0]),
.fgallag( Ic3e3b4cba05d80c0ceaa6e25a906a602 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie2ad82bbff584541911e13b90a5d15a0 = (Iec48da6882325d8a33e0e0e845eb18a0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic3e3b4cba05d80c0ceaa6e25a906a602 ;

Ic9c2f173881d25f8976d723957809f51 Ifada4981b64ccb6947d4de0cc39acf3e (
.fgallag_sel( I0fd05e46862fdf8e614afaa3fd478602[fgallag_SEL-1:0]),
.fgallag( Ife0830e12b8bbb5aa0b8c2c0e4191e59 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If6243c5fc2ec9a15eecf227b234434d1 = (I0fd05e46862fdf8e614afaa3fd478602[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ife0830e12b8bbb5aa0b8c2c0e4191e59 ;

Ic9c2f173881d25f8976d723957809f51 I692e1ad2d52079514c739f09a57f82a9 (
.fgallag_sel( I6253a59dca81842d9ab6e58cf204abbf[fgallag_SEL-1:0]),
.fgallag( I95eaa4ac5199ebbb06f780d1376062ec ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I41f34c28805f2653586d89312f73237f = (I6253a59dca81842d9ab6e58cf204abbf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I95eaa4ac5199ebbb06f780d1376062ec ;

Ic9c2f173881d25f8976d723957809f51 I8d6dd6556c44a63b919a1072d2b83a95 (
.fgallag_sel( Ib18d64bc58b354358ee6ac16785880e2[fgallag_SEL-1:0]),
.fgallag( Ib40ccfdb9ea28f333a7cc67f2446c923 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie2031e8a9632f0b98f617232f7c462e6 = (Ib18d64bc58b354358ee6ac16785880e2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib40ccfdb9ea28f333a7cc67f2446c923 ;

Ic9c2f173881d25f8976d723957809f51 If2fb76b7d99f8cc9d42604f0e0f0e7e9 (
.fgallag_sel( I28689b693a7a5f761a1f252aa3ef3b67[fgallag_SEL-1:0]),
.fgallag( I507515355429e697cd5496809aa03cfb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9d706a29e764935ac3cabdac4e95af1d = (I28689b693a7a5f761a1f252aa3ef3b67[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I507515355429e697cd5496809aa03cfb ;

Ic9c2f173881d25f8976d723957809f51 I66b621ae2fcc3dec67c83912b1a671e7 (
.fgallag_sel( I1a4e6d12f9776d5e61094e0b5edf71d9[fgallag_SEL-1:0]),
.fgallag( I6bcc3a323e67f95eb4bf28a0704d3c50 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7a2e1620640d2060cbb0a1bef5eb79c0 = (I1a4e6d12f9776d5e61094e0b5edf71d9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6bcc3a323e67f95eb4bf28a0704d3c50 ;

Ic9c2f173881d25f8976d723957809f51 I23482376cfd437061474738d2688c9e2 (
.fgallag_sel( I8e1ad23b7ac662bb827a83d3709f0adb[fgallag_SEL-1:0]),
.fgallag( I55e3a2566ef3ac257021a294376be634 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2795513c5d99dc8e09be4bebb4d12944 = (I8e1ad23b7ac662bb827a83d3709f0adb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I55e3a2566ef3ac257021a294376be634 ;

Ic9c2f173881d25f8976d723957809f51 Ie58023cf606921b44793ee9cb50f9d23 (
.fgallag_sel( I000ad2287813072cc18dad933758f2ab[fgallag_SEL-1:0]),
.fgallag( I40f10dc3289ea8a59f593f62066aaff8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I03cb6aeff54e7e9e2ee809f8bea621bc = (I000ad2287813072cc18dad933758f2ab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I40f10dc3289ea8a59f593f62066aaff8 ;

Ic9c2f173881d25f8976d723957809f51 Ic3aad8eda928211e1e38deea87cbaa64 (
.fgallag_sel( I7bc3698b51b89ac38ba5f4b5428a0c96[fgallag_SEL-1:0]),
.fgallag( Ieeabde5600d81208346ebd50d4a95d83 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I78c43fed329002e5ab9a0e429fb3b769 = (I7bc3698b51b89ac38ba5f4b5428a0c96[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ieeabde5600d81208346ebd50d4a95d83 ;

Ic9c2f173881d25f8976d723957809f51 Ie733758b1a0e59c1760f4f9a10d7f0f7 (
.fgallag_sel( I78aea1705621e2845a331c3e61a8055b[fgallag_SEL-1:0]),
.fgallag( Ibb9220dcdd6d7fc2b6d6ca5f4cc93a8b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I639755c3c20317c18359e96fce8e2f2e = (I78aea1705621e2845a331c3e61a8055b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibb9220dcdd6d7fc2b6d6ca5f4cc93a8b ;

Ic9c2f173881d25f8976d723957809f51 I1084c1dc44a714a40184f88a216249a4 (
.fgallag_sel( I0a31314c3580f5f9e61e79c133e5d794[fgallag_SEL-1:0]),
.fgallag( I05a3aebc90966144a6809e460d6ceda1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I68c7cb0d5275b576e4021c8aedda4646 = (I0a31314c3580f5f9e61e79c133e5d794[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I05a3aebc90966144a6809e460d6ceda1 ;

Ic9c2f173881d25f8976d723957809f51 Ib3284ee9b23df00773c8538306bae7a4 (
.fgallag_sel( I0e274fd7bfc0388fef95a8ceb939ee91[fgallag_SEL-1:0]),
.fgallag( I7e3150622eb318e94f99b36016ac7d2f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2bd974f363231ecfaa9ef8d018a02936 = (I0e274fd7bfc0388fef95a8ceb939ee91[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7e3150622eb318e94f99b36016ac7d2f ;

Ic9c2f173881d25f8976d723957809f51 I778ca73573d9ad6578f4c6c7248aa2f0 (
.fgallag_sel( Id6f39ddcb73d3f4ec081a365d11d1ef4[fgallag_SEL-1:0]),
.fgallag( Ifb146b2073d447377a1b21fe21baa4da ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I675d5b900c6a4bbdb8f14db50b873893 = (Id6f39ddcb73d3f4ec081a365d11d1ef4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifb146b2073d447377a1b21fe21baa4da ;

Ic9c2f173881d25f8976d723957809f51 I0069104a64f16be3605fef279b326deb (
.fgallag_sel( I807770bfa86d160459d6ec3c0f4d6a0b[fgallag_SEL-1:0]),
.fgallag( Ifa5048ac43025e9cdf3f3436c37bb835 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I36b68c4fcf7a2adafce004ec0e231209 = (I807770bfa86d160459d6ec3c0f4d6a0b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifa5048ac43025e9cdf3f3436c37bb835 ;

Ic9c2f173881d25f8976d723957809f51 Ie01f7781ca23c7222a89c17e4bda03f4 (
.fgallag_sel( I31c89b8a11a3090bfd74b112cbc474bb[fgallag_SEL-1:0]),
.fgallag( I837ba4049e4973924e51d642f7f481ad ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iea5c378e0635e3bb31343988c4dc6259 = (I31c89b8a11a3090bfd74b112cbc474bb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I837ba4049e4973924e51d642f7f481ad ;

Ic9c2f173881d25f8976d723957809f51 I896baab163d64cb884f8f8262ae4453a (
.fgallag_sel( I79b82cb1bfc72bd5a9d313b9e9c9203c[fgallag_SEL-1:0]),
.fgallag( I2910e5e74ca008b7e5502d787cb88a6d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2edf197a22f055871ed9b54f9e1a874a = (I79b82cb1bfc72bd5a9d313b9e9c9203c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2910e5e74ca008b7e5502d787cb88a6d ;

Ic9c2f173881d25f8976d723957809f51 I905e845141c115272695782bf0e65841 (
.fgallag_sel( Ib1046ae03c9a77fd2c0b3e9838e9af87[fgallag_SEL-1:0]),
.fgallag( Ia24816d601e29172628cad0c364b47e9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie80e559352812ffe4d9cf6006af19e85 = (Ib1046ae03c9a77fd2c0b3e9838e9af87[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia24816d601e29172628cad0c364b47e9 ;

Ic9c2f173881d25f8976d723957809f51 I6c39d48f442e45b3ae700e791dc9b71b (
.fgallag_sel( Ic63723fd43cbbbde51c233a3cca15d3f[fgallag_SEL-1:0]),
.fgallag( I8f99af880f329241cfc9616ff9859091 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id2f23da93344ae523d495478dd559ded = (Ic63723fd43cbbbde51c233a3cca15d3f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8f99af880f329241cfc9616ff9859091 ;

Ic9c2f173881d25f8976d723957809f51 I5a99ffd937a6e270674894d1a8d703da (
.fgallag_sel( I3abbb59abada1aec6941185f95f738bd[fgallag_SEL-1:0]),
.fgallag( Iea7c2970a7d80c55c1a6d6933c6c81c9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If18e431ab87f137467f6f87e40b9c27e = (I3abbb59abada1aec6941185f95f738bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iea7c2970a7d80c55c1a6d6933c6c81c9 ;

Ic9c2f173881d25f8976d723957809f51 I2b77d60a0bb9aa7d5697610dbc78d45d (
.fgallag_sel( I8d5bd7039a77ce82ce0f6cbba9c2a076[fgallag_SEL-1:0]),
.fgallag( I75a12697a4ee6de46fc098b0f02b8349 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3f5b5d6b646070d84f2fb963f3824ce1 = (I8d5bd7039a77ce82ce0f6cbba9c2a076[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I75a12697a4ee6de46fc098b0f02b8349 ;

Ic9c2f173881d25f8976d723957809f51 I82faa1701b787abfe4b0973d9beb735c (
.fgallag_sel( I527ad0b9382dd7b6e657dc1a32d8e472[fgallag_SEL-1:0]),
.fgallag( I623d1f0b6829caf5dc0f0eab0ca47f74 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie964e5a463904ac52c4529ffb3ebaf65 = (I527ad0b9382dd7b6e657dc1a32d8e472[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I623d1f0b6829caf5dc0f0eab0ca47f74 ;

Ic9c2f173881d25f8976d723957809f51 I99d16c18fd1091e4e3edbb5297cf5ad2 (
.fgallag_sel( I8de02f32e14e719f4930d99743c04a20[fgallag_SEL-1:0]),
.fgallag( Ieabf207f10f7df1e9059f1e953d7b399 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia74858d5df6a76635e6ba60d0b1a63ea = (I8de02f32e14e719f4930d99743c04a20[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ieabf207f10f7df1e9059f1e953d7b399 ;

Ic9c2f173881d25f8976d723957809f51 I5aae665de42b0494945968f54222a007 (
.fgallag_sel( I7614dd5e9628c761dd9b2a512cb1da98[fgallag_SEL-1:0]),
.fgallag( I1399b55530e343bd85606e7c7529d453 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id9c69999bee621002fa9b387aa809dc5 = (I7614dd5e9628c761dd9b2a512cb1da98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1399b55530e343bd85606e7c7529d453 ;

Ic9c2f173881d25f8976d723957809f51 I2812bd03880296afeb09a82345224d8b (
.fgallag_sel( Icae7efa4742dd0ad943ee1f67b0c9b14[fgallag_SEL-1:0]),
.fgallag( I39ee898ed8a8af64552e1aa145437310 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie9e8ae352a1699484f85ae1e7b7f9246 = (Icae7efa4742dd0ad943ee1f67b0c9b14[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I39ee898ed8a8af64552e1aa145437310 ;

Ic9c2f173881d25f8976d723957809f51 I788db48a598355f85e9bd0ca823aefaf (
.fgallag_sel( Ieb1854b79e9a2bc6cf5aa1c319e8e753[fgallag_SEL-1:0]),
.fgallag( I0af241f9f65af3bff2bb0d69977bb0c6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5a006c73dcb7807d5943857199cc3535 = (Ieb1854b79e9a2bc6cf5aa1c319e8e753[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0af241f9f65af3bff2bb0d69977bb0c6 ;

Ic9c2f173881d25f8976d723957809f51 I6cb9bf0d87818528e564076d819cc8f1 (
.fgallag_sel( Iff50b77f300183ca59a67ccbcc9573c4[fgallag_SEL-1:0]),
.fgallag( I9de68705b5430023d2eb5554370bb188 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idfb53869ea5692adddb6f7452d44effa = (Iff50b77f300183ca59a67ccbcc9573c4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9de68705b5430023d2eb5554370bb188 ;

Ic9c2f173881d25f8976d723957809f51 I7b99a256c8598b0060a3f37b69ed6912 (
.fgallag_sel( I4868604f8178663de759d4c63dc6c4bd[fgallag_SEL-1:0]),
.fgallag( Icdf7ba01c4813abe3cfa760f2d8d5c84 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0d11a8980f8fd7aadc8e48e62a653aa6 = (I4868604f8178663de759d4c63dc6c4bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Icdf7ba01c4813abe3cfa760f2d8d5c84 ;

Ic9c2f173881d25f8976d723957809f51 I8705924ee7188be5c5de6b55b966dcfd (
.fgallag_sel( Ife992a151986c58df4cba79b6bc4ac0a[fgallag_SEL-1:0]),
.fgallag( Ia6b995eb6bbaad8a638c80d587d45ab9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib843721cd2106b7e5cc21812aeb374eb = (Ife992a151986c58df4cba79b6bc4ac0a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia6b995eb6bbaad8a638c80d587d45ab9 ;

Ic9c2f173881d25f8976d723957809f51 Ifc82648fa5aa0d28da501a0927ac34a1 (
.fgallag_sel( I9ab973fb74d9fac5d78eb8fc2c7ecf36[fgallag_SEL-1:0]),
.fgallag( I75c2987dcebc9cdca578aeebec96fccc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I400d30374ae90fa066db0f5a29195e4e = (I9ab973fb74d9fac5d78eb8fc2c7ecf36[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I75c2987dcebc9cdca578aeebec96fccc ;

Ic9c2f173881d25f8976d723957809f51 I9fefbe9fc9b7c7fe92a4e955137b5db9 (
.fgallag_sel( I5ee7916e859b86a98538659401685016[fgallag_SEL-1:0]),
.fgallag( I6fab90e9a0f606d7c26346c89c6f1d47 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I49316949f603c233556dfe520b9e1a61 = (I5ee7916e859b86a98538659401685016[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6fab90e9a0f606d7c26346c89c6f1d47 ;

Ic9c2f173881d25f8976d723957809f51 Ie8e321169776dd0533e472dc4263470d (
.fgallag_sel( I48c284cefb8cfb5a938a8f23ce4d7f03[fgallag_SEL-1:0]),
.fgallag( Iab2f70a1d3093b3194e9047a8fe8e487 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I57c335ac00303b6df3bb5bc5a1b1bcb6 = (I48c284cefb8cfb5a938a8f23ce4d7f03[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iab2f70a1d3093b3194e9047a8fe8e487 ;

Ic9c2f173881d25f8976d723957809f51 I3fcf37dcb28dce06e13be02b3d198ff2 (
.fgallag_sel( I5c1fc666b77a689478654dd29519f458[fgallag_SEL-1:0]),
.fgallag( Ic84b6224be8eb8eefc9ad9bcc2280291 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I177fce9af9d7a8e9e9dfe423c8abe225 = (I5c1fc666b77a689478654dd29519f458[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic84b6224be8eb8eefc9ad9bcc2280291 ;

Ic9c2f173881d25f8976d723957809f51 I34856b40f036cbd78477d71779e982ed (
.fgallag_sel( I38bba98b59184c75ba3b27e1dcf52182[fgallag_SEL-1:0]),
.fgallag( I64a0e60fdcc93d84606774196b2b7598 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I335535f77c13df799b6e5f9613607a9b = (I38bba98b59184c75ba3b27e1dcf52182[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I64a0e60fdcc93d84606774196b2b7598 ;

Ic9c2f173881d25f8976d723957809f51 I28247ab7b49bb8bcc9b5c63f2491c80a (
.fgallag_sel( I6905b65403c16b0211643227ece536f6[fgallag_SEL-1:0]),
.fgallag( Iaa6a4f3826d87e43dd3213dc5083184b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icbe54351ad1360193ea28dc76e073f23 = (I6905b65403c16b0211643227ece536f6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaa6a4f3826d87e43dd3213dc5083184b ;

Ic9c2f173881d25f8976d723957809f51 Ib824a6c02cc6ad60af6b950a37a0ffc0 (
.fgallag_sel( I3ed34401bba9d5f229bc98480aedd9a5[fgallag_SEL-1:0]),
.fgallag( I94fd5b790a9dceab1b4b3f1b5e30a0d9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I812a6ce8adb2ef9a2a9eb7e7e8cc96f1 = (I3ed34401bba9d5f229bc98480aedd9a5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I94fd5b790a9dceab1b4b3f1b5e30a0d9 ;

Ic9c2f173881d25f8976d723957809f51 I5f3d33b3a52acc415c733101b700a1e5 (
.fgallag_sel( Ib4d05804277cddc7f00ac17ac14f5325[fgallag_SEL-1:0]),
.fgallag( I9c8c1d22021bbe798b1863ae1dfc3965 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I87a99623e8305e331ca590dc62df5252 = (Ib4d05804277cddc7f00ac17ac14f5325[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9c8c1d22021bbe798b1863ae1dfc3965 ;

Ic9c2f173881d25f8976d723957809f51 Id1f60f2bf97e2b1c41124c22e6f010fe (
.fgallag_sel( I41babdca6d3fa462849592d37b0a7998[fgallag_SEL-1:0]),
.fgallag( I870366e9c3b29c1683a7528f4b5d5329 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I130df8a2e7e3e33055f2f2997e6d5716 = (I41babdca6d3fa462849592d37b0a7998[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I870366e9c3b29c1683a7528f4b5d5329 ;

Ic9c2f173881d25f8976d723957809f51 Idbf4e860c56db5381781e8d467721aea (
.fgallag_sel( I58cfec706dc929ebfdeaca6e01b00c0a[fgallag_SEL-1:0]),
.fgallag( I066db3b79f8b4581f96567d943a7e7db ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I07ee1ac328d24e8fa9862659903fd379 = (I58cfec706dc929ebfdeaca6e01b00c0a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I066db3b79f8b4581f96567d943a7e7db ;

Ic9c2f173881d25f8976d723957809f51 I3a98a5a8a463b424f00cd3239f8147d0 (
.fgallag_sel( I7efe3c5b2fc69840a79545e0399ce749[fgallag_SEL-1:0]),
.fgallag( Iabd6f58c4760c939dfd58e4f426bcab9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idd74d5e61d5397193aaf3cdb96dbc84b = (I7efe3c5b2fc69840a79545e0399ce749[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iabd6f58c4760c939dfd58e4f426bcab9 ;

Ic9c2f173881d25f8976d723957809f51 I67c0b8b12739e8c4b382ce6fb961eb92 (
.fgallag_sel( I70e3eeb2b3966676d16a6aa4c85753ab[fgallag_SEL-1:0]),
.fgallag( Ia3505661cb9b7eacbd47774346d12f5b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id74f690142fb1e4a04fa3dca841979a6 = (I70e3eeb2b3966676d16a6aa4c85753ab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia3505661cb9b7eacbd47774346d12f5b ;

Ic9c2f173881d25f8976d723957809f51 I802e13c43ce86fbbe9b0a016f60f6356 (
.fgallag_sel( I2a32d545d1e7beecc7531174c7e8dfbc[fgallag_SEL-1:0]),
.fgallag( I4e7245fc882e3e284d8c152c8998b028 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8327851510864c943e64c3d22b456152 = (I2a32d545d1e7beecc7531174c7e8dfbc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4e7245fc882e3e284d8c152c8998b028 ;

Ic9c2f173881d25f8976d723957809f51 I2928494ba451ec10d9c5cc52bef878fd (
.fgallag_sel( Ib8fb40e4ba0ba1f5e9f5a99d1271ed06[fgallag_SEL-1:0]),
.fgallag( Ibe962754759204890883a6de0993a64b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4f37cf4b922e288365376a45753c4a38 = (Ib8fb40e4ba0ba1f5e9f5a99d1271ed06[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibe962754759204890883a6de0993a64b ;

Ic9c2f173881d25f8976d723957809f51 I1185cfafc4a35cab3313c02b12aabed0 (
.fgallag_sel( Ica792cb9850a61fa4a8bd8a4b6c6ca05[fgallag_SEL-1:0]),
.fgallag( Id2ef1e193163adc702763541f37fec4d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If50168d2535d752dd95301bfe723db9a = (Ica792cb9850a61fa4a8bd8a4b6c6ca05[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id2ef1e193163adc702763541f37fec4d ;

Ic9c2f173881d25f8976d723957809f51 I69677fd02e4058e63683fb89e8bcaed0 (
.fgallag_sel( I779e5997c66649d6d54fd7f0514c47bd[fgallag_SEL-1:0]),
.fgallag( I8a925721cf106d4e6ca1f69bbc2f53d4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6eb5641a21e34b4ced1cf124c3f23646 = (I779e5997c66649d6d54fd7f0514c47bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8a925721cf106d4e6ca1f69bbc2f53d4 ;

Ic9c2f173881d25f8976d723957809f51 I7419d5fb278a3481e7770e72c6e6a823 (
.fgallag_sel( I5aa578b0c2831453683fa44af1878cb8[fgallag_SEL-1:0]),
.fgallag( Ib97671e4daa1b606aa01c5e8f753a9e8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I94da98c2f9e0c8be8ab8f23a2a10095b = (I5aa578b0c2831453683fa44af1878cb8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib97671e4daa1b606aa01c5e8f753a9e8 ;

Ic9c2f173881d25f8976d723957809f51 I685b7482e4fc2b9aaa713b611788a7af (
.fgallag_sel( I735d6229ef1a4ecda0a1f1dbdfb53fc1[fgallag_SEL-1:0]),
.fgallag( Icdd0962fd06355a7dcbb491543eb9cb6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I339ec0bef37cb2e72e8e8795686da0c4 = (I735d6229ef1a4ecda0a1f1dbdfb53fc1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Icdd0962fd06355a7dcbb491543eb9cb6 ;

Ic9c2f173881d25f8976d723957809f51 I9522583999e15d4303351ee93d9a7eb8 (
.fgallag_sel( I62affd47512c5e8f0979244115624d97[fgallag_SEL-1:0]),
.fgallag( I003f9dc1b83f386f070b0a2e8c7ce4f4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If7c621d8183ce83092644a1d80d6c77b = (I62affd47512c5e8f0979244115624d97[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I003f9dc1b83f386f070b0a2e8c7ce4f4 ;

Ic9c2f173881d25f8976d723957809f51 I1a7205d4e2d08226dd95883a761e9345 (
.fgallag_sel( I14fe27afb3df5531b18dc9604e8dbe65[fgallag_SEL-1:0]),
.fgallag( I66e8ad34c764833f038cff700a237fcb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icb4d6012447eb0d6bfa8e8b3f88f0ff9 = (I14fe27afb3df5531b18dc9604e8dbe65[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I66e8ad34c764833f038cff700a237fcb ;

Ic9c2f173881d25f8976d723957809f51 I0ee8b1e1f6eedd5ddc1aa524695c8aa9 (
.fgallag_sel( Ib1b1626c84dad8ad13c058f921ffd57d[fgallag_SEL-1:0]),
.fgallag( I614bddda696787a552e28cfaa81a3aa3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If7c3b54bc0cce4eecf8f55fcf4a5a588 = (Ib1b1626c84dad8ad13c058f921ffd57d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I614bddda696787a552e28cfaa81a3aa3 ;

Ic9c2f173881d25f8976d723957809f51 Ib617d09840f4c0e115a4e7444158ee00 (
.fgallag_sel( Idf4a4bdddb88c21c5afe10a02373a6eb[fgallag_SEL-1:0]),
.fgallag( I38c22e6b7c066be10ec1f8929dbf88f9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1ffe02eedf41df8b947a285adc220fea = (Idf4a4bdddb88c21c5afe10a02373a6eb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I38c22e6b7c066be10ec1f8929dbf88f9 ;

Ic9c2f173881d25f8976d723957809f51 Ife5ac9ba42c4ed053033434b51475069 (
.fgallag_sel( Iadefc2a3d07ed4b2c3c46b2ab5dec252[fgallag_SEL-1:0]),
.fgallag( I245816ec4a0392af2cfa4b44a4e93610 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icd8c721f78cfbefbf25c2e094927401a = (Iadefc2a3d07ed4b2c3c46b2ab5dec252[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I245816ec4a0392af2cfa4b44a4e93610 ;

Ic9c2f173881d25f8976d723957809f51 I5df1cbdbc3e1f426b7330bb21dc4da7a (
.fgallag_sel( I19315957077b037ffc6415dbb06ef789[fgallag_SEL-1:0]),
.fgallag( I83253182662d56779685c9742f55789f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie139a6a80ab0051c5d951103b1554338 = (I19315957077b037ffc6415dbb06ef789[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I83253182662d56779685c9742f55789f ;

Ic9c2f173881d25f8976d723957809f51 I3912fb7493a803bd1dcf13d453763182 (
.fgallag_sel( I1f9be09334407fc86c83a7c127e17bbe[fgallag_SEL-1:0]),
.fgallag( I963a4391dba3d12756b89dda1e962c3f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I993fd34b89fe9b0af3348cdd91ecf025 = (I1f9be09334407fc86c83a7c127e17bbe[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I963a4391dba3d12756b89dda1e962c3f ;

Ic9c2f173881d25f8976d723957809f51 Ia1fafa5d6d7bde1e7bf227b0687ebeed (
.fgallag_sel( I28e17a5af7a7286a2643100d6d058dc0[fgallag_SEL-1:0]),
.fgallag( Ie959690f46f82cbb15ae0cee69f3135f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib5d321981c2997b3635fd0b342993d38 = (I28e17a5af7a7286a2643100d6d058dc0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie959690f46f82cbb15ae0cee69f3135f ;

Ic9c2f173881d25f8976d723957809f51 I46672afa95bec8767585f4d0bedeef80 (
.fgallag_sel( Icb2297c397bfe56be251ffb6b249a020[fgallag_SEL-1:0]),
.fgallag( Ic475c578935fa69db2b1c834539750af ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If1660e858bdb3b0c8a4c1f93f4fe037a = (Icb2297c397bfe56be251ffb6b249a020[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic475c578935fa69db2b1c834539750af ;

Ic9c2f173881d25f8976d723957809f51 Ic75469b06325133a70e411106676b96c (
.fgallag_sel( I64a48984527d660002f1f82c376c7a84[fgallag_SEL-1:0]),
.fgallag( I4f9bc0f2aeafb89fbaa0d0af7dbda06a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7d9ab0daacce00542083a30a35297207 = (I64a48984527d660002f1f82c376c7a84[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4f9bc0f2aeafb89fbaa0d0af7dbda06a ;

Ic9c2f173881d25f8976d723957809f51 Iee4ea7243a35c90a4d8997fa5f1db552 (
.fgallag_sel( I238b5fc70ce9f05b6322a2691b3a0207[fgallag_SEL-1:0]),
.fgallag( I393fa73117dcbf1fb1b74ea1fc7e6c99 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9761f2282bcb9637892cf898b928126c = (I238b5fc70ce9f05b6322a2691b3a0207[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I393fa73117dcbf1fb1b74ea1fc7e6c99 ;

Ic9c2f173881d25f8976d723957809f51 I8dd142af5e4e73055bfe517ce5df7d29 (
.fgallag_sel( I00c16e7ad3821981032a42d5baa767b3[fgallag_SEL-1:0]),
.fgallag( I95836c571386b3b6de07c9195932fe22 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I25de2ab105b6cdb0e30ca97822109fbd = (I00c16e7ad3821981032a42d5baa767b3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I95836c571386b3b6de07c9195932fe22 ;

Ic9c2f173881d25f8976d723957809f51 I261eadaec5d888737a083566e0357d40 (
.fgallag_sel( I42fd5b094da200b33036e6cb8c7d0286[fgallag_SEL-1:0]),
.fgallag( I6dd6f9abc962974c292d22f17a21a936 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I23c14408deedeecba4753f182549adf7 = (I42fd5b094da200b33036e6cb8c7d0286[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6dd6f9abc962974c292d22f17a21a936 ;

Ic9c2f173881d25f8976d723957809f51 I9b821574f18208fdbac6287e4803d1a4 (
.fgallag_sel( I98b7e26a0e9ec9ad750ff87cc0641a73[fgallag_SEL-1:0]),
.fgallag( I9f9e6bc8d2cc6e41813d42ffcd5cff01 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id208387ab734f8ccfaf1567e6b00a4a6 = (I98b7e26a0e9ec9ad750ff87cc0641a73[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9f9e6bc8d2cc6e41813d42ffcd5cff01 ;

Ic9c2f173881d25f8976d723957809f51 I25eb8ba807b33f50d0c5128d114bd2d3 (
.fgallag_sel( I3ec904916870171bf837e162d1030052[fgallag_SEL-1:0]),
.fgallag( I2ba75ccf97b5caf5aa676a9e3c42a366 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I54e43b8da49648867403cf839e87a9ec = (I3ec904916870171bf837e162d1030052[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2ba75ccf97b5caf5aa676a9e3c42a366 ;

Ic9c2f173881d25f8976d723957809f51 I46661d94a102017ccb9c2d06b884a1d1 (
.fgallag_sel( Iedb11b97900b7dd769d31f8a89521975[fgallag_SEL-1:0]),
.fgallag( I006699f0e016e7022b2706751965c42c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I66c8b8649e7997b7e4c9c17f7c0b17b7 = (Iedb11b97900b7dd769d31f8a89521975[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I006699f0e016e7022b2706751965c42c ;

Ic9c2f173881d25f8976d723957809f51 Ia66fa1ec5a72391302d5c5ddcfbdeb60 (
.fgallag_sel( Id0dceec6497c9f13ada07138986d4145[fgallag_SEL-1:0]),
.fgallag( I66d5992f4f39337782cfbbb9fec3b2c8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9a0093065fb4cf517f1e7b75b3080b1c = (Id0dceec6497c9f13ada07138986d4145[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I66d5992f4f39337782cfbbb9fec3b2c8 ;

Ic9c2f173881d25f8976d723957809f51 I7db4d75fc23b77d4b5013c95e9469f8a (
.fgallag_sel( Ibfe7d9bac29b8838f20cdcfe8ef7da0c[fgallag_SEL-1:0]),
.fgallag( Ie5f503c91ddf6eff2b9645e6e3c22b2e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I72d18b26784448b5514e66251bb19ebd = (Ibfe7d9bac29b8838f20cdcfe8ef7da0c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie5f503c91ddf6eff2b9645e6e3c22b2e ;

Ic9c2f173881d25f8976d723957809f51 I13229e09321219c7a9d179fefd0ef804 (
.fgallag_sel( I4d6c95605595942a34573d6ed55eb326[fgallag_SEL-1:0]),
.fgallag( Ieb7e6a2425e93a2b96a94f0e2c4442c3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icec022a0de167257d08e0b2beb6ba8f5 = (I4d6c95605595942a34573d6ed55eb326[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ieb7e6a2425e93a2b96a94f0e2c4442c3 ;

Ic9c2f173881d25f8976d723957809f51 If3f716acc8533596e27e2cc682681416 (
.fgallag_sel( Id6d8f32958dfa1a98958a84e7f1aed02[fgallag_SEL-1:0]),
.fgallag( I4a0483f2d2585cd44fe35191d7cd88b1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3d8a7850f0080b0d6068d58837e3294f = (Id6d8f32958dfa1a98958a84e7f1aed02[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4a0483f2d2585cd44fe35191d7cd88b1 ;

Ic9c2f173881d25f8976d723957809f51 I69246a60a1fc2696f930a33a5c1b0574 (
.fgallag_sel( I971cdf9ddd1bfff5664eec35f22da335[fgallag_SEL-1:0]),
.fgallag( I00e8b3cde14889fcb0b40dc5582a58f9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I26b947511e25e51f1bb9728c169e7e64 = (I971cdf9ddd1bfff5664eec35f22da335[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I00e8b3cde14889fcb0b40dc5582a58f9 ;

Ic9c2f173881d25f8976d723957809f51 I28c5363f71df47cd56c7686a04f10bd5 (
.fgallag_sel( Idd8bc1412a0dc5f489ef253a6164ceea[fgallag_SEL-1:0]),
.fgallag( Ib53dbb62231f729a278d2afa3acffdbf ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8baf26027cc707ae93b6c74e2af5f207 = (Idd8bc1412a0dc5f489ef253a6164ceea[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib53dbb62231f729a278d2afa3acffdbf ;

Ic9c2f173881d25f8976d723957809f51 Id2cc079a08a1b14049749cb27092d191 (
.fgallag_sel( Idbeec36de0128e5924e214877c82bf11[fgallag_SEL-1:0]),
.fgallag( I5503d6011d58dfa4e1ec524eb1875c7d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9902253554855a3d12ceaf47f6cc5569 = (Idbeec36de0128e5924e214877c82bf11[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5503d6011d58dfa4e1ec524eb1875c7d ;

Ic9c2f173881d25f8976d723957809f51 I68cf330449a5a5ced3cb923cc1ebf081 (
.fgallag_sel( I50a9cd240979bc56421bf85011ae99ed[fgallag_SEL-1:0]),
.fgallag( Id86fbda00d923c29c99b4a9fe52d513a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I81ab0ce0526dd851c51d5d42f807e62d = (I50a9cd240979bc56421bf85011ae99ed[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id86fbda00d923c29c99b4a9fe52d513a ;

Ic9c2f173881d25f8976d723957809f51 I6310696939f1fe51cffbabc8755b26fc (
.fgallag_sel( I6437095f6bad2d4fb2fbe0361f60bba1[fgallag_SEL-1:0]),
.fgallag( I3ba6e9f7d7fa98ad776299f8cd8a8363 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I51dc4acb242b33bb123f8b106aafbc93 = (I6437095f6bad2d4fb2fbe0361f60bba1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3ba6e9f7d7fa98ad776299f8cd8a8363 ;

Ic9c2f173881d25f8976d723957809f51 Iffb7519a284c80b34de35c957cfb7e2c (
.fgallag_sel( Ie9b6eb3bbac26635aa00c38110958d46[fgallag_SEL-1:0]),
.fgallag( I67b512efbaf9c063a4ac75cb97a8abdb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I32ca8b2806bf397557167b133d1411ab = (Ie9b6eb3bbac26635aa00c38110958d46[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I67b512efbaf9c063a4ac75cb97a8abdb ;

Ic9c2f173881d25f8976d723957809f51 I7ae7a802452f175b8c02fbdadf26b836 (
.fgallag_sel( I9f34e81e3ffb85539a6273babc2a732e[fgallag_SEL-1:0]),
.fgallag( If5f5eecf512463544c8b2419c0a58779 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5c39fac168568808f33fc6be5eec66a7 = (I9f34e81e3ffb85539a6273babc2a732e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If5f5eecf512463544c8b2419c0a58779 ;

Ic9c2f173881d25f8976d723957809f51 I399966b07ebd7bb6a467eea63d1d6598 (
.fgallag_sel( Id0a1ab8472d704001e0eba0317b117d6[fgallag_SEL-1:0]),
.fgallag( I81cdc8b54bc7f98798713985e8f4553e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If355236b8b8375ad095cc46a373ad4d6 = (Id0a1ab8472d704001e0eba0317b117d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I81cdc8b54bc7f98798713985e8f4553e ;

Ic9c2f173881d25f8976d723957809f51 I51f048123e20c267553de3570304de1e (
.fgallag_sel( I9e632217cd0561d8faa28e4b8850d995[fgallag_SEL-1:0]),
.fgallag( I35bb2eb0cb589f694001ba1509cbf7f8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I31fad95729e24c7724a73285e966684f = (I9e632217cd0561d8faa28e4b8850d995[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I35bb2eb0cb589f694001ba1509cbf7f8 ;

Ic9c2f173881d25f8976d723957809f51 I3c10d515e1f4da9fa0b20c7a9688f620 (
.fgallag_sel( Iedeb5b7b2fa8acf1ea083102678710ea[fgallag_SEL-1:0]),
.fgallag( I3bf8f19c98c78f8e1c315e75a533bb1c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0415d9d3687656d7a07ea2c12ba505d1 = (Iedeb5b7b2fa8acf1ea083102678710ea[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3bf8f19c98c78f8e1c315e75a533bb1c ;

Ic9c2f173881d25f8976d723957809f51 I732371e251d462a3436d999a67a7634f (
.fgallag_sel( I972431d1f5af0bdf4828e4f85591e358[fgallag_SEL-1:0]),
.fgallag( I71cbdcd6e3a873851e9084bc9dcd99bd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id54f584cdc590112180e9000e1d015a1 = (I972431d1f5af0bdf4828e4f85591e358[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I71cbdcd6e3a873851e9084bc9dcd99bd ;

Ic9c2f173881d25f8976d723957809f51 Ibfc30160405bd81b86e2a8f2df2ec2be (
.fgallag_sel( I1f41024b715d8312944ccbf70e95bb40[fgallag_SEL-1:0]),
.fgallag( Iebad2e3d84bae3d4807badae823aec52 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If9930e999d72a139c345aeb1c33e51c1 = (I1f41024b715d8312944ccbf70e95bb40[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iebad2e3d84bae3d4807badae823aec52 ;

Ic9c2f173881d25f8976d723957809f51 I56ba239c2adc0054c6f24c72b7164068 (
.fgallag_sel( Ia6bb5ca05f5d0af452c994dd50004e1d[fgallag_SEL-1:0]),
.fgallag( I054f07cdf6a44100034c7e2fb438055f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I28e9624edb8f59290eba51c87f2a88cc = (Ia6bb5ca05f5d0af452c994dd50004e1d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I054f07cdf6a44100034c7e2fb438055f ;

Ic9c2f173881d25f8976d723957809f51 If61bd1ac3e28e35ef68714e50bc2920d (
.fgallag_sel( I9a1d1d1c862808f9a769cbdb3bc634e1[fgallag_SEL-1:0]),
.fgallag( If3b82307d1ad78e262f76ba9b711e1a6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie6c99d8fe1a105832500bf8a722c82c7 = (I9a1d1d1c862808f9a769cbdb3bc634e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If3b82307d1ad78e262f76ba9b711e1a6 ;

Ic9c2f173881d25f8976d723957809f51 I4acf41a29f10e01fb1214cd2afcfd86e (
.fgallag_sel( I9734eb86f4e73ba217739baf5cb1b13c[fgallag_SEL-1:0]),
.fgallag( I0f40c8301521c136b3ede2cc9e8352a3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I24307c47884babba3b0a16a1791c674f = (I9734eb86f4e73ba217739baf5cb1b13c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0f40c8301521c136b3ede2cc9e8352a3 ;

Ic9c2f173881d25f8976d723957809f51 I797de7c977d812a02a60d3b0bc4cf5a8 (
.fgallag_sel( Ifc0fe00f86569956df72d8a960337e8c[fgallag_SEL-1:0]),
.fgallag( I3615a34cbf1646a7cd0f1da43d62faa5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2951bad4b57a2ad6715844998c491ec7 = (Ifc0fe00f86569956df72d8a960337e8c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3615a34cbf1646a7cd0f1da43d62faa5 ;

Ic9c2f173881d25f8976d723957809f51 Ibaf829d5460fb80e0c3f3de8d85566cf (
.fgallag_sel( I223341a807a1d555f759632f67815159[fgallag_SEL-1:0]),
.fgallag( I0bbd697ad8d3877570ab9e200e66164a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie0149abcf22aeff58be4cb418f477239 = (I223341a807a1d555f759632f67815159[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0bbd697ad8d3877570ab9e200e66164a ;

Ic9c2f173881d25f8976d723957809f51 I64ef815a1f17e49adff40f6db6519c33 (
.fgallag_sel( I6c1f5cdf5f2917118941f4af14d67fef[fgallag_SEL-1:0]),
.fgallag( I298f7389a7fd8e927b7e3354f0d32344 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If8ec8dc5888438922c6074ff23eb42c7 = (I6c1f5cdf5f2917118941f4af14d67fef[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I298f7389a7fd8e927b7e3354f0d32344 ;

Ic9c2f173881d25f8976d723957809f51 I72d1764b19886a70ad38dbff9e1ea216 (
.fgallag_sel( Ie84e88fd1aa2a0b90aa1715fcd27a329[fgallag_SEL-1:0]),
.fgallag( I9960d39fce3c5b9945965dedac46dfed ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If969c721b9636b840193a85d8946fc32 = (Ie84e88fd1aa2a0b90aa1715fcd27a329[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9960d39fce3c5b9945965dedac46dfed ;

Ic9c2f173881d25f8976d723957809f51 I10ec0a5da7934dc8736f213d38184fb3 (
.fgallag_sel( I558f70d7039a8bb58d8ea3f72e43dac0[fgallag_SEL-1:0]),
.fgallag( I02f48e93599dc91bb24a144a0ef1a933 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id6dec5f563e485414043770af559ec76 = (I558f70d7039a8bb58d8ea3f72e43dac0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I02f48e93599dc91bb24a144a0ef1a933 ;

Ic9c2f173881d25f8976d723957809f51 Icdfdfd6345b6f635b4d3c38cc193f277 (
.fgallag_sel( I9924269ed3de12f1f2a28893c7f95292[fgallag_SEL-1:0]),
.fgallag( I7e31af1959a0374af6c2767e4837c566 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I79ae237d2105b50c92b8507272bcbd4e = (I9924269ed3de12f1f2a28893c7f95292[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7e31af1959a0374af6c2767e4837c566 ;

Ic9c2f173881d25f8976d723957809f51 I6f34a6fe8ed3d51e2a509889c56f93c8 (
.fgallag_sel( If1153befd1396be2798cc14535ddeb8a[fgallag_SEL-1:0]),
.fgallag( I8d18e2ecaf2bda4a0ba47d9782e9917a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9ea4ebd1f6cea81da598f16b5a7c31f4 = (If1153befd1396be2798cc14535ddeb8a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8d18e2ecaf2bda4a0ba47d9782e9917a ;

Ic9c2f173881d25f8976d723957809f51 I1282506be5bc27e427b17852d68745a6 (
.fgallag_sel( I9bc447b20687fb3e7eff45792bd4dc3a[fgallag_SEL-1:0]),
.fgallag( Id0a13655f967dfd3000b8dcf4a57f555 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id7b8f8df1818623e7a9e897e019a09e7 = (I9bc447b20687fb3e7eff45792bd4dc3a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id0a13655f967dfd3000b8dcf4a57f555 ;

Ic9c2f173881d25f8976d723957809f51 Id0c29936d1efd0200156fc430e489184 (
.fgallag_sel( If590520f01e452db9867a8d6d5dab29b[fgallag_SEL-1:0]),
.fgallag( Ibf384c0b998b5a5f7808c54292c6b844 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia5e1a46c7d21e79ef859b788b27ee3d1 = (If590520f01e452db9867a8d6d5dab29b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibf384c0b998b5a5f7808c54292c6b844 ;

Ic9c2f173881d25f8976d723957809f51 Ica4df665a4d31f49724b730501629167 (
.fgallag_sel( Id93ee7d283016ab9b0aaa21237237c54[fgallag_SEL-1:0]),
.fgallag( I58b8202ae510e96b4f6ae334f3b282c6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If5b0270fa354f64b8b58e5f02353daa4 = (Id93ee7d283016ab9b0aaa21237237c54[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I58b8202ae510e96b4f6ae334f3b282c6 ;

Ic9c2f173881d25f8976d723957809f51 Ia895cbe2c2e8a017267df8cdb1c1fb4f (
.fgallag_sel( Ic1cf03baabaed466fe532e4db3a9ea78[fgallag_SEL-1:0]),
.fgallag( Icbc75d6e4d0bcc42cdf813529b017e0e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie800c32198a9d6181225f2274b301d9d = (Ic1cf03baabaed466fe532e4db3a9ea78[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Icbc75d6e4d0bcc42cdf813529b017e0e ;

Ic9c2f173881d25f8976d723957809f51 Iaa1ce53a9180152b865f3331618e9709 (
.fgallag_sel( If3031f9aa8f6eba90eac12db7839fefd[fgallag_SEL-1:0]),
.fgallag( I6fa1835a8e7f8ea435c4515b1c059cc9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id596782860b623f79a8fd0e83712d9d0 = (If3031f9aa8f6eba90eac12db7839fefd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6fa1835a8e7f8ea435c4515b1c059cc9 ;

Ic9c2f173881d25f8976d723957809f51 Ie93b9eb93e41891f8eee28488389c6c6 (
.fgallag_sel( I0dc2708970ca2b6c092273b6626bacd6[fgallag_SEL-1:0]),
.fgallag( Id3984a3dd1009c9c76347b9843f27b25 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If5a41054200c97e01b9132f7c7ff9793 = (I0dc2708970ca2b6c092273b6626bacd6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id3984a3dd1009c9c76347b9843f27b25 ;

Ic9c2f173881d25f8976d723957809f51 Ic44a6d819cabdabf59becbda5aa34350 (
.fgallag_sel( Ia58944aebf0b4f0a7d76a1444fced9de[fgallag_SEL-1:0]),
.fgallag( Id5fd757abdc0b2e1b1d4c5dab96ee08a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2cf304c8f8efef74593929b1bea0bf91 = (Ia58944aebf0b4f0a7d76a1444fced9de[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id5fd757abdc0b2e1b1d4c5dab96ee08a ;

Ic9c2f173881d25f8976d723957809f51 I8092cf043080b1aa583f2c1a79f30f44 (
.fgallag_sel( Iedd8e69679d10e05f2889f1d71cf0e7b[fgallag_SEL-1:0]),
.fgallag( I98ab1b82b2991b4cb3bec530711bdc43 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id0b597aa1dc456b83d4e38147c97a9fb = (Iedd8e69679d10e05f2889f1d71cf0e7b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I98ab1b82b2991b4cb3bec530711bdc43 ;

Ic9c2f173881d25f8976d723957809f51 I72ca93fa410c42a809e75df860cb45c7 (
.fgallag_sel( I90f0d471914a2333b9dc14d6d01cf927[fgallag_SEL-1:0]),
.fgallag( I610d0ed6f55a4906aac1be5823358392 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I318a691d3ffd634a1c5c362d5b3a8c34 = (I90f0d471914a2333b9dc14d6d01cf927[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I610d0ed6f55a4906aac1be5823358392 ;

Ic9c2f173881d25f8976d723957809f51 I6458958320a561220013f59690af9006 (
.fgallag_sel( Idceeb22013af64b6bb9f0d773e9ffe9a[fgallag_SEL-1:0]),
.fgallag( I2ed0ad73f73f9f4e1b7ec38af320ee4d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I881c34f97e2d2f4765cf3cd7cde53c7f = (Idceeb22013af64b6bb9f0d773e9ffe9a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2ed0ad73f73f9f4e1b7ec38af320ee4d ;

Ic9c2f173881d25f8976d723957809f51 I1655b13a2b5678047612684d7f1642fe (
.fgallag_sel( If43574342e60a625fb6bee5a495e88f3[fgallag_SEL-1:0]),
.fgallag( I3dfc4dd447cd1f4e40506f516c106861 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I922d1ac78df6c82308d2028527f8f56c = (If43574342e60a625fb6bee5a495e88f3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3dfc4dd447cd1f4e40506f516c106861 ;

Ic9c2f173881d25f8976d723957809f51 Ifa65c844fb98d311f174248284c4f2c9 (
.fgallag_sel( Id285f055275014d9f23d35f91879afa1[fgallag_SEL-1:0]),
.fgallag( Idfeea354b3f9ca8c671851fd90f4e1bc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I49dbef91e0572ad9296838e769edf0c3 = (Id285f055275014d9f23d35f91879afa1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idfeea354b3f9ca8c671851fd90f4e1bc ;

Ic9c2f173881d25f8976d723957809f51 I2e12317e20353684478288f40f5d3400 (
.fgallag_sel( I8c803ab08db372802117de4fa4e2a187[fgallag_SEL-1:0]),
.fgallag( I415d8306edb869fc838eb518aad75168 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8819e4519e4930d300f5536af5d62a94 = (I8c803ab08db372802117de4fa4e2a187[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I415d8306edb869fc838eb518aad75168 ;

Ic9c2f173881d25f8976d723957809f51 I6e7572da2ac8d09b70f592948fb3e9cc (
.fgallag_sel( I13ba48a6b360f3cff5f37ce60cb735c6[fgallag_SEL-1:0]),
.fgallag( I1dc6b2aef1bb326c3d5c19f97a2e1d4f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4779a6c85288e6dba977cedd1cd3cb6b = (I13ba48a6b360f3cff5f37ce60cb735c6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1dc6b2aef1bb326c3d5c19f97a2e1d4f ;

Ic9c2f173881d25f8976d723957809f51 Ie45735194031f713dcc2d34007404d27 (
.fgallag_sel( I4547cd1dad45dfd01e335e8cf20eadd6[fgallag_SEL-1:0]),
.fgallag( Ie2f47a06ca4b6d5823cbbe099f5de0f0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I934d36f3afd37afdaad46c93f45a044c = (I4547cd1dad45dfd01e335e8cf20eadd6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie2f47a06ca4b6d5823cbbe099f5de0f0 ;

Ic9c2f173881d25f8976d723957809f51 I58ec0adf008a7749a1e3f0aec6505f41 (
.fgallag_sel( I0a305655b815b0cc159ac1c5f4ce30f8[fgallag_SEL-1:0]),
.fgallag( I55b7a58384e50ade254c3c8934c290f6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2667428380ad21221430252aa00402bf = (I0a305655b815b0cc159ac1c5f4ce30f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I55b7a58384e50ade254c3c8934c290f6 ;

Ic9c2f173881d25f8976d723957809f51 If2705d0889007db162471e119b7c8d2e (
.fgallag_sel( I3633737da6b74284b0ea9a06c3f5875f[fgallag_SEL-1:0]),
.fgallag( I53bf5dca5911aec50866be5a720d4aa2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I257185648f29565e2259890a6a70583a = (I3633737da6b74284b0ea9a06c3f5875f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I53bf5dca5911aec50866be5a720d4aa2 ;

Ic9c2f173881d25f8976d723957809f51 Ie9eb0cd07fc71a4a5b04ef829533c021 (
.fgallag_sel( Ia949c1b338d1cba07cf6bb6572c3e322[fgallag_SEL-1:0]),
.fgallag( Ie57f78d4c002e69e0e92b25bad752d3f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I49a61c916eb52d0bfd08700d087d379a = (Ia949c1b338d1cba07cf6bb6572c3e322[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie57f78d4c002e69e0e92b25bad752d3f ;

Ic9c2f173881d25f8976d723957809f51 If4a3a18ce8b017a6522183e2a0fadbf9 (
.fgallag_sel( I9a0185f8400159415bc0ad6c38284041[fgallag_SEL-1:0]),
.fgallag( I2ac511a908c9973254672fd38cabccd3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If180a1b31f53c672e4f05b2aeca3caba = (I9a0185f8400159415bc0ad6c38284041[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2ac511a908c9973254672fd38cabccd3 ;

Ic9c2f173881d25f8976d723957809f51 I54a58a01f0356124cfc2e8d265d7288b (
.fgallag_sel( I3eeffe43e7deed7ee77a7f5a3bce3cd2[fgallag_SEL-1:0]),
.fgallag( I8f06d78dd2e6be736f4e4f41fadf130d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I335057378d9ae46b1e1442fd341fabad = (I3eeffe43e7deed7ee77a7f5a3bce3cd2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8f06d78dd2e6be736f4e4f41fadf130d ;

Ic9c2f173881d25f8976d723957809f51 I10748b83c097e6c9b160bbe68ce6839e (
.fgallag_sel( I85af0c31ca7002ae569d9f5ce39943f7[fgallag_SEL-1:0]),
.fgallag( I65450e396e33720967b7a6271e3a70e1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3027f4cba09ab3eee29cf9b34ed27ae4 = (I85af0c31ca7002ae569d9f5ce39943f7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I65450e396e33720967b7a6271e3a70e1 ;

Ic9c2f173881d25f8976d723957809f51 I699af38b26169827d819760d675d989a (
.fgallag_sel( I3dfb8d2fad83fbd807fbfc6330c5b857[fgallag_SEL-1:0]),
.fgallag( I876c6361d2164d03cad2ffc8bf920ac0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9ac1c5487994b853d666af93d35c82cc = (I3dfb8d2fad83fbd807fbfc6330c5b857[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I876c6361d2164d03cad2ffc8bf920ac0 ;

Ic9c2f173881d25f8976d723957809f51 I2f23ce24b0b2c5994c478d30d437ffff (
.fgallag_sel( Ic12be21bcba5fa49437cc44dd8a7f064[fgallag_SEL-1:0]),
.fgallag( Id3b8e1157a3e9eea4d210f466740f673 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I099f1e1b4eb55718dd73dff7efc16ae9 = (Ic12be21bcba5fa49437cc44dd8a7f064[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id3b8e1157a3e9eea4d210f466740f673 ;

Ic9c2f173881d25f8976d723957809f51 I41d370caf3dd1684803c304ff1fc9541 (
.fgallag_sel( I713a384d022d3012e3d0019f5c4ac077[fgallag_SEL-1:0]),
.fgallag( I6973de59fb6014d7c4bf5b982cddc4d8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie9ebb06f41fbc042867ee14d8f4090f2 = (I713a384d022d3012e3d0019f5c4ac077[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6973de59fb6014d7c4bf5b982cddc4d8 ;

Ic9c2f173881d25f8976d723957809f51 I49b594b182849355991fb1f245e64197 (
.fgallag_sel( I80550019479d0323d0dd7e7d0f767d83[fgallag_SEL-1:0]),
.fgallag( I26cb99c4cc37be5f52dfeeca60d5d102 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2647305e100a9fb38fbf290f12778d49 = (I80550019479d0323d0dd7e7d0f767d83[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I26cb99c4cc37be5f52dfeeca60d5d102 ;

Ic9c2f173881d25f8976d723957809f51 I0c06eb001db09660d3e6991b41a018e1 (
.fgallag_sel( Ib8a866f080dd997e0b6c93b6c844d1bc[fgallag_SEL-1:0]),
.fgallag( Ie9835b1d512d9c9c4f2801956fbf13cb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iae4b5e5348101abc4640c84686ddad69 = (Ib8a866f080dd997e0b6c93b6c844d1bc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie9835b1d512d9c9c4f2801956fbf13cb ;

Ic9c2f173881d25f8976d723957809f51 I571a230e6fe8a8f0fe37c70cb3b37c7f (
.fgallag_sel( Id542de206d736ee3769ea0bd037cb627[fgallag_SEL-1:0]),
.fgallag( I89057e4e979b903ae1f10f9dd2f196fe ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibeba1d51f76197f960672ea90dabfb75 = (Id542de206d736ee3769ea0bd037cb627[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I89057e4e979b903ae1f10f9dd2f196fe ;

Ic9c2f173881d25f8976d723957809f51 I3a85255c65a60c09fe6c379792ca3cc7 (
.fgallag_sel( I77e6cdb09c92492c3303d0213de9c291[fgallag_SEL-1:0]),
.fgallag( If1299e6b34cd1f2239d64ade23f33f01 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I83ebb6a41c9d866a8ff3fe3fa0b5321f = (I77e6cdb09c92492c3303d0213de9c291[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If1299e6b34cd1f2239d64ade23f33f01 ;

Ic9c2f173881d25f8976d723957809f51 I1dcf8fbf22ec227f2cace6cf4782a1bf (
.fgallag_sel( I788c33a9f94b26f4ce0f515891d06f90[fgallag_SEL-1:0]),
.fgallag( I3f106ef1876021bb3cc5866d2b5698f4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iedc551659ac328435c906b5748c9790f = (I788c33a9f94b26f4ce0f515891d06f90[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3f106ef1876021bb3cc5866d2b5698f4 ;

Ic9c2f173881d25f8976d723957809f51 I1f3d48668704adf4b983c7b518d7013d (
.fgallag_sel( Iaf7074c2b570a296fe2ea8a5a7097ca0[fgallag_SEL-1:0]),
.fgallag( If6cb9fec3dc380f1c4894bccfa35b33c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I95e1540f2a2eadf6fb80e3519a1d9d5c = (Iaf7074c2b570a296fe2ea8a5a7097ca0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If6cb9fec3dc380f1c4894bccfa35b33c ;

Ic9c2f173881d25f8976d723957809f51 I6c6d416f221b844573ca78121bcaff8e (
.fgallag_sel( I8964c6d3f8e02866a6ad86553ab05d99[fgallag_SEL-1:0]),
.fgallag( I313980f8406e9f26d5eaa53270a23b9e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3587e6334c7c3f23bee5675353bbeaba = (I8964c6d3f8e02866a6ad86553ab05d99[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I313980f8406e9f26d5eaa53270a23b9e ;

Ic9c2f173881d25f8976d723957809f51 I358c73fdfa019b0722c6eea408aa2303 (
.fgallag_sel( I2aa25edaca90c9dae8ed63b48d333c17[fgallag_SEL-1:0]),
.fgallag( I792b5aea212da69a9c18f5723e820432 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4e71cbc9773ff4abc24804d39a64abf8 = (I2aa25edaca90c9dae8ed63b48d333c17[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I792b5aea212da69a9c18f5723e820432 ;

Ic9c2f173881d25f8976d723957809f51 I286ce711ac39c767450bec155eabde5c (
.fgallag_sel( I51a440917c7ae23339bec6f8a745c103[fgallag_SEL-1:0]),
.fgallag( I98f245ec9b667dc065c9494c00ecdf88 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I884dc79c03a585814e9d058ef7669ed8 = (I51a440917c7ae23339bec6f8a745c103[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I98f245ec9b667dc065c9494c00ecdf88 ;

Ic9c2f173881d25f8976d723957809f51 I709b4a08ab654b0493ba0a499e9b5cc0 (
.fgallag_sel( I56ce875e4619d4d8d6ca2fa0ddee91b1[fgallag_SEL-1:0]),
.fgallag( I15254b39b6e136520a9497d8684f9d94 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0b2b9b8f1d6c6d5c6c5a8bd883d3ea5c = (I56ce875e4619d4d8d6ca2fa0ddee91b1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I15254b39b6e136520a9497d8684f9d94 ;

Ic9c2f173881d25f8976d723957809f51 Ic9f40fdeaa3fe76bac17d1a73d86fdbb (
.fgallag_sel( I80607da8f92f5a5d2e4798a62a7b1c5c[fgallag_SEL-1:0]),
.fgallag( I6c8312a9d655f143a0b65d91907ce533 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I645a63009d5be827b30fa02df646c872 = (I80607da8f92f5a5d2e4798a62a7b1c5c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6c8312a9d655f143a0b65d91907ce533 ;

Ic9c2f173881d25f8976d723957809f51 I1c4cca7a75e3210e395f405da58b4a2c (
.fgallag_sel( Ic4dcaa520e26bac40b3876f02074f856[fgallag_SEL-1:0]),
.fgallag( Ie6df2f89b05947f6be3b64e3b4f23df3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If4630c847d9890c2b93acbaa6c9bd392 = (Ic4dcaa520e26bac40b3876f02074f856[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie6df2f89b05947f6be3b64e3b4f23df3 ;

Ic9c2f173881d25f8976d723957809f51 I84c869a3b831703f927e4249b074c6fc (
.fgallag_sel( I3b2714d34081a3b6cccc47fa1638e72e[fgallag_SEL-1:0]),
.fgallag( Ia71232b0b468b729fa1262957cbe9faa ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I49c56ae29a27e764325a9dcacb99f907 = (I3b2714d34081a3b6cccc47fa1638e72e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia71232b0b468b729fa1262957cbe9faa ;

Ic9c2f173881d25f8976d723957809f51 I40616fb30c05844cd94cb489af13493c (
.fgallag_sel( I2db1d1ee8f546c00e512875ce2e13cee[fgallag_SEL-1:0]),
.fgallag( If75d8d882c6afc3df62096486b8e5b80 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie5272faa6aabb6e8d0720cdb7ec98358 = (I2db1d1ee8f546c00e512875ce2e13cee[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If75d8d882c6afc3df62096486b8e5b80 ;

Ic9c2f173881d25f8976d723957809f51 Iab3b2f015f705de6906548127d248a31 (
.fgallag_sel( If80a6bb104ff3b2020e909103c104063[fgallag_SEL-1:0]),
.fgallag( I7ed551b891500784c827992eb53f9ef9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I92779ca466dbced9070a774d84439921 = (If80a6bb104ff3b2020e909103c104063[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7ed551b891500784c827992eb53f9ef9 ;

Ic9c2f173881d25f8976d723957809f51 Ic63c09031ec9cc940ae59d68c671fca7 (
.fgallag_sel( Iadb72cc5444816fbd132256493930bb4[fgallag_SEL-1:0]),
.fgallag( I5b5a24fd7116acd8ad2161513848c6a2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I037e8ab38d779544d25ca5a4bfadeade = (Iadb72cc5444816fbd132256493930bb4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5b5a24fd7116acd8ad2161513848c6a2 ;

Ic9c2f173881d25f8976d723957809f51 I505b37e353f9cfbee0354750227eb861 (
.fgallag_sel( I3a8ec1ad07bfada3d2c6ffca88b8b678[fgallag_SEL-1:0]),
.fgallag( Id7055f4e578533dbd25d0505f8e47f34 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3001e26d13b0cca9bc53d24324ac44d4 = (I3a8ec1ad07bfada3d2c6ffca88b8b678[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id7055f4e578533dbd25d0505f8e47f34 ;

Ic9c2f173881d25f8976d723957809f51 Ib8a15e1f561a3e3b672177f83841687b (
.fgallag_sel( I0aa042b86d9f68d22a49b4eb480a9088[fgallag_SEL-1:0]),
.fgallag( I9c78f3a2aa3986718caf8e70d4d939d4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I933465899e56523ce1c470cad8dbd229 = (I0aa042b86d9f68d22a49b4eb480a9088[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9c78f3a2aa3986718caf8e70d4d939d4 ;

Ic9c2f173881d25f8976d723957809f51 Ia3cb95f1bef810d10df8981c546db030 (
.fgallag_sel( I89a387374771b68d87d7ff2dcc810829[fgallag_SEL-1:0]),
.fgallag( I2def789e23f8ea0edee6f58200144096 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id8b135f08d0464f9e308e25b8df2eb1d = (I89a387374771b68d87d7ff2dcc810829[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2def789e23f8ea0edee6f58200144096 ;

Ic9c2f173881d25f8976d723957809f51 I4dfc00b6ef6585c9e750cbcc1ab54936 (
.fgallag_sel( I2935b3d5c3bba4dddfc7ae03fa77b229[fgallag_SEL-1:0]),
.fgallag( I319c2cb3a815a6347511f0c398876a3c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I938596dee81ba14870ee4acfabce5e7b = (I2935b3d5c3bba4dddfc7ae03fa77b229[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I319c2cb3a815a6347511f0c398876a3c ;

Ic9c2f173881d25f8976d723957809f51 I6090f87a806b2f91b4cc4dfd13a87799 (
.fgallag_sel( I4e0c0248f4aa97d263d64dfec36e3aa2[fgallag_SEL-1:0]),
.fgallag( I0603434655e30a66d4e00b2bc2c878c0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I61599f00ae7d6964dd40c96edefd6f67 = (I4e0c0248f4aa97d263d64dfec36e3aa2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0603434655e30a66d4e00b2bc2c878c0 ;

Ic9c2f173881d25f8976d723957809f51 I04d101af8edca0a2207b3dc92a941799 (
.fgallag_sel( Ia2871d7493b2727d2cb2fbab596b7e6a[fgallag_SEL-1:0]),
.fgallag( Ia6f16190b83b661f68a7a217bb356bdc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic847a85de8e8ba2df520b737ea004374 = (Ia2871d7493b2727d2cb2fbab596b7e6a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia6f16190b83b661f68a7a217bb356bdc ;

Ic9c2f173881d25f8976d723957809f51 I6f0b3b19976429feb08fdc13b862383a (
.fgallag_sel( Ie57adae8873946d6c706074b52a49786[fgallag_SEL-1:0]),
.fgallag( I68fc61dbee0900bd66be7c7f5aaf8825 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifb0f088bf5bbf1884e1f27ed9808c273 = (Ie57adae8873946d6c706074b52a49786[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I68fc61dbee0900bd66be7c7f5aaf8825 ;

Ic9c2f173881d25f8976d723957809f51 Idd1840488db271e8ab174cd13a6f75d0 (
.fgallag_sel( If5ac85646e4b339a19af658f01d0a17f[fgallag_SEL-1:0]),
.fgallag( I4ddd7ecf84b4ee4a4b6290f3d362f190 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8705aa11e5ada7ec6e5431292d83fc54 = (If5ac85646e4b339a19af658f01d0a17f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4ddd7ecf84b4ee4a4b6290f3d362f190 ;

Ic9c2f173881d25f8976d723957809f51 I2708f58ef92fd13a8c4208de4e6481a2 (
.fgallag_sel( I1c092426f34be030b3e020f40517b0e1[fgallag_SEL-1:0]),
.fgallag( I8e60b67eb6a187737de2717ebb95cf6c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ieaa7babedd5bfa1c8e1eb50d62ad9682 = (I1c092426f34be030b3e020f40517b0e1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8e60b67eb6a187737de2717ebb95cf6c ;

Ic9c2f173881d25f8976d723957809f51 I16c384056ef91a5199775a3e8ca6393f (
.fgallag_sel( Ic719b72ad271bc7c077067518e6bbb98[fgallag_SEL-1:0]),
.fgallag( I7e17264500cb48d228c20542c40169cb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9eb9f7a6fe5932b574084bb18ce44e78 = (Ic719b72ad271bc7c077067518e6bbb98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7e17264500cb48d228c20542c40169cb ;

Ic9c2f173881d25f8976d723957809f51 Iddaceb076abba584a78455f669757bd4 (
.fgallag_sel( Ib87362230682c88d68a0ba70e25f3c20[fgallag_SEL-1:0]),
.fgallag( I6bddfc7b277ff042899fb2acd5625c5e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic4b80e5673ad931188a2edfa1119e139 = (Ib87362230682c88d68a0ba70e25f3c20[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6bddfc7b277ff042899fb2acd5625c5e ;

Ic9c2f173881d25f8976d723957809f51 I01d6c756f4aafe13ad7748e75f183c93 (
.fgallag_sel( Ifcf097a102f8dc1f912022fed893d222[fgallag_SEL-1:0]),
.fgallag( I6daafbc7b14e2736b2a4e29c5f6fc5ff ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5cdaf1ff24d7fb2bb4411b63a0a4488a = (Ifcf097a102f8dc1f912022fed893d222[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6daafbc7b14e2736b2a4e29c5f6fc5ff ;

Ic9c2f173881d25f8976d723957809f51 Ic8ae1111d27a9e4901fd15642a77fd67 (
.fgallag_sel( I56483ca3fa550dc59bfa347780cfef7b[fgallag_SEL-1:0]),
.fgallag( I29df797d4c3ebd64fb088660bf89e922 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7db6dcc03117fef703f20919a3c2ee89 = (I56483ca3fa550dc59bfa347780cfef7b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I29df797d4c3ebd64fb088660bf89e922 ;

Ic9c2f173881d25f8976d723957809f51 Ib9106c1a678fc1b9b9829cabdea83244 (
.fgallag_sel( I4aa9f61be376458185c3235442c8fda0[fgallag_SEL-1:0]),
.fgallag( I9418cc6766916bf1afc1f8a01feaad4e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3d2a8a166ccade50e320baaa68b40954 = (I4aa9f61be376458185c3235442c8fda0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9418cc6766916bf1afc1f8a01feaad4e ;

Ic9c2f173881d25f8976d723957809f51 I6a7082be9b8f50a7758e5357591e8604 (
.fgallag_sel( Id91fde1007d47258273299de80721390[fgallag_SEL-1:0]),
.fgallag( I90e1a5b43e93c02512a76c5cab15c5ad ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3356737fddf6440f36fde442d29bb860 = (Id91fde1007d47258273299de80721390[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I90e1a5b43e93c02512a76c5cab15c5ad ;

Ic9c2f173881d25f8976d723957809f51 Id22e79a1fb5d3c86b1f93f3cde917799 (
.fgallag_sel( Id58498c34aff2e1216c189b9df88822c[fgallag_SEL-1:0]),
.fgallag( I26977fe4cdb2f9714fae2f12ca4a809b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I13d6fc4a99a3a9989e655c417552fdb1 = (Id58498c34aff2e1216c189b9df88822c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I26977fe4cdb2f9714fae2f12ca4a809b ;

Ic9c2f173881d25f8976d723957809f51 Icd76d0eef001cafc53cf157be58b7246 (
.fgallag_sel( Ib52e0c68caadcf4dd9636a84f5460e53[fgallag_SEL-1:0]),
.fgallag( I59775b68e199902c38d62e28cff01393 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8a508ec5f2c2aaa05b632f422e67394f = (Ib52e0c68caadcf4dd9636a84f5460e53[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I59775b68e199902c38d62e28cff01393 ;

Ic9c2f173881d25f8976d723957809f51 I510935920615ecb5a4a8c098cef7f089 (
.fgallag_sel( Ie19679053b289bb5a0aad570cc81bd14[fgallag_SEL-1:0]),
.fgallag( I9470ef82dad13754d8d061b5fd00a667 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I451fd82336efc778a51debf10f7cf325 = (Ie19679053b289bb5a0aad570cc81bd14[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9470ef82dad13754d8d061b5fd00a667 ;

Ic9c2f173881d25f8976d723957809f51 Icf2ff70eb60a57de80df87cb50f9e633 (
.fgallag_sel( I8862c5ef45b723c9abf5d0ab6854a900[fgallag_SEL-1:0]),
.fgallag( I62eb7a176351be84d086ce3c463214e8 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I76637de9be7c2c0dd0c324b4327a6184 = (I8862c5ef45b723c9abf5d0ab6854a900[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I62eb7a176351be84d086ce3c463214e8 ;

Ic9c2f173881d25f8976d723957809f51 I1f7453d914c019158d04a4325f1b7a22 (
.fgallag_sel( I30db951a07af96a8ddf59360141b9a6a[fgallag_SEL-1:0]),
.fgallag( I106eb0d8f9ea92cda7bec4fe4aed6409 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6e6d24ccb985ade6f058ce459592dfb0 = (I30db951a07af96a8ddf59360141b9a6a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I106eb0d8f9ea92cda7bec4fe4aed6409 ;

Ic9c2f173881d25f8976d723957809f51 I620a8a348cfee9072c6eb17223bf47cc (
.fgallag_sel( I4855a0a0c6426d33014ce6a4c96965ce[fgallag_SEL-1:0]),
.fgallag( Id0c12bc1a2139e57ea40c3254f30de7b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If379a7696fdd0afebcb8ca169bb8f34a = (I4855a0a0c6426d33014ce6a4c96965ce[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id0c12bc1a2139e57ea40c3254f30de7b ;

Ic9c2f173881d25f8976d723957809f51 Id3f5457f9b246f05a41d4a60d20dcb47 (
.fgallag_sel( I362e8db1791718290bd33a79b4fc0855[fgallag_SEL-1:0]),
.fgallag( Ib809a6099992799ce0235f22ce798c9a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idbd1062a6090858034185f1d5d503adf = (I362e8db1791718290bd33a79b4fc0855[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib809a6099992799ce0235f22ce798c9a ;

Ic9c2f173881d25f8976d723957809f51 I2eaca010067c4a853ee9290425265eae (
.fgallag_sel( I773f0508440fb71d73fd82a372cc0a00[fgallag_SEL-1:0]),
.fgallag( I1a9be3897e044e9b24ac330ef3a20419 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iea3c638b692d2540c1c8c81a6308673d = (I773f0508440fb71d73fd82a372cc0a00[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1a9be3897e044e9b24ac330ef3a20419 ;

Ic9c2f173881d25f8976d723957809f51 I3902718ac6db47e234ce9700441801c1 (
.fgallag_sel( I792891cecae468d7a87e12f2da62a718[fgallag_SEL-1:0]),
.fgallag( I6e87b3400b7ddab94faf11c3910fa534 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icd9e1d048d56d5d8557f80329bc6ffcc = (I792891cecae468d7a87e12f2da62a718[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6e87b3400b7ddab94faf11c3910fa534 ;

Ic9c2f173881d25f8976d723957809f51 Idd04b3258e1b5f9c6ccd1d29ce7d6180 (
.fgallag_sel( I33303820ad094d7a0ab53bca722fc609[fgallag_SEL-1:0]),
.fgallag( I51e0ff0f52ca609663781545174b763d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6f0de2d570fa0245666c834b823e545b = (I33303820ad094d7a0ab53bca722fc609[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I51e0ff0f52ca609663781545174b763d ;

Ic9c2f173881d25f8976d723957809f51 I1944c42bb915dc71bf7c2d6a95564332 (
.fgallag_sel( Iff98739de575e25104c0dc30f08912a5[fgallag_SEL-1:0]),
.fgallag( I5c523df1fb2161ab4efd1c9b3e6b7aef ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ief41e2502056d029a0c8bea8c052700c = (Iff98739de575e25104c0dc30f08912a5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5c523df1fb2161ab4efd1c9b3e6b7aef ;

Ic9c2f173881d25f8976d723957809f51 Ic7988087e6f2bece4415f3e2c989b3a6 (
.fgallag_sel( I1952614b64ea451e9d0646dcce5dd1cd[fgallag_SEL-1:0]),
.fgallag( Ia307e5901694783f7761cdf724b767d0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7cd5df0d2845c7ed9f336a7940c7256e = (I1952614b64ea451e9d0646dcce5dd1cd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia307e5901694783f7761cdf724b767d0 ;

Ic9c2f173881d25f8976d723957809f51 I599ddd152d17afff0bad8b0d29bd9108 (
.fgallag_sel( I49c1a7d1c20a25496821ad80c7eff790[fgallag_SEL-1:0]),
.fgallag( Ia47164e8ba831b85e696e30ff59ceab1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5471bcc8bf4f4d0fab46d549b43113ef = (I49c1a7d1c20a25496821ad80c7eff790[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia47164e8ba831b85e696e30ff59ceab1 ;

Ic9c2f173881d25f8976d723957809f51 Ibcf651f8df3cf78743f39d7be7214a8c (
.fgallag_sel( Ie2be17a55e79ca76350e033f227800de[fgallag_SEL-1:0]),
.fgallag( Ic217af0cb9728801034fdcb273a577fc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I599b8e0677efc1541283c2d7bf84809f = (Ie2be17a55e79ca76350e033f227800de[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic217af0cb9728801034fdcb273a577fc ;

Ic9c2f173881d25f8976d723957809f51 I4a4287dab4fb632c05278dab5ef93c28 (
.fgallag_sel( I737a5b06f848cacf0c8da4985c73c66b[fgallag_SEL-1:0]),
.fgallag( Id5c8ea61025914f6e5a9b5eab9269261 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4e4829b24a42e96e5c8399156aa61786 = (I737a5b06f848cacf0c8da4985c73c66b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id5c8ea61025914f6e5a9b5eab9269261 ;

Ic9c2f173881d25f8976d723957809f51 I94fa40e833e09dc4a711b7a4894dbbe3 (
.fgallag_sel( Iab160609bb21501aa55b662d2010357b[fgallag_SEL-1:0]),
.fgallag( I924ef8499a83579e3449bbac0994775e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1cda8d902f71f780775c85f38f9e799e = (Iab160609bb21501aa55b662d2010357b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I924ef8499a83579e3449bbac0994775e ;

Ic9c2f173881d25f8976d723957809f51 Ia9cbceaf4e13cd3122bcf0d3ee99e0d0 (
.fgallag_sel( Ief74f1a9d4a43ee5c9def7b83369bb21[fgallag_SEL-1:0]),
.fgallag( Ia8da4833c93e9ef6188709e7082092de ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic0b2c3e49d55853bc705021e5c0a2b06 = (Ief74f1a9d4a43ee5c9def7b83369bb21[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia8da4833c93e9ef6188709e7082092de ;

Ic9c2f173881d25f8976d723957809f51 I7f70a8d18281c7c1acffa18669e134cd (
.fgallag_sel( Id144423f50751e661db3860a8487d004[fgallag_SEL-1:0]),
.fgallag( Icd8516e6bf231bce29ebefbc7c97bff7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6235ba2f129cfbcff36b368a39312bd7 = (Id144423f50751e661db3860a8487d004[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Icd8516e6bf231bce29ebefbc7c97bff7 ;

Ic9c2f173881d25f8976d723957809f51 Id0999532bede9fce3e12ef52e3ba608b (
.fgallag_sel( I623352a4f6705b21d461d6b32e85c12b[fgallag_SEL-1:0]),
.fgallag( I76c6762c515d0c9de1d777c0868b20af ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6804a691f5de298ab553ee66c3e9610c = (I623352a4f6705b21d461d6b32e85c12b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I76c6762c515d0c9de1d777c0868b20af ;

Ic9c2f173881d25f8976d723957809f51 Ib4537744b241a8d73272690a47c98789 (
.fgallag_sel( I28d1dc8dc594977b5058b5bb9f6bfc66[fgallag_SEL-1:0]),
.fgallag( If5da296bcf91d370f8341fc402eed6df ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I973825f628679f8bbaf0650136e7259b = (I28d1dc8dc594977b5058b5bb9f6bfc66[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If5da296bcf91d370f8341fc402eed6df ;

Ic9c2f173881d25f8976d723957809f51 I0d709f9957d11cd5e8381f666f45c7d5 (
.fgallag_sel( I5371a83bf9d6f334cf8d1c5b082527e9[fgallag_SEL-1:0]),
.fgallag( I64673b4b013682f9ce54925853c06ca4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibfa3babbd7909dfada58a7f579281b8c = (I5371a83bf9d6f334cf8d1c5b082527e9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I64673b4b013682f9ce54925853c06ca4 ;

Ic9c2f173881d25f8976d723957809f51 Id43872f1a59191d4f673c93263fdd384 (
.fgallag_sel( If1605d6646fd267e701668a7245b3b44[fgallag_SEL-1:0]),
.fgallag( Iabfccf7b60f9be4e3714ad753cd8922a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0aa6569579526ac14e0d55caa4cef2a7 = (If1605d6646fd267e701668a7245b3b44[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iabfccf7b60f9be4e3714ad753cd8922a ;

Ic9c2f173881d25f8976d723957809f51 I89ccfeda71dbfd799a31c8a03f729136 (
.fgallag_sel( Idf5eb1ac2c5bd92fa08ed935ae298255[fgallag_SEL-1:0]),
.fgallag( I73ab1f85232818929b1b2e9d343584a3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I87c99b1e08ca19dea7ffbfa15ecc2db9 = (Idf5eb1ac2c5bd92fa08ed935ae298255[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I73ab1f85232818929b1b2e9d343584a3 ;

Ic9c2f173881d25f8976d723957809f51 Id537e736da638ec2d96503d9bdccd750 (
.fgallag_sel( I44ce30330c4d2d6033a0a970dd2bdd68[fgallag_SEL-1:0]),
.fgallag( I06f989f65e614903ffba3594e8112235 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I40ba1533f32b981c4e937b2e48f38ea0 = (I44ce30330c4d2d6033a0a970dd2bdd68[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I06f989f65e614903ffba3594e8112235 ;

Ic9c2f173881d25f8976d723957809f51 I75fae94751eb53fdadbd7315a342ba33 (
.fgallag_sel( Ic101b8f56ea1e25c6b752583a1b01242[fgallag_SEL-1:0]),
.fgallag( I0391247480cb6bd6bda2c59dcf8f7607 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I83483243e11dd867b1eea10b6ef0dbd2 = (Ic101b8f56ea1e25c6b752583a1b01242[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0391247480cb6bd6bda2c59dcf8f7607 ;

Ic9c2f173881d25f8976d723957809f51 I73fb1489837099d536418e33ab049dc3 (
.fgallag_sel( Ib7cf44e681881e55d2d353280a6319d6[fgallag_SEL-1:0]),
.fgallag( Iee114a92d2238e4b8fcdfa79c4c99d6a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8265d9994495dbe871b565be6710b428 = (Ib7cf44e681881e55d2d353280a6319d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iee114a92d2238e4b8fcdfa79c4c99d6a ;

Ic9c2f173881d25f8976d723957809f51 I7e8af7d5cbc961cf91c973279881b474 (
.fgallag_sel( I35690f724e964248dbb1e80fb1ea49f8[fgallag_SEL-1:0]),
.fgallag( Ida429b8e252b80b45435af1c6522f783 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3d4ee0ad8461c2ac5128adc9c231f465 = (I35690f724e964248dbb1e80fb1ea49f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ida429b8e252b80b45435af1c6522f783 ;

Ic9c2f173881d25f8976d723957809f51 I558b57199e5e1044b10136f4be3bd2f9 (
.fgallag_sel( I5affa2759148a6baf5b9f0cd3122348c[fgallag_SEL-1:0]),
.fgallag( Id3849d43e39d78fd2428109bf9677e0d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib609900664dc10ef97873cccb161c320 = (I5affa2759148a6baf5b9f0cd3122348c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id3849d43e39d78fd2428109bf9677e0d ;

Ic9c2f173881d25f8976d723957809f51 I3e05ab9ef97382c792226fcba43e35ae (
.fgallag_sel( Iaeea1f06ff0c6e9cfa43ba14420c3adc[fgallag_SEL-1:0]),
.fgallag( I5e51799e585f3dbef5e64908bcfc3e7a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If8b44d90a4ef1715e9144255d606a27e = (Iaeea1f06ff0c6e9cfa43ba14420c3adc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5e51799e585f3dbef5e64908bcfc3e7a ;

Ic9c2f173881d25f8976d723957809f51 I8384fe686d2fbeb6911ae3ec3ed4db87 (
.fgallag_sel( Iac5a23266c3b038b4b54a916dccdf3a8[fgallag_SEL-1:0]),
.fgallag( I6d12e4545b8befb8d09545ea00c8ea96 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I06715db3159c94a5913c05e9827cddd1 = (Iac5a23266c3b038b4b54a916dccdf3a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6d12e4545b8befb8d09545ea00c8ea96 ;

Ic9c2f173881d25f8976d723957809f51 If06073d8fd7050d37d23dda31b8fb14f (
.fgallag_sel( Icdfb7f52cc27b1cfcde90a100d29af13[fgallag_SEL-1:0]),
.fgallag( I98d04e6bae91796784a864c5bed637cb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia295ba836438cd4e7c1b03b4261949ed = (Icdfb7f52cc27b1cfcde90a100d29af13[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I98d04e6bae91796784a864c5bed637cb ;

Ic9c2f173881d25f8976d723957809f51 I3ceb4032cc7e18993dd228850e65d119 (
.fgallag_sel( I71484d7e00efa02a08b54a1405f2902c[fgallag_SEL-1:0]),
.fgallag( I83b3247bed67d1e2ed488d5b7812851d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5f9c502cdffe77bb7e298a9bfdd325b1 = (I71484d7e00efa02a08b54a1405f2902c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I83b3247bed67d1e2ed488d5b7812851d ;

Ic9c2f173881d25f8976d723957809f51 I00d8590a5195956af795376c91f1a381 (
.fgallag_sel( I68a9b0607e69e8b3dae64689eb288a33[fgallag_SEL-1:0]),
.fgallag( I868021f44830a9d81c4ba3dad804f889 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3f13e4887f4982583fe615807c42d121 = (I68a9b0607e69e8b3dae64689eb288a33[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I868021f44830a9d81c4ba3dad804f889 ;

Ic9c2f173881d25f8976d723957809f51 Id3bdb11d564326449ba4eddad1254134 (
.fgallag_sel( I2598c48aad48072a7f216b2ab56ee532[fgallag_SEL-1:0]),
.fgallag( I685e59e3865058f29978a8cc2f1b6c7c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie1a491c10dad8dfd4b0fe42977d625b6 = (I2598c48aad48072a7f216b2ab56ee532[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I685e59e3865058f29978a8cc2f1b6c7c ;

Ic9c2f173881d25f8976d723957809f51 I993ea1e9de62d8edd5124dae5f019758 (
.fgallag_sel( I796e3a193b1b66fa9a04ca60aee11ea1[fgallag_SEL-1:0]),
.fgallag( I5a76dd9f4a2078dee81102a9f205ca53 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id2334d193c70ad43e5b7cdcd923e364a = (I796e3a193b1b66fa9a04ca60aee11ea1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5a76dd9f4a2078dee81102a9f205ca53 ;

Ic9c2f173881d25f8976d723957809f51 Ib7e3526ef4c618e2f966fa48822ed800 (
.fgallag_sel( Ic96be7e69faf0f43b92618131cf0c98a[fgallag_SEL-1:0]),
.fgallag( Ice3bd7a4bbf0705a3dc1f89c5ceca084 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I621999a98b66cc50cf7732668af444e0 = (Ic96be7e69faf0f43b92618131cf0c98a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ice3bd7a4bbf0705a3dc1f89c5ceca084 ;

Ic9c2f173881d25f8976d723957809f51 Ic95efcba247a69eedc0bdb007ccb8f98 (
.fgallag_sel( I648afe4114ce435bf1d13e0ad54425cf[fgallag_SEL-1:0]),
.fgallag( I5f741a3213cecdf58440120c2ea78e87 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8c5fe32c1860a2beb9c14634c62a95aa = (I648afe4114ce435bf1d13e0ad54425cf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5f741a3213cecdf58440120c2ea78e87 ;

Ic9c2f173881d25f8976d723957809f51 I7aa67413dda82b41698253c375ed7609 (
.fgallag_sel( If05d7e30b4717e0a1bfd20b90d0539bd[fgallag_SEL-1:0]),
.fgallag( Idad89ade7f96091abfea876b3af0d5b4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5cc33aeefc2bbf0d777b4b59bcba7ec4 = (If05d7e30b4717e0a1bfd20b90d0539bd[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idad89ade7f96091abfea876b3af0d5b4 ;

Ic9c2f173881d25f8976d723957809f51 I46c8308b812c7eb242bc2442b1772e30 (
.fgallag_sel( I5fc356af8a62a1d739cb375fb851e90f[fgallag_SEL-1:0]),
.fgallag( Ie0ab4b7c79196195db0971e7c7a85adb ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5a2f74df4050f2898061471586f3fb63 = (I5fc356af8a62a1d739cb375fb851e90f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie0ab4b7c79196195db0971e7c7a85adb ;

Ic9c2f173881d25f8976d723957809f51 I242a7ea3c0be277aa8bc2656f0da14a4 (
.fgallag_sel( I22f4c5403fbe33d18f97cf21786cdd80[fgallag_SEL-1:0]),
.fgallag( I0093585d710940feaa8ebdc5fb000806 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I54c68d66f2692522fdd982a31ff0b3a8 = (I22f4c5403fbe33d18f97cf21786cdd80[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0093585d710940feaa8ebdc5fb000806 ;

Ic9c2f173881d25f8976d723957809f51 If986be5291767e6dfe5052c9e18368b2 (
.fgallag_sel( I9a1b2b9f924099f1e57fa501ba2e33ba[fgallag_SEL-1:0]),
.fgallag( I76a0b74bb633743ac56cf4a0d52f80c0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I98b0bc583105e551a5c1c7a8b6de61e1 = (I9a1b2b9f924099f1e57fa501ba2e33ba[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I76a0b74bb633743ac56cf4a0d52f80c0 ;

Ic9c2f173881d25f8976d723957809f51 I8ae501a70118506340bd05253f4c55e1 (
.fgallag_sel( If6253af4ebc430e4937269a5f4989b29[fgallag_SEL-1:0]),
.fgallag( I11931fd13219c1ae615d164a8f4130f9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3ca304e8b6c5440935c6944b64ddde65 = (If6253af4ebc430e4937269a5f4989b29[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I11931fd13219c1ae615d164a8f4130f9 ;

Ic9c2f173881d25f8976d723957809f51 Ic0f4425bc017a531980fc4b84c9ece99 (
.fgallag_sel( I0427d17423548dbb33cf792883b4be8c[fgallag_SEL-1:0]),
.fgallag( I6de7a344ae1574e551c7c10a1773d880 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I33c7b994472de0942347e9b06ed9f59c = (I0427d17423548dbb33cf792883b4be8c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6de7a344ae1574e551c7c10a1773d880 ;

Ic9c2f173881d25f8976d723957809f51 I6eb3466f656864350dd5d0c45b4e8544 (
.fgallag_sel( Ie539faf01ae85253e399308fef98afd6[fgallag_SEL-1:0]),
.fgallag( I4920b0740cb56988ba4fc10b86195cdd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id5395616ea942f63477bffe5c17560e3 = (Ie539faf01ae85253e399308fef98afd6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4920b0740cb56988ba4fc10b86195cdd ;

Ic9c2f173881d25f8976d723957809f51 Icdea5aa4feee7a36ebf3f5b7ef913b69 (
.fgallag_sel( Iae6e7c42f250cd9223f18f8830fb177d[fgallag_SEL-1:0]),
.fgallag( I37d27fda03770ad37a1fbad835c076c3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If90e3127bcb3ed51a225ce72afb0a793 = (Iae6e7c42f250cd9223f18f8830fb177d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I37d27fda03770ad37a1fbad835c076c3 ;

Ic9c2f173881d25f8976d723957809f51 I0f1e8b13dca3874c77169a917560481f (
.fgallag_sel( Iff47ec1743b59d7f90e9042af7ce44cb[fgallag_SEL-1:0]),
.fgallag( Ib868fcb71300c09a49719e0b0459ca06 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia6ff80807e320ef75fbdad7c86add89d = (Iff47ec1743b59d7f90e9042af7ce44cb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib868fcb71300c09a49719e0b0459ca06 ;

Ic9c2f173881d25f8976d723957809f51 I67f40c7f4ae4bc02db3592f9e145dc95 (
.fgallag_sel( I1cf4a55ebab332defa32d2922b885285[fgallag_SEL-1:0]),
.fgallag( I2c67e89b58d7f998c43c68d857fa2381 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If8a6eb502f55f58090ffd901b27086c2 = (I1cf4a55ebab332defa32d2922b885285[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2c67e89b58d7f998c43c68d857fa2381 ;

Ic9c2f173881d25f8976d723957809f51 I542df8a53caf77a72557ec959532c0a3 (
.fgallag_sel( I284913858691ad5724073b73a820047a[fgallag_SEL-1:0]),
.fgallag( Idb770d9fc630f77beca27c3182279001 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If10a93a95dd1f3e7117e64ae2915bcd5 = (I284913858691ad5724073b73a820047a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idb770d9fc630f77beca27c3182279001 ;

Ic9c2f173881d25f8976d723957809f51 Ie3757c301a45e6b57e3e1ee5eb9c7638 (
.fgallag_sel( I35626ca53adbbf0a3a71cc6fcf43bcb1[fgallag_SEL-1:0]),
.fgallag( I6ab74c183d97a5df7a336c6c66c66e2e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id86eeb13a357d077460584e1941e74a7 = (I35626ca53adbbf0a3a71cc6fcf43bcb1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6ab74c183d97a5df7a336c6c66c66e2e ;

Ic9c2f173881d25f8976d723957809f51 I4360aa193a2a1845707a71a49e3e0ad0 (
.fgallag_sel( I0d74ef22d31abcec73c7c582310b1e6d[fgallag_SEL-1:0]),
.fgallag( Ic4fc6d6a69dccb796d208aba87ec002c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5d7e70c0e768f5868bf9fa07111036e7 = (I0d74ef22d31abcec73c7c582310b1e6d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic4fc6d6a69dccb796d208aba87ec002c ;

Ic9c2f173881d25f8976d723957809f51 I5ab4a5cfd310d07f1857eea12cf25fcb (
.fgallag_sel( I15f4cf1aa0ad5ce2bda52df338e677e3[fgallag_SEL-1:0]),
.fgallag( I450cd05f0109ad62ae4ca7f540ac7505 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I48f780aaedbd67e6342d9e0232635ac8 = (I15f4cf1aa0ad5ce2bda52df338e677e3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I450cd05f0109ad62ae4ca7f540ac7505 ;

Ic9c2f173881d25f8976d723957809f51 Id5cd920a43f37c4fb9d878da3311e4b4 (
.fgallag_sel( I6c5ca5e68c8844bb1617a2288b5bbc37[fgallag_SEL-1:0]),
.fgallag( Ia6f1bdee90a01ee3f3e59eec00689d50 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia9a47dd6aa0313a806147f2c4a91df0b = (I6c5ca5e68c8844bb1617a2288b5bbc37[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia6f1bdee90a01ee3f3e59eec00689d50 ;

Ic9c2f173881d25f8976d723957809f51 Iad85a44693e128c44e42161bff51f9c2 (
.fgallag_sel( I44343a9491069c3c8ea4fbd6255a5a6c[fgallag_SEL-1:0]),
.fgallag( I33193403a8d72dcd02e87ae03b668e09 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id0a9c8069c91546ee6dcdcca1dbddd61 = (I44343a9491069c3c8ea4fbd6255a5a6c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I33193403a8d72dcd02e87ae03b668e09 ;

Ic9c2f173881d25f8976d723957809f51 I5cc3fa29daa1c95948fc1f1e62d829d6 (
.fgallag_sel( I1d8318b94d86e1fd28323a5e5684a37b[fgallag_SEL-1:0]),
.fgallag( I5208f3202b32a30c4abaca4c617d3b3b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3e30cc2747c9a7dd9c4fcd144f640552 = (I1d8318b94d86e1fd28323a5e5684a37b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5208f3202b32a30c4abaca4c617d3b3b ;

Ic9c2f173881d25f8976d723957809f51 I638fbbd9b1e7705cb12fbd5f090a66e1 (
.fgallag_sel( I825e83bd88575868f4fcc9a8b8729663[fgallag_SEL-1:0]),
.fgallag( Ib607167c806dd831aaed4a42b9cf4349 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia4433ae2b484d7bfff269cb336831628 = (I825e83bd88575868f4fcc9a8b8729663[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib607167c806dd831aaed4a42b9cf4349 ;

Ic9c2f173881d25f8976d723957809f51 Ic013e6787c92269fdec37a1e89bf977a (
.fgallag_sel( I3184a16c71cff80c8c90b40e45f114b8[fgallag_SEL-1:0]),
.fgallag( I42b87e52c168abb775c1e1e5ddfc1958 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7aef236fed5567b77c8a3f5c22e3bff3 = (I3184a16c71cff80c8c90b40e45f114b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I42b87e52c168abb775c1e1e5ddfc1958 ;

Ic9c2f173881d25f8976d723957809f51 Ia423392d98ec42ff08c1c54ac992c9c6 (
.fgallag_sel( Iae133550f8bad8357a73e7de1372faa3[fgallag_SEL-1:0]),
.fgallag( Ifc4e50801a1606717efd57bd5ac6f41f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iff3859ddd94ff25ba5a08a367baf602b = (Iae133550f8bad8357a73e7de1372faa3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifc4e50801a1606717efd57bd5ac6f41f ;

Ic9c2f173881d25f8976d723957809f51 Idca921760380e112e9eacfe8ad3576d3 (
.fgallag_sel( Ibccb4a43c410f698e0fff68553326a77[fgallag_SEL-1:0]),
.fgallag( I5e7282e9a35cead2f4d1d9860d45852c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4c0c110a6f362969bce6db69cb1c0bfc = (Ibccb4a43c410f698e0fff68553326a77[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5e7282e9a35cead2f4d1d9860d45852c ;

Ic9c2f173881d25f8976d723957809f51 Ib14e467f2d8f26417f8de35834f59764 (
.fgallag_sel( I72dc7aa294a3af89101ea62a4223170e[fgallag_SEL-1:0]),
.fgallag( I8503b90594f3d4b492cca9cf154fc3d3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I51225282195bed9916ae55ae7887c1d2 = (I72dc7aa294a3af89101ea62a4223170e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I8503b90594f3d4b492cca9cf154fc3d3 ;

Ic9c2f173881d25f8976d723957809f51 I2091bf71229d2522e513073498f2742d (
.fgallag_sel( I91eb3e70921e0b141a344bc57dfbc934[fgallag_SEL-1:0]),
.fgallag( I95010cdf08c373916ab02e3794afa77a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I58380b8eb6332c81366215b1dd60cea5 = (I91eb3e70921e0b141a344bc57dfbc934[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I95010cdf08c373916ab02e3794afa77a ;

Ic9c2f173881d25f8976d723957809f51 I1def8e7b129515d2d9d8db8033630810 (
.fgallag_sel( I1986f22f2269cc135c6ed28d35fb0bd1[fgallag_SEL-1:0]),
.fgallag( I832fdc71e665ad2acac2576188e0d65b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I55df86c0751564116c4f1a65de2ac9fa = (I1986f22f2269cc135c6ed28d35fb0bd1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I832fdc71e665ad2acac2576188e0d65b ;

Ic9c2f173881d25f8976d723957809f51 I5be00e1a7e227309c0f9d5d2e38354f1 (
.fgallag_sel( Ibef24017bc71de9c002aafa7ce9a784c[fgallag_SEL-1:0]),
.fgallag( Ic21a6f1abcecf14acaf2aa23b7dcdb6b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0bc0390d7c9b369ebc92e9547b87b9df = (Ibef24017bc71de9c002aafa7ce9a784c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic21a6f1abcecf14acaf2aa23b7dcdb6b ;

Ic9c2f173881d25f8976d723957809f51 I5c042480a9a07232c1fe8121400909b0 (
.fgallag_sel( Ieae3ed78fa2c45507066f4e20d96e956[fgallag_SEL-1:0]),
.fgallag( I49847c8c979d9ed82be80f62552e97bf ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icfe3de1a8dc46c883a65345392921c50 = (Ieae3ed78fa2c45507066f4e20d96e956[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I49847c8c979d9ed82be80f62552e97bf ;

Ic9c2f173881d25f8976d723957809f51 Id4f7280f983b15241a0d3b45fa6343a8 (
.fgallag_sel( I730fd25ffc7778fd4bb02d33cb3870d6[fgallag_SEL-1:0]),
.fgallag( I7a2bfe5efbe1d0dc222bff675c621485 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4c0e5a2ba1c2b42970f41699d5ddcb9a = (I730fd25ffc7778fd4bb02d33cb3870d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7a2bfe5efbe1d0dc222bff675c621485 ;

Ic9c2f173881d25f8976d723957809f51 Ic481b87b83ebc908134c69bfcdfdce20 (
.fgallag_sel( I9a32313f2911b797fb0848f7d97e62b9[fgallag_SEL-1:0]),
.fgallag( Ie0d874ce4b0713de7d087396a1879c54 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib81161d68b741b2656196d7284209d58 = (I9a32313f2911b797fb0848f7d97e62b9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie0d874ce4b0713de7d087396a1879c54 ;

Ic9c2f173881d25f8976d723957809f51 I82b04b98f5c24aed5e76bce1f3b8bc9b (
.fgallag_sel( I6373e2d64fdb5dd77733b3e4bb405121[fgallag_SEL-1:0]),
.fgallag( Iaf4c12394552f42e476b70f6c75003d7 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib98bf53c446dcc7920b842d29191fe0a = (I6373e2d64fdb5dd77733b3e4bb405121[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaf4c12394552f42e476b70f6c75003d7 ;

Ic9c2f173881d25f8976d723957809f51 I6134adccaaa6acaebbf26b9c4f575a9d (
.fgallag_sel( Ib437aa67ab7c13b45d7a4d56ce9e79b8[fgallag_SEL-1:0]),
.fgallag( I64d7f4a0df87ce07ce49350610122f79 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I31c34cf26a3890305171a6beca791fa3 = (Ib437aa67ab7c13b45d7a4d56ce9e79b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I64d7f4a0df87ce07ce49350610122f79 ;

Ic9c2f173881d25f8976d723957809f51 I92378486628266460af4c20f5f2a7b97 (
.fgallag_sel( I0cb5c7a759f4c75d4a675f9777f15c5f[fgallag_SEL-1:0]),
.fgallag( If51795ea140bec96fdefbc52291801b5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idc436d6b98d48c479d762c31bb55e071 = (I0cb5c7a759f4c75d4a675f9777f15c5f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If51795ea140bec96fdefbc52291801b5 ;

Ic9c2f173881d25f8976d723957809f51 Ieb6bb58bb679f765a9596c3b1c606590 (
.fgallag_sel( I0ca91c1426ba14a7b47a081cb3becd19[fgallag_SEL-1:0]),
.fgallag( Ib0a0f80cb818018b2fe0fd4597325bb4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I49300b5a8d4f2ce3ef7238f75a2800a9 = (I0ca91c1426ba14a7b47a081cb3becd19[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib0a0f80cb818018b2fe0fd4597325bb4 ;

Ic9c2f173881d25f8976d723957809f51 I03ef5580ac8c5f47afc1d4339bc154a4 (
.fgallag_sel( I0737e0cc7453e328efab2277bb712ea8[fgallag_SEL-1:0]),
.fgallag( If01a65e097f026a816133c34d73ccff1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4c1b051c518c4fa2e042e11cae60de02 = (I0737e0cc7453e328efab2277bb712ea8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If01a65e097f026a816133c34d73ccff1 ;

Ic9c2f173881d25f8976d723957809f51 I975a0d37c6e9ecbd273646b349aa3d10 (
.fgallag_sel( I456af863661122cc303fccb235f3c7a1[fgallag_SEL-1:0]),
.fgallag( Ida9ed61c543afde2257053443d133119 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3ccb0a4c235cd79c6c11271aa1aeb8af = (I456af863661122cc303fccb235f3c7a1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ida9ed61c543afde2257053443d133119 ;

Ic9c2f173881d25f8976d723957809f51 I6e8db33c89a9f7af7f5d336dfb2cfeae (
.fgallag_sel( Idc5916c4800e9f647d51c52444ab6fff[fgallag_SEL-1:0]),
.fgallag( I983a5656d68192a7a3d5a78f17f12ff0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8a2e9aba30b284e87bdbb6e91a30d9a6 = (Idc5916c4800e9f647d51c52444ab6fff[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I983a5656d68192a7a3d5a78f17f12ff0 ;

Ic9c2f173881d25f8976d723957809f51 Ib91d65750d256c04ff51fff7e3294dc6 (
.fgallag_sel( I57aca70e2b8d126c120736b2606ed333[fgallag_SEL-1:0]),
.fgallag( I315445ad2d762b66f94a75d76fbfb839 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I29d269323cfbc900f3868dde96e8da48 = (I57aca70e2b8d126c120736b2606ed333[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I315445ad2d762b66f94a75d76fbfb839 ;

Ic9c2f173881d25f8976d723957809f51 I20ef21b81718a1b8c5ee21ea8966eb90 (
.fgallag_sel( Ic6650a6d092b749b4498c08d69cf815e[fgallag_SEL-1:0]),
.fgallag( I7a97a8fe65e56b0a80c242e13e70db09 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I39a53ef95ccd9c8b1b85e3214af441f3 = (Ic6650a6d092b749b4498c08d69cf815e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7a97a8fe65e56b0a80c242e13e70db09 ;

Ic9c2f173881d25f8976d723957809f51 I0c454713281701cceab8e0d0c447aced (
.fgallag_sel( Ic2e3b8f91eb218650c7b9c515c7efe97[fgallag_SEL-1:0]),
.fgallag( I2243095f420e4d996f1c69c965932778 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id64ff7aeff6f73342f863be760a32a16 = (Ic2e3b8f91eb218650c7b9c515c7efe97[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2243095f420e4d996f1c69c965932778 ;

Ic9c2f173881d25f8976d723957809f51 I010b3a4893a69b888c132f486d05ffa2 (
.fgallag_sel( I93a084aa1e6881ab8dc905dcdcdfd7ee[fgallag_SEL-1:0]),
.fgallag( I0154a19f9adb43089080304978256c09 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I083900fbd062835b505165f1da19e228 = (I93a084aa1e6881ab8dc905dcdcdfd7ee[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0154a19f9adb43089080304978256c09 ;

Ic9c2f173881d25f8976d723957809f51 I589691139218824954a774b3ccec6ede (
.fgallag_sel( I8cba172573be52c5a90bd40e6f40a508[fgallag_SEL-1:0]),
.fgallag( Ib8bdc3b41b3cc7132c43833802115880 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7cf9dee91f849e28b2b2b38d2df00dfd = (I8cba172573be52c5a90bd40e6f40a508[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib8bdc3b41b3cc7132c43833802115880 ;

Ic9c2f173881d25f8976d723957809f51 Id1167d87a9926ce2ba4fb3c63a8574d7 (
.fgallag_sel( I1cccfd1516af59265731121dde878116[fgallag_SEL-1:0]),
.fgallag( I167586906b601ffc473a5b856b213f2b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If54b33370dcdf69c464c92dab1248828 = (I1cccfd1516af59265731121dde878116[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I167586906b601ffc473a5b856b213f2b ;

Ic9c2f173881d25f8976d723957809f51 I159ae5326f6e85c2cb000d19b9124483 (
.fgallag_sel( Ia171bbefe2d20b4c058126c33ef28eb8[fgallag_SEL-1:0]),
.fgallag( I094a6ac91aacfdd2f8de8a0d776f732b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I79c5230097571dcdf6ec2a15d633cdba = (Ia171bbefe2d20b4c058126c33ef28eb8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I094a6ac91aacfdd2f8de8a0d776f732b ;

Ic9c2f173881d25f8976d723957809f51 I46bc456dc38ad6c0b23ad70bd3994be9 (
.fgallag_sel( I84bc44a5d53a8f66b985b70c7ec1ae7c[fgallag_SEL-1:0]),
.fgallag( I9d4437c250c28653bbccdea6af8b6280 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I71efb4b4bb9b37a4e9b717282c5fbb03 = (I84bc44a5d53a8f66b985b70c7ec1ae7c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9d4437c250c28653bbccdea6af8b6280 ;

Ic9c2f173881d25f8976d723957809f51 If433b113c5e173e1dc0b5ea79c999e58 (
.fgallag_sel( I321b104ca3c818018d4b03adfe1110b9[fgallag_SEL-1:0]),
.fgallag( I4afab82ea1a6ad0a36fea0692de1d106 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0cc336baadd473b40a866cb2944eb719 = (I321b104ca3c818018d4b03adfe1110b9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4afab82ea1a6ad0a36fea0692de1d106 ;

Ic9c2f173881d25f8976d723957809f51 I5276b246863da0d3ae3c601016d0fb71 (
.fgallag_sel( Ia79b8994da536c86634bf6f54a21145d[fgallag_SEL-1:0]),
.fgallag( I864d41b77a51fda97ea7017ed18b5fea ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I42d8c11aefc92acf389d12e26217e867 = (Ia79b8994da536c86634bf6f54a21145d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I864d41b77a51fda97ea7017ed18b5fea ;

Ic9c2f173881d25f8976d723957809f51 I6fd8a3cd7231f43975c57b9e29a785ab (
.fgallag_sel( I4df55ce80eec5fee295b5a0ae92bd6c8[fgallag_SEL-1:0]),
.fgallag( I758ee12b430cda151b452699eb2039dc ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I40412ee4da7bae7c7745064488928be1 = (I4df55ce80eec5fee295b5a0ae92bd6c8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I758ee12b430cda151b452699eb2039dc ;

Ic9c2f173881d25f8976d723957809f51 If0c68128f1c6dc2a77eed22084ba5800 (
.fgallag_sel( I46593a7956590d870fe680228081a6d2[fgallag_SEL-1:0]),
.fgallag( I134cd61326b70030c027a3821d98a994 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7f6fc13ef5b20f9f1646a608b63f6f77 = (I46593a7956590d870fe680228081a6d2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I134cd61326b70030c027a3821d98a994 ;

Ic9c2f173881d25f8976d723957809f51 I2f982a5b45c20f43db618e3dee62f94a (
.fgallag_sel( I906e9da31de73ae45579607a014e8b54[fgallag_SEL-1:0]),
.fgallag( I99951d295b9065614c103b3e43fa255c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iddd6e6676bf1c96936bb1dbecf6fd805 = (I906e9da31de73ae45579607a014e8b54[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I99951d295b9065614c103b3e43fa255c ;

Ic9c2f173881d25f8976d723957809f51 Ie8053fbbcedbb617f26b6e37c2ba4559 (
.fgallag_sel( If5dd1a1b9e3fc0e67a85da3183480aed[fgallag_SEL-1:0]),
.fgallag( I31a4e4f3eac271c84b36c84d7de338fd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id0a701ba3adbf20de140020b675cc363 = (If5dd1a1b9e3fc0e67a85da3183480aed[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I31a4e4f3eac271c84b36c84d7de338fd ;

Ic9c2f173881d25f8976d723957809f51 If3148152dae0fa41bc06f0b9505f58ef (
.fgallag_sel( Iadfb1571c78c3f0c05e4ef498267df24[fgallag_SEL-1:0]),
.fgallag( Id36c36d2b2dd9a79f9887c9950b385c3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7e8db4d3310c345d7ada4c2fe05cf9b6 = (Iadfb1571c78c3f0c05e4ef498267df24[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id36c36d2b2dd9a79f9887c9950b385c3 ;

Ic9c2f173881d25f8976d723957809f51 I0bfa01a1f14953ae1eb71058f7320e35 (
.fgallag_sel( Icebb43b184c2745cc9da9d01b06bc62f[fgallag_SEL-1:0]),
.fgallag( I59455b0e53bac4fe6b1cbf609cb03da5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3fba42f5d091f0b7a5d8b4d099f72284 = (Icebb43b184c2745cc9da9d01b06bc62f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I59455b0e53bac4fe6b1cbf609cb03da5 ;

Ic9c2f173881d25f8976d723957809f51 Id6db3285ea0a8a85ea247bc993d4a525 (
.fgallag_sel( I6e4b0489ec7333abf2245a1b72a8923d[fgallag_SEL-1:0]),
.fgallag( Ifd633f2ea91cb88aaa2a0bf5579ed1e0 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia12c6ec292c6e9fdf58fe58a2af18a53 = (I6e4b0489ec7333abf2245a1b72a8923d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifd633f2ea91cb88aaa2a0bf5579ed1e0 ;

Ic9c2f173881d25f8976d723957809f51 I52518990a693861548758e440ad7a4bd (
.fgallag_sel( I24ac5dd30526c1d3bc7b941103a66804[fgallag_SEL-1:0]),
.fgallag( I87218b174c1db735ac153604b5ff3e15 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I37448ddc452e005ec974628ade793433 = (I24ac5dd30526c1d3bc7b941103a66804[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I87218b174c1db735ac153604b5ff3e15 ;

Ic9c2f173881d25f8976d723957809f51 If44ee0e04b5c92d80f41c75e8eb9dd35 (
.fgallag_sel( I33681b2292c086fe536dae2aec70903a[fgallag_SEL-1:0]),
.fgallag( I4608c92d52306432c114f31b9ba6dd69 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4dee5017c9b71edda82d50b867879afd = (I33681b2292c086fe536dae2aec70903a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4608c92d52306432c114f31b9ba6dd69 ;

Ic9c2f173881d25f8976d723957809f51 I5ab5070def1078571d6c4438c2a764a6 (
.fgallag_sel( Ia373ca76c3b15a4148532b3822f82ba5[fgallag_SEL-1:0]),
.fgallag( Iba3f6cde40827d82bc32078344b9bd81 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2115d9af1cbecde8b5e89c70e582de00 = (Ia373ca76c3b15a4148532b3822f82ba5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iba3f6cde40827d82bc32078344b9bd81 ;

Ic9c2f173881d25f8976d723957809f51 I7f4228ac2fd344a5e1be2fc8c91fa44e (
.fgallag_sel( I7d08adbaf66cea04be4891db610bca3f[fgallag_SEL-1:0]),
.fgallag( Ib987bde3ee5a0256d0b8b3aa7357cdb2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0e2c6c08e1bcd629678ff57f6bf23be5 = (I7d08adbaf66cea04be4891db610bca3f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib987bde3ee5a0256d0b8b3aa7357cdb2 ;

Ic9c2f173881d25f8976d723957809f51 I67298566fd91c0dec771f226471a7464 (
.fgallag_sel( Ic09ed51b20f411683a801eaad61657a3[fgallag_SEL-1:0]),
.fgallag( I3c33a2bfaa82172457b15f4f621eefee ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I00a3c15421af76c65865ff21d2598055 = (Ic09ed51b20f411683a801eaad61657a3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3c33a2bfaa82172457b15f4f621eefee ;

Ic9c2f173881d25f8976d723957809f51 I6df6597f22915996d5a9507aa66210a1 (
.fgallag_sel( I6a9af8c9009b5de47ebe9ee8b79d3831[fgallag_SEL-1:0]),
.fgallag( I7ce33eb337b6cacaea13f748061e338a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I9fa21fd04ffc0a7dc281717e599fd443 = (I6a9af8c9009b5de47ebe9ee8b79d3831[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7ce33eb337b6cacaea13f748061e338a ;

Ic9c2f173881d25f8976d723957809f51 Ifdbb60bb17060ff7394f0578884c4701 (
.fgallag_sel( Ife18e8a16d4437161b75a93e3dff1b5b[fgallag_SEL-1:0]),
.fgallag( I7a8c5be75d87552ca717a87d1a832d21 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I66231fd914db4a60705f1d6de751077d = (Ife18e8a16d4437161b75a93e3dff1b5b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7a8c5be75d87552ca717a87d1a832d21 ;

Ic9c2f173881d25f8976d723957809f51 I869a679dd2b6e83b5dc89daab8944600 (
.fgallag_sel( I0cde86532c8db1a32d9fbe38a40b91b8[fgallag_SEL-1:0]),
.fgallag( Id9c9cebf44647040da33567d815c261f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1142cf230d2632a5972a95316f2fa15f = (I0cde86532c8db1a32d9fbe38a40b91b8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id9c9cebf44647040da33567d815c261f ;

Ic9c2f173881d25f8976d723957809f51 I6110ea6b5b20ab24f4d4ab29ada8c4d6 (
.fgallag_sel( I49c8ec4cd33e6caed8ed7dab779e7ebb[fgallag_SEL-1:0]),
.fgallag( I6c522c28a0dc265facb1f21ebe51c564 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibe1b4cc79b063aafddadcfdb5bc4a694 = (I49c8ec4cd33e6caed8ed7dab779e7ebb[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6c522c28a0dc265facb1f21ebe51c564 ;

Ic9c2f173881d25f8976d723957809f51 Id09365d68f7ee2f0a3f5d15b1194aee7 (
.fgallag_sel( Idb86f95570587a0711d796aac7004c25[fgallag_SEL-1:0]),
.fgallag( I86c367b0fd4548d5edfb8863f454653e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5371e6575d8bdc6f72cb08beca627fec = (Idb86f95570587a0711d796aac7004c25[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I86c367b0fd4548d5edfb8863f454653e ;

Ic9c2f173881d25f8976d723957809f51 I9590c0120faaa50974110a72630aaf74 (
.fgallag_sel( I2d1373d0b18992fa46a9607a86d21520[fgallag_SEL-1:0]),
.fgallag( I800271efe85fcbaee8fe733190e90f6d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5e78e43fbf13f79a885bb3cee615d926 = (I2d1373d0b18992fa46a9607a86d21520[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I800271efe85fcbaee8fe733190e90f6d ;

Ic9c2f173881d25f8976d723957809f51 I68839d3864f567fdea045324b6782f8e (
.fgallag_sel( I30f26e090ab14551cbac41883ad8a152[fgallag_SEL-1:0]),
.fgallag( Ia5172996abb4a6bc50046d36ec033c7f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I735298e3ea4442615df21b3699c94a7d = (I30f26e090ab14551cbac41883ad8a152[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia5172996abb4a6bc50046d36ec033c7f ;

Ic9c2f173881d25f8976d723957809f51 If5221554fef224a107bd55fdeb5e3fd4 (
.fgallag_sel( Ib1b4e41ab25733d1d6dd54e1fe81a419[fgallag_SEL-1:0]),
.fgallag( Ibe20363746d437eef2c85360425739d1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1f2f072bb15b57b5437572b156499e12 = (Ib1b4e41ab25733d1d6dd54e1fe81a419[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibe20363746d437eef2c85360425739d1 ;

Ic9c2f173881d25f8976d723957809f51 Iaf2cd419671cb542c16743a2d2c7b921 (
.fgallag_sel( I146c0d5154a6de44c0536de873904ccf[fgallag_SEL-1:0]),
.fgallag( Iee695b22e8a55479dfcbaa68f5c8b6c9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0344e18f3a5fe97467ba8e6641562f92 = (I146c0d5154a6de44c0536de873904ccf[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iee695b22e8a55479dfcbaa68f5c8b6c9 ;

Ic9c2f173881d25f8976d723957809f51 I24b77aaf5f9d7b4bcae5cd804cf5e45b (
.fgallag_sel( I8eb9d4839a478a4e28b45a549b5682a4[fgallag_SEL-1:0]),
.fgallag( I7cdb0bf6c7195df38d701768e655af70 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8aedaf42a56212b44d820d704945cb99 = (I8eb9d4839a478a4e28b45a549b5682a4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7cdb0bf6c7195df38d701768e655af70 ;

Ic9c2f173881d25f8976d723957809f51 I6555238dc6b5abb09d90cc9a157a33c8 (
.fgallag_sel( I2501ef991a59512c43693ba9d7db8571[fgallag_SEL-1:0]),
.fgallag( I1057373671fd4cfba6696f8e88a2d740 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If267b8451ce8bfd1c33273a9c5d08233 = (I2501ef991a59512c43693ba9d7db8571[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1057373671fd4cfba6696f8e88a2d740 ;

Ic9c2f173881d25f8976d723957809f51 Iba5d5e99f6ada37414e148588aed5c65 (
.fgallag_sel( I38213f78fd4dc52f9d2c9b7b22136c1c[fgallag_SEL-1:0]),
.fgallag( I7dd9da64c1516e6ae1b703defc4cdc55 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie90356409910181f0ffbfdbfea6a47b2 = (I38213f78fd4dc52f9d2c9b7b22136c1c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7dd9da64c1516e6ae1b703defc4cdc55 ;

Ic9c2f173881d25f8976d723957809f51 Ie8eeefbd835bd32725592c37eac588ac (
.fgallag_sel( I49ce91ac152279af421bbc6c4d9b8087[fgallag_SEL-1:0]),
.fgallag( I58bf5f51208a98b2448e2b4fad3f63ac ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I43a2d55679515c4766a6e7c19c3ba1e0 = (I49ce91ac152279af421bbc6c4d9b8087[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I58bf5f51208a98b2448e2b4fad3f63ac ;

Ic9c2f173881d25f8976d723957809f51 Ie551a2d96d31e139ccf96150bf80395c (
.fgallag_sel( I6a2b7bb2cb3ca2ab932c211a68dded55[fgallag_SEL-1:0]),
.fgallag( Icb8281c05ea7168d39d6012a1d622e15 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2b1e17eeb208749a9c320187e98f3c50 = (I6a2b7bb2cb3ca2ab932c211a68dded55[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Icb8281c05ea7168d39d6012a1d622e15 ;

Ic9c2f173881d25f8976d723957809f51 Ib441a835fe7d91e57ec34a8de3089e09 (
.fgallag_sel( Idaae6ba9da8754615a2c34ef859492db[fgallag_SEL-1:0]),
.fgallag( I5b16ad2952938bc64f6c9f5ff1ab5a0b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib9c8fc92cd361858e4fb1ddc6dcab191 = (Idaae6ba9da8754615a2c34ef859492db[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5b16ad2952938bc64f6c9f5ff1ab5a0b ;

Ic9c2f173881d25f8976d723957809f51 I435d71506982ba90da657ea137e2d63d (
.fgallag_sel( Icaca9fc70a3ec6c48c0e41f8168e2bb9[fgallag_SEL-1:0]),
.fgallag( I5d5790b480d08bf6c957f26e24467b9a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7ef5a40bcc9976da690ae85ee866b2d0 = (Icaca9fc70a3ec6c48c0e41f8168e2bb9[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5d5790b480d08bf6c957f26e24467b9a ;

Ic9c2f173881d25f8976d723957809f51 I213684e46324a3ff95a4ee51ba067fbe (
.fgallag_sel( I4f69b8ff834c7ab3194bc9390ce0f5f6[fgallag_SEL-1:0]),
.fgallag( Ieb32ca618265eed3419f01907f48527d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia52b8e11416781165d713f38018047d6 = (I4f69b8ff834c7ab3194bc9390ce0f5f6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ieb32ca618265eed3419f01907f48527d ;

Ic9c2f173881d25f8976d723957809f51 Iebc9408ba0214534b1a6d33f560628ba (
.fgallag_sel( I037cb596cd48c5533ed22bc32518d992[fgallag_SEL-1:0]),
.fgallag( Ief90415b272ce5707ba28a8470132f5e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ibb05d1616c4b57cdf6a268fe16bb9ef9 = (I037cb596cd48c5533ed22bc32518d992[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ief90415b272ce5707ba28a8470132f5e ;

Ic9c2f173881d25f8976d723957809f51 I22e82d556852a28ef200935edf5193fe (
.fgallag_sel( I94a89577951de90edc4f73b281ad7364[fgallag_SEL-1:0]),
.fgallag( I386c79f4301dea9a37c9ce283e8050e4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3be04ed5b262f461ad65b860adc6c601 = (I94a89577951de90edc4f73b281ad7364[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I386c79f4301dea9a37c9ce283e8050e4 ;

Ic9c2f173881d25f8976d723957809f51 I5b41d68c073243e5ae729ef9d4cf97ae (
.fgallag_sel( Ib7493a1a384aebaa7999ff1fb867fc6b[fgallag_SEL-1:0]),
.fgallag( I0d113fab9d7095f8d1693fec58b7c5a6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0bcc8dd8d2adfb33dace6c005377ef97 = (Ib7493a1a384aebaa7999ff1fb867fc6b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0d113fab9d7095f8d1693fec58b7c5a6 ;

Ic9c2f173881d25f8976d723957809f51 I88219dfbe8661aaa58d2198fbf8ba1e6 (
.fgallag_sel( I2ceb9e423696539135c5bae5cc2d8d98[fgallag_SEL-1:0]),
.fgallag( I2bbbe9e5d322d9cee76903fa813765ae ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iad8fd338d5a105b6fe3a3a021f96f317 = (I2ceb9e423696539135c5bae5cc2d8d98[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2bbbe9e5d322d9cee76903fa813765ae ;

Ic9c2f173881d25f8976d723957809f51 Ic7dfdaf75266325d4e76042ac6c06b6c (
.fgallag_sel( Ia6bbf236436b2ed22bbaae3b8849de6d[fgallag_SEL-1:0]),
.fgallag( If5317506b6ab92c946af745a65b9e86a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I46f7c02eeea9f5a0058da869a84e57d4 = (Ia6bbf236436b2ed22bbaae3b8849de6d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If5317506b6ab92c946af745a65b9e86a ;

Ic9c2f173881d25f8976d723957809f51 I19a8c895bfa5733d8850f95258a5640c (
.fgallag_sel( I33cdaee4676d546dd5507df4704ea1f8[fgallag_SEL-1:0]),
.fgallag( Ib61ddb3ef6c7239bfc720b1761cc0221 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie8e3dd32f3ccf581400d8dd0fd5daea7 = (I33cdaee4676d546dd5507df4704ea1f8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib61ddb3ef6c7239bfc720b1761cc0221 ;

Ic9c2f173881d25f8976d723957809f51 I9890884d78850f0d13ecba0d2f56b907 (
.fgallag_sel( Ia44daa9ddc3e4d377267333813d4675f[fgallag_SEL-1:0]),
.fgallag( I70d669976b271b2319d60114c468cae5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic23bbefb8e8e80ac5df4ef8a50aa5c83 = (Ia44daa9ddc3e4d377267333813d4675f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I70d669976b271b2319d60114c468cae5 ;

Ic9c2f173881d25f8976d723957809f51 I015a4348e263d8baa48dec35756820ab (
.fgallag_sel( Ie1f8fff3f43426d6bc39e45322a532ca[fgallag_SEL-1:0]),
.fgallag( I96cb81892e2d1737d6cb25522ea2d9e4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7c56e54d472bc2301521ecb93aed0ea2 = (Ie1f8fff3f43426d6bc39e45322a532ca[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I96cb81892e2d1737d6cb25522ea2d9e4 ;

Ic9c2f173881d25f8976d723957809f51 Id3d58bc2ba46c1a500292b1051be6789 (
.fgallag_sel( I4ee181895efc22862b6e85802a944095[fgallag_SEL-1:0]),
.fgallag( I6c87926b040d4006c2294c516a3c46fd ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4979d09a4bf88992a280e598841f5e50 = (I4ee181895efc22862b6e85802a944095[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6c87926b040d4006c2294c516a3c46fd ;

Ic9c2f173881d25f8976d723957809f51 I4ecd0d1de0e5723dff1b42a974feb232 (
.fgallag_sel( I5c24ea83cabbb6be089ac084732cb9d6[fgallag_SEL-1:0]),
.fgallag( I549670efc854cdc29bad1d9bc03e9f5e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I15264bbbe49fff9c53b8066414264010 = (I5c24ea83cabbb6be089ac084732cb9d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I549670efc854cdc29bad1d9bc03e9f5e ;

Ic9c2f173881d25f8976d723957809f51 Ia5eb6ebf84dbd8a9e4191edab70e98d0 (
.fgallag_sel( Ifee2342449a3b3d0036ce2ecbc9ae189[fgallag_SEL-1:0]),
.fgallag( If54c0c169048bb3e8a1423a58aed0e70 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I32293d41086053c7055fa40ce224631e = (Ifee2342449a3b3d0036ce2ecbc9ae189[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If54c0c169048bb3e8a1423a58aed0e70 ;

Ic9c2f173881d25f8976d723957809f51 I1462d1260cf75ce4e7760a38bd918441 (
.fgallag_sel( I70a9a9b8f25066612a50e411ad68e6c4[fgallag_SEL-1:0]),
.fgallag( I5c956f39031611db595fbc34e6edad65 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4bd0008f9e9598e9f60a0aa8c2aa2da5 = (I70a9a9b8f25066612a50e411ad68e6c4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5c956f39031611db595fbc34e6edad65 ;

Ic9c2f173881d25f8976d723957809f51 I1d12b2cb36a10b9475f6d36ac19efd6f (
.fgallag_sel( I1870059af857c79d444bef948bb536ef[fgallag_SEL-1:0]),
.fgallag( I86851725f5d424c4636f9f41e5a7c7e9 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I584861d31ee7ff0efc61b192c64bca32 = (I1870059af857c79d444bef948bb536ef[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I86851725f5d424c4636f9f41e5a7c7e9 ;

Ic9c2f173881d25f8976d723957809f51 Ie3ac3567e9a6289fbe772e115fb3cb79 (
.fgallag_sel( Iafe61ab12e232a1090123a0f16eefaca[fgallag_SEL-1:0]),
.fgallag( Ibec300322cef05615c818b163f8a1fef ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I64f092a873fee78a333072d8c5bbddf8 = (Iafe61ab12e232a1090123a0f16eefaca[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibec300322cef05615c818b163f8a1fef ;

Ic9c2f173881d25f8976d723957809f51 Id2b71fd2e51212154de024a9836061d1 (
.fgallag_sel( I10ca809fe9a04eaf5d7784ba69314178[fgallag_SEL-1:0]),
.fgallag( I09cc443ecf3811a8a672c4aec1f7d6d4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idd6f95a4386cbea3c1533683854a4c75 = (I10ca809fe9a04eaf5d7784ba69314178[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I09cc443ecf3811a8a672c4aec1f7d6d4 ;

Ic9c2f173881d25f8976d723957809f51 I17fd994c1119f7c9ddc3be4595e3bab5 (
.fgallag_sel( I7a1bd0a115b3a1f85cb9c54840f5bf9b[fgallag_SEL-1:0]),
.fgallag( Iaaf5b9288b4eb557d56908bf072cc642 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I32710d1855b18d6c70f6e23a0a440a69 = (I7a1bd0a115b3a1f85cb9c54840f5bf9b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iaaf5b9288b4eb557d56908bf072cc642 ;

Ic9c2f173881d25f8976d723957809f51 I13260b5b97c2a18aef5893601275c0e9 (
.fgallag_sel( I986a564393d944d7d202414431c6d165[fgallag_SEL-1:0]),
.fgallag( Ib224ff2bea17f6e694b10bc7cfdb898d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I32cc6023f28c6dee2b4b097f1fe890d6 = (I986a564393d944d7d202414431c6d165[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib224ff2bea17f6e694b10bc7cfdb898d ;

Ic9c2f173881d25f8976d723957809f51 I4dabb2412daef4712958ca6250645619 (
.fgallag_sel( I464042aaa60a41c7e1faf3d16eeb121d[fgallag_SEL-1:0]),
.fgallag( Ide7d6472bf33f8dcf5c6397c7d7fb733 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Id91b5daa1685f0e3d492f0c3c8306f8e = (I464042aaa60a41c7e1faf3d16eeb121d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ide7d6472bf33f8dcf5c6397c7d7fb733 ;

Ic9c2f173881d25f8976d723957809f51 Id028fce86a2691dab71412b8b4ad7bd8 (
.fgallag_sel( I34b9a0bf2b6b562fb36291022ddf5179[fgallag_SEL-1:0]),
.fgallag( Ie6193636ea1cba8b71e1d0d5f2e3c1b2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icfdd224aa430648d4afe7b224340b91d = (I34b9a0bf2b6b562fb36291022ddf5179[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie6193636ea1cba8b71e1d0d5f2e3c1b2 ;

Ic9c2f173881d25f8976d723957809f51 I9f02d3be67cbe16c9123384cbd4c102c (
.fgallag_sel( I17dd8612b5c7f9dcc90f17e584aab2d3[fgallag_SEL-1:0]),
.fgallag( Id631b0a4de889a3c3eff4df79367d3d4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icbcaa7780b1ad02e07cbbc871b0c2729 = (I17dd8612b5c7f9dcc90f17e584aab2d3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id631b0a4de889a3c3eff4df79367d3d4 ;

Ic9c2f173881d25f8976d723957809f51 I9b4df2dbbc89b68f1b735a4bca80ea16 (
.fgallag_sel( Id77cf7c05844d83e808a694971145261[fgallag_SEL-1:0]),
.fgallag( I93d80b8bfb77e7af4d9ac734f26c4e62 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I587b0b57b4f95e8533842965674d1416 = (Id77cf7c05844d83e808a694971145261[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I93d80b8bfb77e7af4d9ac734f26c4e62 ;

Ic9c2f173881d25f8976d723957809f51 I230f298160d73fb907087a727b8fae7e (
.fgallag_sel( I276c1155d766437253f12b25066b84e4[fgallag_SEL-1:0]),
.fgallag( I7fba5fee37c5912e7f635feb8c111b3a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1188961bb659f61f0749a27f4ee5c62d = (I276c1155d766437253f12b25066b84e4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7fba5fee37c5912e7f635feb8c111b3a ;

Ic9c2f173881d25f8976d723957809f51 I5380abd15601365f1b6c392348ce409b (
.fgallag_sel( Id75b386d8076893cb73baca69c3eff59[fgallag_SEL-1:0]),
.fgallag( I22c14ad43399d8a1aee258826a71f50e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4ed124c919ba9e29d61a5f771b554ead = (Id75b386d8076893cb73baca69c3eff59[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I22c14ad43399d8a1aee258826a71f50e ;

Ic9c2f173881d25f8976d723957809f51 I618657ae53efd25255efe715e3596a8c (
.fgallag_sel( If62ddbe87274965cfd83189c6666401e[fgallag_SEL-1:0]),
.fgallag( I3bdc4806c5c09de9a7de8d3601c57bfe ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I735b52f16a8beb195d3e7332f39a1c86 = (If62ddbe87274965cfd83189c6666401e[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3bdc4806c5c09de9a7de8d3601c57bfe ;

Ic9c2f173881d25f8976d723957809f51 I50943a2e35d7f91e5e297acb5b48ccce (
.fgallag_sel( I4f73a07452638a610b31e3ee52cb5639[fgallag_SEL-1:0]),
.fgallag( Id451569510e0d1bbba9002c2b27bb3d4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I626977a5bbbdb2da503472e8fe6c9569 = (I4f73a07452638a610b31e3ee52cb5639[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Id451569510e0d1bbba9002c2b27bb3d4 ;

Ic9c2f173881d25f8976d723957809f51 Ibf7f0e15ce49042f297d3039f3a4afd9 (
.fgallag_sel( I2a4faf3344d9bf4ee71da0be8994788a[fgallag_SEL-1:0]),
.fgallag( I16753a377bced0688797a464157d847b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8f2450ac5c97afe557d068ee5760b527 = (I2a4faf3344d9bf4ee71da0be8994788a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I16753a377bced0688797a464157d847b ;

Ic9c2f173881d25f8976d723957809f51 I29f9d5575c7a1f4ac9e0ff546a9923e1 (
.fgallag_sel( I7d7ad0cbb962a47e229fe9d8406e6fe1[fgallag_SEL-1:0]),
.fgallag( I76fd17f22401b66bfc0a6239a0518157 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I13834193a9eb2706cdc680b303efbcf4 = (I7d7ad0cbb962a47e229fe9d8406e6fe1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I76fd17f22401b66bfc0a6239a0518157 ;

Ic9c2f173881d25f8976d723957809f51 Iecd52fca7eeea3bd155a25098ee8baaf (
.fgallag_sel( I82988dc2dc83ac61380d2a5cb6551768[fgallag_SEL-1:0]),
.fgallag( Ie56f8b245ab7833b6939cfea43a99874 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I798a185688b52e59c92b42161b3da7e7 = (I82988dc2dc83ac61380d2a5cb6551768[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie56f8b245ab7833b6939cfea43a99874 ;

Ic9c2f173881d25f8976d723957809f51 I0066620f14ea9cec68706bf1c59bfb04 (
.fgallag_sel( I058c3a9848fd30010e4742d8682081ac[fgallag_SEL-1:0]),
.fgallag( I668f8103700f044c7764f2281a5b457e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib695cf55b921ed43db22362a28761714 = (I058c3a9848fd30010e4742d8682081ac[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I668f8103700f044c7764f2281a5b457e ;

Ic9c2f173881d25f8976d723957809f51 I0391d29c781ac99c264636c4ddcb6757 (
.fgallag_sel( I368121c2534820a7147858c06e58b3fc[fgallag_SEL-1:0]),
.fgallag( Ib75c0ca4f8b59afc2fdd7793bff7ad16 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1dd0afb6f1a979176d01ab7d37f39bed = (I368121c2534820a7147858c06e58b3fc[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib75c0ca4f8b59afc2fdd7793bff7ad16 ;

Ic9c2f173881d25f8976d723957809f51 Id2ba0e2207bb2242027b02463f8bb759 (
.fgallag_sel( I03d4541eeb1440aa72ee490c49977e32[fgallag_SEL-1:0]),
.fgallag( I3d39fa04d24aa69d19a2db8da00eb0d3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I559878eee7f3bee345a0f0e891dd2c05 = (I03d4541eeb1440aa72ee490c49977e32[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I3d39fa04d24aa69d19a2db8da00eb0d3 ;

Ic9c2f173881d25f8976d723957809f51 I676651d40efa36606ddd64f3490d1e9e (
.fgallag_sel( I75fdf5a355949a87b768b1e67db674e4[fgallag_SEL-1:0]),
.fgallag( I284b4ccbcb23293efe64fa45b2e0ad98 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6c688b7c6f01ae353117029f80487ec4 = (I75fdf5a355949a87b768b1e67db674e4[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I284b4ccbcb23293efe64fa45b2e0ad98 ;

Ic9c2f173881d25f8976d723957809f51 I8fd3ef8ffc5ab44d7c28c2a1aa635388 (
.fgallag_sel( I088f4a0af0239602d422324549cb9799[fgallag_SEL-1:0]),
.fgallag( I689ac029a268fe244a8793367c900602 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I62ad8f36d1e0b80d0d04a326d80e1729 = (I088f4a0af0239602d422324549cb9799[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I689ac029a268fe244a8793367c900602 ;

Ic9c2f173881d25f8976d723957809f51 Ic5c5d93d488f1c29e28b1496d31561a4 (
.fgallag_sel( I787fe66b38237caf805ec14970d154c7[fgallag_SEL-1:0]),
.fgallag( If53dace3e8a7be2524d711de84855015 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icf1eb32cfc4a48f7e53c180aa94f5833 = (I787fe66b38237caf805ec14970d154c7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If53dace3e8a7be2524d711de84855015 ;

Ic9c2f173881d25f8976d723957809f51 Ie115e9e1e43ecc22abc68d9d823c8443 (
.fgallag_sel( Icef176cff3ae503dbbe2af9ecfc4c859[fgallag_SEL-1:0]),
.fgallag( Ie3fe635b63e13732c17ae2076b807b4d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I8bdfadcfa5cb308e6e254d42997340fd = (Icef176cff3ae503dbbe2af9ecfc4c859[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie3fe635b63e13732c17ae2076b807b4d ;

Ic9c2f173881d25f8976d723957809f51 Id6b1d065dab621ac94eb885f1645587d (
.fgallag_sel( Ie0a66e4871bfe94f6716279ecc9ef21c[fgallag_SEL-1:0]),
.fgallag( I1e196a61113d4db7b51f3d6b18c33da3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I6ceae370fa59e601566286b127dec684 = (Ie0a66e4871bfe94f6716279ecc9ef21c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I1e196a61113d4db7b51f3d6b18c33da3 ;

Ic9c2f173881d25f8976d723957809f51 Ie8ce0795f61db0b467a4bfbfc6784f9e (
.fgallag_sel( I474adf7a975b405c288058139a08be38[fgallag_SEL-1:0]),
.fgallag( Ic80e494400a5d7dcfdbf96424391e596 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifcf5bef8ae2998f0bd3d270e98acc1c5 = (I474adf7a975b405c288058139a08be38[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic80e494400a5d7dcfdbf96424391e596 ;

Ic9c2f173881d25f8976d723957809f51 I4831974ec4260337376913a53b391a6b (
.fgallag_sel( Iebeadb39658f41dcf8719ed413e46144[fgallag_SEL-1:0]),
.fgallag( I69d20a7aaf2c66ed9b41fdeff0d5c6ec ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic1c8e5992501f0e04191fe6dadd2d56c = (Iebeadb39658f41dcf8719ed413e46144[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I69d20a7aaf2c66ed9b41fdeff0d5c6ec ;

Ic9c2f173881d25f8976d723957809f51 I87fec69bdb0bd3eb8587f427c27baf20 (
.fgallag_sel( Ie018b0d9f05a86207ae09ca2efac54e2[fgallag_SEL-1:0]),
.fgallag( I19b667bdb053ebd555aaa540d3a76f95 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I3f88a35a94c77ca32f3b58c4b509b21c = (Ie018b0d9f05a86207ae09ca2efac54e2[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I19b667bdb053ebd555aaa540d3a76f95 ;

Ic9c2f173881d25f8976d723957809f51 I63933085bfd52b8589c425e4d1880505 (
.fgallag_sel( I51ee69807609fca0f332c8bc31afd632[fgallag_SEL-1:0]),
.fgallag( Ifc3d9cc420aa1274fed24b38c4d9fd8a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib875be40a1b73b1583cfc9cfec760e31 = (I51ee69807609fca0f332c8bc31afd632[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifc3d9cc420aa1274fed24b38c4d9fd8a ;

Ic9c2f173881d25f8976d723957809f51 I427eb756e21fbc83d63602102f423723 (
.fgallag_sel( Iee1cb471704b2a8718a68ef93fd2e356[fgallag_SEL-1:0]),
.fgallag( Ie8a6ed15370edd38bfc92290bf7bb55a ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I15eae5f35300569305dc03e24d1cdd7f = (Iee1cb471704b2a8718a68ef93fd2e356[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie8a6ed15370edd38bfc92290bf7bb55a ;

Ic9c2f173881d25f8976d723957809f51 I2001703c2fc4e81de149127b3811614b (
.fgallag_sel( I1731c0e3be86eec142c3732ee836e4d5[fgallag_SEL-1:0]),
.fgallag( Ife5a1b49d4b0342f06ef83750ab914d4 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Idffbcb47f4a04fc71d1406e46f4ab6c4 = (I1731c0e3be86eec142c3732ee836e4d5[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ife5a1b49d4b0342f06ef83750ab914d4 ;

Ic9c2f173881d25f8976d723957809f51 I141fe3b3fc14f9f4a3710ba55df6fa72 (
.fgallag_sel( Id3b8c0ca32331f94fd98c8dae72bb15d[fgallag_SEL-1:0]),
.fgallag( I9906c49536062867b98ed290e49bbe50 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ifaf09d72a75fd4f9948e997b8a8388f4 = (Id3b8c0ca32331f94fd98c8dae72bb15d[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9906c49536062867b98ed290e49bbe50 ;

Ic9c2f173881d25f8976d723957809f51 I0e2ba3cfb7dabc7ad578ff3a0f1a7152 (
.fgallag_sel( I6a86b0a82441c6c14436a3e0af6b0fb7[fgallag_SEL-1:0]),
.fgallag( I41be66295070bec696e91d0f9efdc233 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I661c1624e4d13ba49efc3fb608ba84ed = (I6a86b0a82441c6c14436a3e0af6b0fb7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I41be66295070bec696e91d0f9efdc233 ;

Ic9c2f173881d25f8976d723957809f51 Ic49593b29bb52ef4ccd4fa76fa0b8dd0 (
.fgallag_sel( I8c92ff598084da7a50f7c68da96620b3[fgallag_SEL-1:0]),
.fgallag( I4838b956d8a597e78bef9a0fce82542e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iaa8bf572a01757f5e9321e6ff7364d7e = (I8c92ff598084da7a50f7c68da96620b3[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4838b956d8a597e78bef9a0fce82542e ;

Ic9c2f173881d25f8976d723957809f51 Ibd04af4e95d6959272321b69d0e8b063 (
.fgallag_sel( I8bd1862e7bc2e83e9863389d532e6623[fgallag_SEL-1:0]),
.fgallag( Ia06cb40e9a3341f34625c5804e02c07f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I7ef389b5ce4bdcca7fab9e9ec2bfa3a9 = (I8bd1862e7bc2e83e9863389d532e6623[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ia06cb40e9a3341f34625c5804e02c07f ;

Ic9c2f173881d25f8976d723957809f51 Ie4af77771bdc7fe3b128bbfe73b03891 (
.fgallag_sel( I8053269f8bd78a931878c8350693e1d6[fgallag_SEL-1:0]),
.fgallag( I4eaad70758412eab097822b2feda7a57 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4e7823ff42f8f44a21778dc4b3633a67 = (I8053269f8bd78a931878c8350693e1d6[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I4eaad70758412eab097822b2feda7a57 ;

Ic9c2f173881d25f8976d723957809f51 I6cafdc41428d4ef02166506e9f177213 (
.fgallag_sel( I2ff66cdd7314276232715ef2361ad184[fgallag_SEL-1:0]),
.fgallag( If89e1da3daa6fd3090781723173b140b ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icf5823b64f3a9b7d2656656b61724bcd = (I2ff66cdd7314276232715ef2361ad184[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If89e1da3daa6fd3090781723173b140b ;

Ic9c2f173881d25f8976d723957809f51 I21d7c3c44854d7cd2e9fcdd1a05195c7 (
.fgallag_sel( Icf541c76bfaf37fe6111de037d205f15[fgallag_SEL-1:0]),
.fgallag( I9ac67c519fd5a55d0ffb727389781492 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If77f93c61b38d10360f7dd382686d91c = (Icf541c76bfaf37fe6111de037d205f15[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9ac67c519fd5a55d0ffb727389781492 ;

Ic9c2f173881d25f8976d723957809f51 I7c54785ad1983edede61607f2eaabe02 (
.fgallag_sel( I68319c8b9febef9f564832429c91b85a[fgallag_SEL-1:0]),
.fgallag( I73799799e5469ae887dec9b46c9c965d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iede699ff40abf5838b54678df24ff29d = (I68319c8b9febef9f564832429c91b85a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I73799799e5469ae887dec9b46c9c965d ;

Ic9c2f173881d25f8976d723957809f51 I062cc69bd2d35df46712ae449cdf6fc4 (
.fgallag_sel( I127772614218dd7c50d3136b4f174d7a[fgallag_SEL-1:0]),
.fgallag( I7ebd7c3f0617cf500deeb8c152c09af2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia1c9e86b6112a18e7aa613315343e696 = (I127772614218dd7c50d3136b4f174d7a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7ebd7c3f0617cf500deeb8c152c09af2 ;

Ic9c2f173881d25f8976d723957809f51 I0edf3f4b59b3a14b3f2b6ca4623a9eb8 (
.fgallag_sel( Ib8d1aea4ad24c6ceb44f2cc672e1ff90[fgallag_SEL-1:0]),
.fgallag( I2ee7d4f522ba17ca941c67079309c398 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iad94272a2a302f4b6b963e71ccd64ccb = (Ib8d1aea4ad24c6ceb44f2cc672e1ff90[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I2ee7d4f522ba17ca941c67079309c398 ;

Ic9c2f173881d25f8976d723957809f51 Ib31105edeec2e178ca9e1f11bef1ed65 (
.fgallag_sel( I9ca26c8104bf15f48b19dc3256914544[fgallag_SEL-1:0]),
.fgallag( I62d13683ba05cfc27d9ae9a82fb04689 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If4d54d2b483d85b0c4f31db721b14323 = (I9ca26c8104bf15f48b19dc3256914544[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I62d13683ba05cfc27d9ae9a82fb04689 ;

Ic9c2f173881d25f8976d723957809f51 I0577d005af2354173029c2b12b454900 (
.fgallag_sel( Icc76d9ffc3f3d7b410205eeb8232a33b[fgallag_SEL-1:0]),
.fgallag( Ic06032eaed49f01d3d5513b2d145eaaf ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ia3b12887d984da936d88d657090f8972 = (Icc76d9ffc3f3d7b410205eeb8232a33b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ic06032eaed49f01d3d5513b2d145eaaf ;

Ic9c2f173881d25f8976d723957809f51 Ic42dac21bec10ba6d167380493515694 (
.fgallag_sel( I7fc4551d8a0445f79b87b4ba5f2ffeaa[fgallag_SEL-1:0]),
.fgallag( Idba6350812d3c90bee79636db48257e2 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib23dbfa64e4a9364e0c1dbbc6b2ff001 = (I7fc4551d8a0445f79b87b4ba5f2ffeaa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Idba6350812d3c90bee79636db48257e2 ;

Ic9c2f173881d25f8976d723957809f51 I3f6c1df4c11a063825289c5a4b20bc65 (
.fgallag_sel( I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8[fgallag_SEL-1:0]),
.fgallag( I6e7ed391604c7e0ff7cca99d5aeddc9f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ic8d47dcabda3b23d4451e609395c4698 = (I6b3c66c4e3fa0ef0cf0b52eaa4dac7a8[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6e7ed391604c7e0ff7cca99d5aeddc9f ;

Ic9c2f173881d25f8976d723957809f51 I956083b6b145aa35a105fa009b67c625 (
.fgallag_sel( Ie34c07af9f6adb9e4b636dce3d0682c0[fgallag_SEL-1:0]),
.fgallag( Ib78d45cc282f110ed3ddaeb706a0fc12 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5d4903ecdf83967c7f60d876bcd0b215 = (Ie34c07af9f6adb9e4b636dce3d0682c0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ib78d45cc282f110ed3ddaeb706a0fc12 ;

Ic9c2f173881d25f8976d723957809f51 I1f1684e97785eb48b33bff508ba4f2a1 (
.fgallag_sel( Ib869a349250a765d2f8660e0dbdcf312[fgallag_SEL-1:0]),
.fgallag( I0f5d081f9846ad888eac13d4916f5b8c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ief11c4434035425db82902c38e47be48 = (Ib869a349250a765d2f8660e0dbdcf312[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0f5d081f9846ad888eac13d4916f5b8c ;

Ic9c2f173881d25f8976d723957809f51 If3d55d4971a02fde1f02a4bac705f901 (
.fgallag_sel( I1a4fb631fdc7b5454c266589962ff5f0[fgallag_SEL-1:0]),
.fgallag( I607bdd63c3ee70e2721de3f994d2923e ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I1c3a6173bb59263a31998a5a69aaa38c = (I1a4fb631fdc7b5454c266589962ff5f0[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I607bdd63c3ee70e2721de3f994d2923e ;

Ic9c2f173881d25f8976d723957809f51 I9ee458d02fe4b8453ed5c0c58cb12b8a (
.fgallag_sel( I9de4e0e86e9edcf948d9eddf0401b94a[fgallag_SEL-1:0]),
.fgallag( I5453775d628c6c01c088278b6e090ddf ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2d77f481539c1258b61c2a6ca7208455 = (I9de4e0e86e9edcf948d9eddf0401b94a[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I5453775d628c6c01c088278b6e090ddf ;

Ic9c2f173881d25f8976d723957809f51 I32accd4e82357e8dae06d15e6f5bb7ac (
.fgallag_sel( Iee7b4838986c962969c00a0bbe53ce0b[fgallag_SEL-1:0]),
.fgallag( Iff51257cd95c2f3a38c64ae872317410 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ie88dbc3340cd953d819e7fa12d1fe3fb = (Iee7b4838986c962969c00a0bbe53ce0b[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Iff51257cd95c2f3a38c64ae872317410 ;

Ic9c2f173881d25f8976d723957809f51 I2fdd2d0fce79203f0eba35d81ea12805 (
.fgallag_sel( Id81b11a8ca1dd8989e36cef637ae6aab[fgallag_SEL-1:0]),
.fgallag( Ie5faf4f522c8d24bc2d3725be57453e3 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Icad54aaa6f380f2808749db56b76a959 = (Id81b11a8ca1dd8989e36cef637ae6aab[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ie5faf4f522c8d24bc2d3725be57453e3 ;

Ic9c2f173881d25f8976d723957809f51 I63a611b4c490a11cfc891ba79ea3e2b9 (
.fgallag_sel( Ibe96deab015b799fe7f69bae8432952c[fgallag_SEL-1:0]),
.fgallag( I7952b4b62af35c930dcffe35b1629100 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign If41dd08de4b2e28dae0404832fa0edd4 = (Ibe96deab015b799fe7f69bae8432952c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I7952b4b62af35c930dcffe35b1629100 ;

Ic9c2f173881d25f8976d723957809f51 I7a3efc8e0b278353ef0a94ac956c42d9 (
.fgallag_sel( I986b52155cc1470299321a4933241ed7[fgallag_SEL-1:0]),
.fgallag( I47337a0b371f749c3f7f5118362c2301 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I161c799aa59a0d82ca4db2b7b0293fdc = (I986b52155cc1470299321a4933241ed7[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I47337a0b371f749c3f7f5118362c2301 ;

Ic9c2f173881d25f8976d723957809f51 Ic619667eb623b8deaed02e3dc2ef9ea6 (
.fgallag_sel( I04be63a04f3942ce749cc9bd7540e055[fgallag_SEL-1:0]),
.fgallag( I21ea597751b3243936aea7c07cc90f70 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I911555064a463cd6a7ebdb4de801b8fb = (I04be63a04f3942ce749cc9bd7540e055[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I21ea597751b3243936aea7c07cc90f70 ;

Ic9c2f173881d25f8976d723957809f51 Ic65fb4662fd9c90ae7995ecfbf755d69 (
.fgallag_sel( Ia7adea5b0ec86e9fcd427a5468d72b64[fgallag_SEL-1:0]),
.fgallag( Ibdce05e98adef0314000dba3c482ace6 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib2fce59707fcc6d804b748678d3fa03a = (Ia7adea5b0ec86e9fcd427a5468d72b64[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ibdce05e98adef0314000dba3c482ace6 ;

Ic9c2f173881d25f8976d723957809f51 Iab78edd07ff3b17736ff42fbd54ff6d4 (
.fgallag_sel( Ie8990d8abd23f8f9f79d7fe38c57fa8c[fgallag_SEL-1:0]),
.fgallag( If0dbc84f59311eeabfb57b5fd0c3b632 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5d40a4f6c096b4962285bee680a366c0 = (Ie8990d8abd23f8f9f79d7fe38c57fa8c[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : If0dbc84f59311eeabfb57b5fd0c3b632 ;

Ic9c2f173881d25f8976d723957809f51 I2c0523be42b7ebb5765b2bb78fa1260f (
.fgallag_sel( I9d2f90ddddbdbb525d5f070f32546b64[fgallag_SEL-1:0]),
.fgallag( I74f2e7798a8383b78a5e7b816c2370af ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I692db6abe25b064802b76618cfd8d151 = (I9d2f90ddddbdbb525d5f070f32546b64[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I74f2e7798a8383b78a5e7b816c2370af ;

Ic9c2f173881d25f8976d723957809f51 I43edee0c8658a3feb993056f28a691f2 (
.fgallag_sel( I905256d73bdb63bf860e15687350795f[fgallag_SEL-1:0]),
.fgallag( I58ee302a3a1faa2b44d9052bffbc2a03 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I396539ceb8b33c1dfe096f71954586e7 = (I905256d73bdb63bf860e15687350795f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I58ee302a3a1faa2b44d9052bffbc2a03 ;

Ic9c2f173881d25f8976d723957809f51 Iad4036ae1dcc88bb2ca7f3e872c1d7e6 (
.fgallag_sel( I9adcfc18e4471209edbe9a379e996067[fgallag_SEL-1:0]),
.fgallag( I979a71fc0942bf62c06405bb63a717c5 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I4335c153299e851249a1492c14987447 = (I9adcfc18e4471209edbe9a379e996067[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I979a71fc0942bf62c06405bb63a717c5 ;

Ic9c2f173881d25f8976d723957809f51 Id9715c339baab9b2009c99139fcf3bd2 (
.fgallag_sel( I3d7d048348bf833f744a9f73889b7802[fgallag_SEL-1:0]),
.fgallag( I30be0ac758b5a0fbacb1c51a36ca8a73 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I5d81087b001624992357f909d2d7e9e2 = (I3d7d048348bf833f744a9f73889b7802[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I30be0ac758b5a0fbacb1c51a36ca8a73 ;

Ic9c2f173881d25f8976d723957809f51 I67e8b6d4723e8d1b75ba3309d518d694 (
.fgallag_sel( Id619e8d4040014d0e415ff71c5e0591f[fgallag_SEL-1:0]),
.fgallag( I9c50e0a8a01aaed98ae54530d5c76ba1 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I2b8539d21de88ded1152a26741003b99 = (Id619e8d4040014d0e415ff71c5e0591f[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9c50e0a8a01aaed98ae54530d5c76ba1 ;

Ic9c2f173881d25f8976d723957809f51 Ia2fba685f0a146057648e36cb4e11506 (
.fgallag_sel( Iaf3de2ef283e03dd72002026e1299224[fgallag_SEL-1:0]),
.fgallag( I0daac80ebeec26e428328344a398ce57 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Ib5f0b838019cb6c583e7aae384a7ffba = (Iaf3de2ef283e03dd72002026e1299224[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I0daac80ebeec26e428328344a398ce57 ;

Ic9c2f173881d25f8976d723957809f51 I4eef322451039cc1003bd4f4f51a6364 (
.fgallag_sel( I64551529c0028ec145407be7f5dfef71[fgallag_SEL-1:0]),
.fgallag( I6739f13ea431943bb5bacb4a05140063 ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign Iee7fb9e4ff68c15395c13083bb14e8af = (I64551529c0028ec145407be7f5dfef71[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6739f13ea431943bb5bacb4a05140063 ;

Ic9c2f173881d25f8976d723957809f51 I47dec328c368e176b4229850c113cfd9 (
.fgallag_sel( I5ebe580a943b65fb16ea722ba101fd05[fgallag_SEL-1:0]),
.fgallag( Ifa0e560fe6445b006ab74096a807b90f ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I18176a5b74de8d98a21cbbbfd35b0bdd = (I5ebe580a943b65fb16ea722ba101fd05[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : Ifa0e560fe6445b006ab74096a807b90f ;

Ic9c2f173881d25f8976d723957809f51 Ie4105e6adc5c2497769a3520c88146d5 (
.fgallag_sel( I0921901599c43b27e701758026dd3ee1[fgallag_SEL-1:0]),
.fgallag( I9595c0fd77d6a0610eb859dcd2b67d1d ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I033c58d2361a232bcfa2eda4ac665761 = (I0921901599c43b27e701758026dd3ee1[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I9595c0fd77d6a0610eb859dcd2b67d1d ;

Ic9c2f173881d25f8976d723957809f51 I633ef32ea8838c0fccb232dafe5c2e47 (
.fgallag_sel( I6033532f27c26b2d42bb3ea128f80dfa[fgallag_SEL-1:0]),
.fgallag( I6f3e685e70fa700b52bec62d0aed942c ),
.start_in(Iac11baea9832d6493626d2fe40fd385f && ~converged_loops_ended),
.start_out(),
.rstn(rstn),
.clk(clk)
);


assign I0ddecbd9a2e867e3bf8a447434f626a1 = (I6033532f27c26b2d42bb3ea128f80dfa[MAX_SUM_WDTH:0] > fgallag_LEN) ? 'h0 : I6f3e685e70fa700b52bec62d0aed942c ;







   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
               I18d11d94a39d5d7687736d266d3e1902  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib64114b4af6a37b3d52bd38cb83459ee  <=  0;
               I6b9ffa985ece553b83f7227e7a85141b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I06ed412c4554e98837146a5c7a6c4789  <=  0;
               I49fdba80df1c667dd264e5105a530332  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iefa11849e46b6ccd923e622fdb878315  <=  0;
               Ibf4fc04c9e0aa536a8e4b8a6192d8498  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia4245ce0efa56b1234283f4969246280  <=  0;
               I899abb7dcba235ff2afb410a87e16973  <= {(MAX_SUM_WDTH_L){1'b0}};
               I671b766473f67c92b75716e2bd9a9596  <=  0;
               Iab322f0da75316ca9937802a327dd537  <= {(MAX_SUM_WDTH_L){1'b0}};
               I24b5cce7252356b606027b301ac6bf48  <=  0;
               Iba0a4530bce787d70253a92c123f589e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2f0d19d012f0bd45308356fce1a50049  <=  0;
               I4475d6a1e59d35444a6a2d9647c6761a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I939c483ddfc18ee8dca73a1c98e6ec4d  <=  0;
               I217e2e1eb3404ba9ff06d284a18256b6  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ife63de208f77b322e1c885e78790f997  <=  0;
               I2003418e663144ee49f1ed044f6a0062  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia065f925c78015a3736219a5c7129439  <=  0;
               I4496255218b6d0f5374328803aeeb412  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie02e0e9e2627b178d6c54ea743b3993b  <=  0;
               Iecbb3f290db6dad3393b592ca946fa13  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib1e432e0b2d7979227d2cc591ed8e383  <=  0;
               I9f88e23f2a17035b31840356a5d0bfde  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib05aef46725afee38240d81738c673f1  <=  0;
               I3fd4a13843fc09ca68b827a8b09e6c49  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie7bea07eac0dc36dbce430e6dd088b5e  <=  0;
               I1530e79da3803bb87787397f19822dbb  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3f42e9b5ae0fc5c9315670cad33374ce  <=  0;
               I613821692bb99a8a6739d3c3ab7211ac  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie6f54d5d349ba8e19295a9ce17ba3f35  <=  0;
               I5ac600834d567934bd2f0b14a3c38ab9  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iab7ce2d8e89a5862f98bd812751d1d17  <=  0;
               I84fe1a1ecad408b16557957b01cc94b9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8a4157cd8206e66109f979bd9bde53b6  <=  0;
               I7d03cdddc264c89446cd80405c34d69a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5f0937deee06e2177807a6d0fbc2e2b0  <=  0;
               I5cf7e3cb90e84c3ac6a66fb6dde220af  <= {(MAX_SUM_WDTH_L){1'b0}};
               I598fa274e3ada377f2e7a43d7dfd9231  <=  0;
               I602c2e5bfa93cb3c87af70dd69b0375d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4a3da449219c7068a0bfd3a192d2ead1  <=  0;
               Id50fe525d660f0bb0ac3bbe6e68758f1  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia7a0522cea2126afdae3fb9f123d51fb  <=  0;
               I6a68067b177340dbea2c53f7d8bd5f14  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5d901ed468b60a31e199d12612a0b396  <=  0;
               I9efdcdeee8883d30159881f8831a2c03  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iceced38b8b522d1679ed4e1cad38c282  <=  0;
               I46290d63552b8cac8d22358cb38c5887  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7d3d6075ca3828a533b52dc3cac3a652  <=  0;
               I6435c7b1b3bfc5dae42cb1b3b03aefc5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0869d337e6cce62a05b29c5baa4ed436  <=  0;
               I63b2f1c2148e595a40bb41968e4b9a65  <= {(MAX_SUM_WDTH_L){1'b0}};
               I36ae963a57878d2c5b647910e003dea0  <=  0;
               Iafb6296c59c2dd241c880c6d57352617  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5851ca9a7e932378c2bdf2c118b498dd  <=  0;
               I0b982beca6221db7b3ec2afb3833a60e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia5597b68eb3f1c1d371cda63fa1fe034  <=  0;
               Iece8968796771c1ef094808823da8962  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icc939d3c403d238cf5c9c196cac91886  <=  0;
               I05c7cb4a076239b8976a76d418ad6149  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0bd90c7dbb94917bb46a3e008484f582  <=  0;
               I9076162e7b10bffbc9473e35b407e986  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6ec7620a49b53a8377767e363e88d471  <=  0;
               If702042844ed38f5e7103382ef4263eb  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie512ccdcaff0cc5c29277e28f1ba5fa8  <=  0;
               Ide63b2762649761944db237c8efe69ae  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia115f92bd6dcb4167f0771941a18ad59  <=  0;
               I1cec628c6d6e22895a0f0c0258851171  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7c8174a3579ed90c0ec89941ac53e287  <=  0;
               I46b0b74552e89df91c0027f0f093e1f5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7d6b68dbc5ac773ce97df3a6726c6836  <=  0;
               I68dbff67a1910346ddc0281b445f4439  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5045f1311d1e891577f3f8a09078fe79  <=  0;
               Ia42f547c0b02c2de66f2ff383ca1741b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I105c3326421f25d3b9931e2178c794d4  <=  0;
               If456045711d535cea07d9dd5ef9b04c6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I838c5c183e758ef4f28ad86d16befd87  <=  0;
               I9585ff28ce0f3bca71d582b1cb8937d7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I33c782b29a89c2ec375038b88919b564  <=  0;
               Iac3dfb28a343cbb391fdf58684e091ef  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia21ec0ad85852d1eea449283d1d45a7c  <=  0;
               I82650d4bf0a9b51e245665259f40fe60  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iae32e0aebc2719c3e476a5300f1bfdea  <=  0;
               Ib21e67aa9696222891a0b33c414b1bbd  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6914a92b8da6d6db6f2e8806c7efc5aa  <=  0;
               I1e168bf1a0dd18ff31d3560be00095f1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I60cad827424e4799360141222a80ac57  <=  0;
               I97e6d2bc8c1ad455f7c61de81e8d4826  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie3389948b5dd781ac9087e62cf93dd2d  <=  0;
               Ie1170db51d408ccc7360ce53c94a9644  <= {(MAX_SUM_WDTH_L){1'b0}};
               I566475d003c9fc40aebaba87655a0668  <=  0;
               If58c2c1e1dffe04295f3313595ffe319  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idb2467b1104f5b924d419208f2573df4  <=  0;
               I9a9fb4da9fdf5bd42cef32c7d8fa65d9  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie0a8d219223bc68ea3040cbbd349caac  <=  0;
               I785e4a1f2556289db0bd024e429bbd3e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ide01b9dcf3a3019d689d79f4d7ce0f32  <=  0;
               Ib6ca0cbcbaadb956d19a482fc099b175  <= {(MAX_SUM_WDTH_L){1'b0}};
               If33bbe9993ff895a7bd07bb8ee4ca970  <=  0;
               Id52b94ae6662bb2137d8b9d53280bcdd  <= {(MAX_SUM_WDTH_L){1'b0}};
               If9a84cb15af69dab2d9e4ed921f4deab  <=  0;
               Ic3975e4171d618ba53e1569e4fc93440  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ieba9f76cfb4c1a8069e2bfae0320ab0d  <=  0;
               Ib4e0f05afd881adf14a5eab850c75a3b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic85dfb2e44272dea346bdb4352a88c44  <=  0;
               Ifb875d675aa28de930d889ae4d37b48e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9f0f8b22b39af997db900c486fc37a18  <=  0;
               If98948e5f60b2c3ba1d7338e24dc0df6  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iebc1dd048a5c7e83175ba1030a4bb587  <=  0;
               I732bb69d248d700bcfdb287932839da8  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie8340c2226ffbab8f79e95ef17594210  <=  0;
               I403a8ece76036b3ce6277435609548a5  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic7dcd6d9c98422e20947712d0f4adc62  <=  0;
               I5a6cf1bdbcb2a342e548fb44c171aaf4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7df25ee69290c62782cd05715b0a6ecb  <=  0;
               I83a16a5be8d92896234bb9f2a36a22c9  <= {(MAX_SUM_WDTH_L){1'b0}};
               If904894b9cd6236c35bd9de268fab07d  <=  0;
               I6cad1cb66561eb6f0e3bfe5070b290c2  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5b890a24c074e7f2ebfee20ce4e15951  <=  0;
               Ia50c447d5838d7979b2e19796be6221b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I22f4468c482ed815d200d72ac2da570a  <=  0;
               Ief62ab0263b74086ae23a208da23e9c7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I091ae78d995382a96c68c47a60844a9b  <=  0;
               I564999dcc2f67c8f82fb5cd16af0ee12  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icbddf0d9df1bad66ea2f7352834bc759  <=  0;
               Ifb0e4775ffb73bb2533844db969ab900  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9a0db2b202a01aad173d2c8109cc596d  <=  0;
               Ib109fcaa55c3094cadb0c1f5f40ca752  <= {(MAX_SUM_WDTH_L){1'b0}};
               I724071f9e582e988d8f2d4c98ab9c070  <=  0;
               I56aeb1bd0b0e9857d9cfd2c6b347fe91  <= {(MAX_SUM_WDTH_L){1'b0}};
               I31e8ca0bb1f64410501bb3c55bbb60fd  <=  0;
               I02651642fc35059fe9b4141c2fa1f34a  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib7b1834c1a9867cb8f42c9ab177dc11c  <=  0;
               I1f1e04979c8a5badc8a103809f76dadb  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iaf22f59aaf7fa5f0e87a8d7504427627  <=  0;
               I19fe22e1104703ddc9bbc94a5368bbc2  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iea702a29812bf0e4b61cf21351648fe4  <=  0;
               I4386a95203c4fe83c6db7e25a288fc4c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I05fa85d0596e05c1df86434a2083c4e1  <=  0;
               I2ddabc0b4bc45698fdd877c93bcbe280  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic61a806c6bc223d2c23cf24dbf3e85db  <=  0;
               I5adddbf99d0d39c5d70ec6a0978f3ef5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8284c12f98671842255420333096213f  <=  0;
               Ia24d776498719aa6cfbdb5df69d648e3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ide2e42206ceb5cc9ddd1646dea75776f  <=  0;
               I038ff8eadf1c551dc42d09fbadaea5b9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I47512947d0532033dfa2b015aa107642  <=  0;
               I102dc8709a274d21c09abae1d2ac1272  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia5ec36569a57a6256966da94a52875d1  <=  0;
               I136256458e71d84e850b61a950f279e7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I07ea72a5755bd2b0da6e89389df44f69  <=  0;
               Icda6fe755f2d840f8e404d84b231e827  <= {(MAX_SUM_WDTH_L){1'b0}};
               I89b6e7810b2a5d45238819a6a171dac6  <=  0;
               I1f6cd53f31f27d86d78d5079e84c9716  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2e6141be9be5edab8e67a1e7f640903f  <=  0;
               Ia1f69042d447cb17772b29f634344b53  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib438d8ef5fdd32b2811e0e755acdfefb  <=  0;
               I84648f139f0fd470a62f0638aeee9e97  <= {(MAX_SUM_WDTH_L){1'b0}};
               I21cc09d0a95b4598c5614b7af3c6fe03  <=  0;
               I6ebc0ad14d76d3a80a4929ba8b5e7848  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia7a6617c92f999d7c19d3c338cc60e8f  <=  0;
               I26cba2d4920ff7fc40b1723c29ed8391  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5ea3e9e13e199daf8df53389a405cd0a  <=  0;
               I27980b3a1936a92a1751588f91a5f542  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5a202e3ec847e13fa21134123db7a027  <=  0;
               I5464cf638e0ca778d4e113b216084180  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie697e69bd62cf7bef4a4934843967cec  <=  0;
               I1804dfc05236c728f563342eb011f4f8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6979425ff99d598782f2a45b1d463f8d  <=  0;
               Id219264de5f6b67cff866b2bafc660b5  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie735fb63c3d40f44ede25d0a213847a8  <=  0;
               I03e4f803d4b82aa774662e02b188b0a6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2f132b8b367a5eb3d7029b1c27991dbe  <=  0;
               I32e079707d9ce4b31aea8fd2c998c27c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I55291a60dc5b1255d71ab749eaba0404  <=  0;
               I488f60405ded7af04c941bdbf55290f8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I804b17fba020affb1ed32666d73607ae  <=  0;
               I26d314b69785bdb0ca8cd52c258c3b35  <= {(MAX_SUM_WDTH_L){1'b0}};
               I478f85d129f1f538304e6cc74b9d2234  <=  0;
               Ia490437ab050e63e611dfb4d9366017c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I71ef5d9d9f272131a3c7bf864c0b4863  <=  0;
               Ia6cc50c8b7f83dd80d7058eea40338e9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I65ed551a24cd36ae20d1ffeac42fb99b  <=  0;
               I3652208cee3ca6dcdef63b7df53e4329  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4c99cb1e56179799079d9a484edf2a02  <=  0;
               Ia9a4760f6a2bf8f8f660e2b0c31dd823  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibd985ec8f6f4eed7f14ae2692367cc00  <=  0;
               I5ec267a535ad08c629940d70c61894a5  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic7eb65782a34589e2b015442172d7568  <=  0;
               I17fadd913ac1008fcbefff48ad366d8f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3bb60f8d4ccc5e40e97af6f6718c90c9  <=  0;
               I275728fecbd15ba77f57860bb329da16  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib109c4220b1113561ec1319a0ac74498  <=  0;
               I8d0bc446761559f2188e78200eb0a895  <= {(MAX_SUM_WDTH_L){1'b0}};
               I91ec97b5793a453f81b1780157e12d47  <=  0;
               If9fc4683c2f0545e1f077541fd25da66  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icae10f8dc7273f91884f011b6a88cf91  <=  0;
               I1c8e7559160d5a1fe1fa0002cc414d1c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8b7efa4f096bf761a8df08d1a3f1b77f  <=  0;
               I059014ede8b9092d817c0aaa1c7ed388  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib0dfb26e39fd974f64d54a0f9c0cd552  <=  0;
               I6294fc2c9181871210e0cfbb9834c3c7  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ida3a51bb8109fd4c3e494b736889efaf  <=  0;
               Id24dd0ede5504678fbd809ffbacd0dcb  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6a47d611882f8af53484f22ce5b74fe6  <=  0;
               I496994e784eb114337ac9e78ec0c4d3f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I52af26697dd18d51e902642e19045d9a  <=  0;
               I44c28351f261765c28a066a581c27c13  <= {(MAX_SUM_WDTH_L){1'b0}};
               I38b0b02379864bed0b097754dac42dec  <=  0;
               I84419e016619a3a33224eeaba85e68b3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic3f80e7837ab46f58cfd4b6c775d4e72  <=  0;
               I67d114d975d5d65f575bbb8c819fa22b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I87b9dff79eb8389488e97e427d59d767  <=  0;
               I6a452adc2501774b55e5fe73c642ea26  <= {(MAX_SUM_WDTH_L){1'b0}};
               I44926d094aefc5aa52713fb52704f84f  <=  0;
               I33792929f4428ddf0629231288e459ec  <= {(MAX_SUM_WDTH_L){1'b0}};
               I57127b05215e4faa4e32d5ca38611eb2  <=  0;
               Id0013f18ab77416e08d994c360b13473  <= {(MAX_SUM_WDTH_L){1'b0}};
               I79aadc384d50af92ae1af6760ffe3b3b  <=  0;
               I5683f67c7d462c01c55b8be9b6d1fca6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I28effe4aa10b24a221d5e1c84f2c21ff  <=  0;
               I4a5e3cf3066a4c2f7f5f8dbe824ff88f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia0d7cfa22522e5b4f7b545aacff7fa59  <=  0;
               I93879adfa4333a80be696d846e34d799  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifdac0b0a75dfcc09291fd95e842e68f1  <=  0;
               I199e944b303446e2cdafb6f34d0d12c7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1bbd0d48cc6bd8a4d4d520d38798f74c  <=  0;
               I91d282de42df72b1c439fede384d6336  <= {(MAX_SUM_WDTH_L){1'b0}};
               I06ede5ab6bc97827c4f866dca1aa17bc  <=  0;
               I8a06d2c278af9d552fa36a61128b8a9b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4b7f22e0b9e1589fbc1d558b37cceb37  <=  0;
               I5a36e45af7599ec00703dfc81f9d1176  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6e63e4047456268e73ad16a5cde93681  <=  0;
               Iae09429ca8733186fdb3c50f36895746  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iec7997b0018f4fb3572579a5bf1e4728  <=  0;
               Ie5f74b33d06ddb8b32b57c8c82392001  <= {(MAX_SUM_WDTH_L){1'b0}};
               I11cb6032d99f05b3f908418a70fd3d6e  <=  0;
               I7d3cdb71cdab3a85122130207d872476  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idba56a073e34e530c36025914f7646d9  <=  0;
               I68ae9f2a14b161c940f6685073eca97e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3a7582a1c86f2b49979372132ce98c87  <=  0;
               I778f907b5eacdfac02b0bc4547af4ea3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifaed912ee00082f8458ae37bd47179a5  <=  0;
               Ibcea5bf1e21fa764ac9f2d2702c8f79a  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibecc30f33083404bf48eb0005e14bb83  <=  0;
               I93a3e1a8e414d4775f19c0c9f16d07a8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I87009d289b53c6e366b73e275e414caf  <=  0;
               I8772034840834e51187950d320f9eb40  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5d5b08cc3fd13b96621143655a806c7d  <=  0;
               I3d0aa00b61d4684ad46f49329197c901  <= {(MAX_SUM_WDTH_L){1'b0}};
               I94ce074b29f44c5e4a63ff6e00d2b9c4  <=  0;
               I146866a6d46604c47d87afa3c88308c6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2fd3e923d1adff22ef7718dae5632b29  <=  0;
               I84cf7aa78617faed2f1762bb1961cc0e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibe2d184a52eb5d33cac0ca4a5dab55f6  <=  0;
               Ib1f43a0b9c86d236b2ed71c35c296b9c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0907dde542619e162f45f3dac8c0c16f  <=  0;
               I88aaa7538f9007ce204319ec639d1c7e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9bdfa0d38ed6d215e7ef7ecb12185b60  <=  0;
               Ie3a171564602e9936d7960e83bb0fb3a  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie0e096809efa587a070562473e9a2fff  <=  0;
               I732b452fd9521b3a13ff1f965c443325  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8c2c0b7861868365bc3935ef8d0fe309  <=  0;
               I16cd75fd747b600e90763d8ce9c08210  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idde6e2f615f8ec0aa66b7397e5581651  <=  0;
               Ic6a7d6bfb12f40ae8823db716cfe017a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3098e45c14ec08213883f7879c30150c  <=  0;
               Iea38a3c260d0caae4ae042264a0f4787  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ide3c2fa1d5da990a0566c65a12d1d7da  <=  0;
               Id6240152bd22a9655b18bdfd91812e03  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6ece8c59f986da73f00e104ff5966189  <=  0;
               I07eeb34c9dfb9baadb9f263b6f095ecc  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5c002c1ec0c63a2c04ca2711fde50254  <=  0;
               Iedb57db3cbaca9f9a469d91ed81466a8  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icb5a521ae9f45d8c9101fdde8925e64f  <=  0;
               I2972b771a4e99ddfa2178349a805b16f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7b72bfdf546647380e6b1f9a810fd1d1  <=  0;
               I6a61cdadaf987763080e6ce4d1605ee6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I84581a99221f2aab1e7cbbcc80296ad4  <=  0;
               I12e430f1ccaa6099ba9ff803c85d9532  <= {(MAX_SUM_WDTH_L){1'b0}};
               I27d48bcfb04bf11d76b496d459ee1b48  <=  0;
               I2cc3c84149c81572357c01219248aa3b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib89fb8b901f12120ab0bdff5207c74f0  <=  0;
               I6d4b18dbba5c2b058f93a8d46bed38ec  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic2324007897bedbb70a77faa1fd301ef  <=  0;
               I32ca5d01c39fe736d6ed57d70fcbd555  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic75af8091015d4615d0c059ceb16371b  <=  0;
               I8807f2f633d64cb064fbc149ebd30412  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5b98fb653fa4d3d4ce2ebccd24085f95  <=  0;
               I822d3b3516499e58ee7777b99259a206  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic9320f9ad332f511422f5b805de9488a  <=  0;
               Ie706bf8dd49322fc1d5d83e40fb20f04  <= {(MAX_SUM_WDTH_L){1'b0}};
               I71574a4f01fc2e2fdd051a90b9115524  <=  0;
               I9975f2ca851119d7ec85cfdefda150f0  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia59c01c2e6f19ee93a091dbd1a1da83c  <=  0;
               I2e0639bf4e48a7b1486beebcc9ad7c0c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5e8e70c7ad583c0c4f09cacb60602c00  <=  0;
               I6131789039de7dc431c3b9b59ecb7654  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia180d785ba74d63500c25e3a04d21c03  <=  0;
               Ia20482fd064712397fe2f9f77f4d854b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4dbcb057b2076d4efd4e05e818d976c9  <=  0;
               If052875ec5a78a68428a1ff09df623df  <= {(MAX_SUM_WDTH_L){1'b0}};
               I24e240c3d018053712e0fb7f861acad7  <=  0;
               I2e27abc9297a3fa647f50859af7cb094  <= {(MAX_SUM_WDTH_L){1'b0}};
               I78d4209646fe0f2b8027988024b947ae  <=  0;
               I5d5e3b64ed1ca16d65d8eadb8100fa06  <= {(MAX_SUM_WDTH_L){1'b0}};
               I62fa50cc71ade42b52be1de668da6b7b  <=  0;
               Ie91a08b49b9bf23270dd3fa331e64968  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5145e1005293c49c849599347a4a2b46  <=  0;
               Ib599712a1e8fadbdf7e3712bca6c0b74  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id77a6df77f3d714b6b1f60bad2462f2b  <=  0;
               I1791c009b0838ef10233015f80a5c4af  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6cbfcd474a5a76538db10b8c3235986b  <=  0;
               I3dead2d8d18ea8503a578469625f3aa3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I17c80f6af6d201a1214d251778a9e534  <=  0;
               I2fc47140b9df2544d7ae9c82cd38ebd6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I468342d7ba88b0a9313f38d0ec2a81e5  <=  0;
               Ice09150d69c67cd2d08d6e63b8a9bbc7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I189be0be892f48991d69acf5a0d42533  <=  0;
               Id67765c4a6b11f6ee0a4524ebb2d1ca7  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib5bdc1c490d7d2fd11359fc6c79372cb  <=  0;
               Ia17bbf4b7f063de0bf0701276b7b0c20  <= {(MAX_SUM_WDTH_L){1'b0}};
               I85e112a43fa9046e94da6bdb7b3a13d7  <=  0;
               I9f9075a7745d475331f0b25bad830421  <= {(MAX_SUM_WDTH_L){1'b0}};
               I03ad487e845cce369a813b0c7f32e59d  <=  0;
               I4d832ef88af4d4244516b0bdfd2b461c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I85aeb073e949fc999464ce61479790db  <=  0;
               Ib2038174dd555b1d058778fa904aee65  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7534524f9d9c64bdf0bb88ba351b3ca5  <=  0;
               I959dff5d57b4c2adb85c3602d5874c90  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic4a902801adb86fdb2481f5b868daa8b  <=  0;
               I30dd112c5a6793cf37bfaaf8dfdebcaf  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1141271b2c1fa529b7f4e4ce9ac10c95  <=  0;
               I4d4a0930420b4d7da8b6e91b2b25bc51  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie62709fd754ca31b0e5d830901bd6433  <=  0;
               I7ae1d318fd0df386e0c8bcf0f0a94e4b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6c6a99a66fe46ca1532fa898123a6131  <=  0;
               I06cc62e12d5a261d672b5428dbc9767b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I963a6698cd1f83ce4e7ecaff7f53ce25  <=  0;
               I9798b16b4658501d739d46182d7ab169  <= {(MAX_SUM_WDTH_L){1'b0}};
               I451d9f14e13b272ea041178627ef7f56  <=  0;
               I90bc85b7a6e56250bf13407ddd32bf11  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3e7f571589d773eaf3435c03bd13c9ca  <=  0;
               I88990d32bd34da606660f1c078b36ce0  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie823a06acbb6935875c5cb9088389b27  <=  0;
               Ib32ce57f2840a45fce8e66f71b37719d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia4c876fe77f09258fb130d03b8cdc67b  <=  0;
               Ib0179c2048d6c9d1865d171b48c521ff  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie6bf8e5060074ce2dfcf7ddcbb158bff  <=  0;
               Icc8ffcc0641f0f9405590338e6b5e517  <= {(MAX_SUM_WDTH_L){1'b0}};
               I706ad22942f1cfbfae4fde958450189b  <=  0;
               I5d6cb688ef094e1f119d8536f0f56766  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic64d1cde239aef0df4f227a64762f9f2  <=  0;
               Ia5aa7c66d2818982a661e4d048876d1c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I719f60bd29522fded995c8230b4f3a34  <=  0;
               I449e514b6afb3e8e337691fc64f7431c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1bd8505e6f316488bb1cdd74932c0314  <=  0;
               Ibbd5f0906646560a903abcf6848ee80e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I63e645f447ddd1fc9409879872479bef  <=  0;
               Iee607ab8132caf0f678324d20394f533  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia8298013e67424c2d5fbe03634170080  <=  0;
               Icc90fd3c992755ac7e4aec1370600e06  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib404a1296714f45ddca6351a918ee875  <=  0;
               I81e0ea92e07ed7d29b4ab769443b55d3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic08905e9ffee26c630277db86cd5be95  <=  0;
               Ie7554e9d2bb6287b440973a9effefb50  <= {(MAX_SUM_WDTH_L){1'b0}};
               I674e937c017f29d18946139b00db02d8  <=  0;
               I3fd483389e4ddb927e7be7636441f0f1  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib3f5f61eaba0c2dfdf6c75e46e4233f0  <=  0;
               I3d7a6bd63d9f66b068c08cf9046474f7  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iff1039ba558287ef96daa7dfd15d6294  <=  0;
               Ifdb5bd8e8237676fd8d2816bfa53f0c0  <= {(MAX_SUM_WDTH_L){1'b0}};
               I017268444024bc19b209dbb4322de15c  <=  0;
               If2865b698bf9c511fcf6724856074335  <= {(MAX_SUM_WDTH_L){1'b0}};
               I22e4741c472c64c846742391d81f682c  <=  0;
               I077ad1ef2fe0a7e791fdb45026788641  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie3c87a536250268b1012b6166173108b  <=  0;
               I4c67ed6284da547b599a4602a3cc51dd  <= {(MAX_SUM_WDTH_L){1'b0}};
               I54204328537dbc383a3a03352e9d6fb6  <=  0;
               I3d0babc64a3400a1ee57fff14920d1e3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic5d81213c2d23b0549006ed162d9e6dd  <=  0;
               Ica1731833fd3d6a881b3a17a5916f7e7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0ac628860f9fb9e6daae572ff007f34a  <=  0;
               Id5705e57bc5c050342e82a302b73902e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2487101836608b77528a49d037c40fb6  <=  0;
               I4606e0ec878c615753206459716b5d25  <= {(MAX_SUM_WDTH_L){1'b0}};
               I99d49fb5c921d2d837ac7b02716d9ada  <=  0;
               I5ac4f231a175a60f63db8d4d71cfabaf  <= {(MAX_SUM_WDTH_L){1'b0}};
               If4d0af4a78a49e861adbdb1a3f6e7ae9  <=  0;
               I26a3cd9ec3a564df04ad20559039598f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iccefd72e7e22a425ced6974251245da8  <=  0;
               I26801bb91e66797982b66ce815da85a8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3fcc5c32415df9710be01f0f35ac68e5  <=  0;
               I3b617a013c15e8b623ad517e08df3a00  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0bf8339802110abb8bc94e481647f25f  <=  0;
               I65f5f9a3f7f68f4b2fd7695ce6bf4629  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6ae57b8d68417d1ea8ef70d43a943e0b  <=  0;
               I7d405b59e360b17d7f2eb1805b796fa9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I07dd0ed55fbdeaace398ab7644a5189f  <=  0;
               I033ad5c570f42830b265d7bf6a102757  <= {(MAX_SUM_WDTH_L){1'b0}};
               I69cfa3967387c5e8e48994b6466673a0  <=  0;
               Ia00376ef5aca6a428280f2dbf25ab1cb  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2ce599e7a40a71d9fe09f80269accc31  <=  0;
               I252b17144e39018fda208bd18b555c09  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id424746e76cc70f9292ed41659973621  <=  0;
               Idb756c313694457c14b02431f3f076c7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I45528f9be6a8f9a0f646d83223307e79  <=  0;
               I0c1545b312d755b14ee27b399a1d3079  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iabcd2910bddf2e544c707c553b2ef370  <=  0;
               I903842d13327b74a952be0aa6c7ab0e8  <= {(MAX_SUM_WDTH_L){1'b0}};
               If01521dbf7dd9aa5196a9130ba47b149  <=  0;
               Ic461c1b7bd09b59297193d388c525ece  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9284cc53534eaf3d6e5b4e9d9d93bea5  <=  0;
               Ia14490057ef27f5df5f1b23ca6440a65  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id5fdf11f0bf10ec37b11ced0a3268ad7  <=  0;
               I2d3c1e36bd952fdbe4fac5f3af07e666  <= {(MAX_SUM_WDTH_L){1'b0}};
               I36cc6827c8e4c7831078c8f9972ee78a  <=  0;
               I7fcea0a5f9987b2414ab443bd07c05ad  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ied6cdc5d7aa6335b2c32d8ab6ee6d889  <=  0;
               If0f5bf08d96033f6281121230c1e47c9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I70709dd8c55168e62143f56d0bda1239  <=  0;
               I19412627d5c573ceaa981cd7f1027e83  <= {(MAX_SUM_WDTH_L){1'b0}};
               I73ce9bd4312ce9a6cdc0c6b6aec72a55  <=  0;
               I7c72a1709b233f745fb0323d04bfeb1a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9d0fc48c488109406aa9cfef80ac3b48  <=  0;
               I2639cefc25ac6f4982e4eeccf8fa810e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie09336ee55ee45ac0297849f7b814f4d  <=  0;
               I76340f05f74b295583bd9353884979be  <= {(MAX_SUM_WDTH_L){1'b0}};
               If919b9778437e1c4366017968d1ea582  <=  0;
               I00974459262f29ec2b5472472e49faf6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I71cdff133cb7a645e623c4bf06588fc3  <=  0;
               I075efbd3c4d87df8d733f0b3db008b1f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie7fd0410103d16e27611f9ac30c657da  <=  0;
               If8bd6a5d380075f1ee7f7a4542531dbe  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iab93975104312336985d4736015098b4  <=  0;
               Ib81b730d107434503c988ab9f00e1605  <= {(MAX_SUM_WDTH_L){1'b0}};
               I564a4d4a94f9951d85287b2ac35479fe  <=  0;
               Ib05cffa1bb31054450391bf9e17f8ef9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I09c5b4146a3c48ae706d3041ddfe074d  <=  0;
               I627097c06e3be5a4385171f3ec7ae5c9  <= {(MAX_SUM_WDTH_L){1'b0}};
               If205c7d745e5372ea61afa389f1af2c2  <=  0;
               I76e2c6001e1ae97670539bd471fc74e8  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ief37a022c34d4e670413f5b7db306876  <=  0;
               I8b4433056d26f4aa60f18418b0114930  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5ac36d471eec2b3ac068a2d20283f674  <=  0;
               I99601176686afd8fb85a85ec43849e6f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I68acc6967dd156d6373abd6cc620f247  <=  0;
               Iad8276d5be3d9c6fc085465f05ac2aed  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic830033c7861645951982dc630e3385b  <=  0;
               I5e5dfce3ceb4fbbfce344bd471901736  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7f9305c8bfe731300ad0a9d1ece97db4  <=  0;
               I22ace766690e445ff36176eac2473368  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0bb61f163279dc993a94e647611f6e06  <=  0;
               I896c57162e4384f021d822789b4c01a3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib5effb1b2c147179bc8c8febce7657c7  <=  0;
               I3d0367a799090b3c9048235436a39063  <= {(MAX_SUM_WDTH_L){1'b0}};
               I81dd944eccdd3dd6fd84727d21efd0ac  <=  0;
               Ic0f25799f0dc7cc33de95e47ebcc083a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I986e7c899df08e35fa2347e282e8c90e  <=  0;
               I7186b368e297d0db1f746c6241eae65d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idb764022b3ae49281c7b82f6e309cca9  <=  0;
               I21d63f6fe5c72798aa4636527c02613d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I311eb64d22cff4b1424f3ccdd33dec45  <=  0;
               I15e0219f2da6f52177e76580198d0e6c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I128183dffb32a1461db0c2b851559f68  <=  0;
               I4cac308bee8801c4f9716673e39da4ab  <= {(MAX_SUM_WDTH_L){1'b0}};
               I817fbe1f44196264e2531197ca8da9ea  <=  0;
               I6f4f7b4e45a495fe139955e0605ff208  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3e74c445193a1c9ec9dcb31f4aef2117  <=  0;
               I79ae5f2981b7dd91141b0a22f012f4b1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I70f3cac8f36ef943672bbe7a9d6be5ed  <=  0;
               Id4b4d757e50bc2721e8725ae10d88c9e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I26b4d738c45246201073f4b4a786078a  <=  0;
               I4513152c34d5d00ddcc4f099481f659d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6c4f341b9eeda21a97806084196421d3  <=  0;
               I7bd4e77993fdd5a0833f1cdc7a382b56  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibdf325321ebd9a7baa25435537c159bb  <=  0;
               I13b0d404e7a96cd53147b574b242ef41  <= {(MAX_SUM_WDTH_L){1'b0}};
               I626a4c66bf0cca36dfa2bcd8c24bff35  <=  0;
               I4acc3bfa99b152c6ef6d11608f639b70  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icd6ab7be501038196ab2674cdf764453  <=  0;
               Ia1ec7ba972ec6f0049c4cf00b9d42125  <= {(MAX_SUM_WDTH_L){1'b0}};
               I31c6d68ecdb4d0a6790a12343f59731b  <=  0;
               I4fb5494e6f04e29d76bb8d3bc8bf6cd9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8eb06ffb6aca72c66cea97d9caa26f1c  <=  0;
               Iaffb0ef4e18bb7b582275b43684fcf3d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I35ecf6ebd98d91d12361beef01dadfbe  <=  0;
               Ia5e3649f8e32a81606ee34353c54350a  <= {(MAX_SUM_WDTH_L){1'b0}};
               If73961b42bf31d49c78c3fbe86f8d2cb  <=  0;
               Ic675cf7eac5ece436feb5a8acd642f6b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I560157aede2c2c3b6dce019e2fb4314c  <=  0;
               I71357943bbe307c9ae9099d4bcbff882  <= {(MAX_SUM_WDTH_L){1'b0}};
               I075a8e7435a4fbe97304b4d379bcfee4  <=  0;
               Ib2684f54caebb1a1c079a2a4f2cf0dab  <= {(MAX_SUM_WDTH_L){1'b0}};
               I09a1ad6a0fba78d4984fee238fd95bd7  <=  0;
               If19836577f9a254b365f0dcfe0ae55ce  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5c03de756d46517f2158e4ffb019edd3  <=  0;
               I2f47a00b58779b836c08b472d305b031  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia897f60b5c256180be523c5ff8ba6b77  <=  0;
               I8b2593fd0e35c37f68097187a41596e2  <= {(MAX_SUM_WDTH_L){1'b0}};
               I81a7d30b51b1d7f9d9bc9a97d2f3caac  <=  0;
               Ibbcdc1c30d3333cbec65d264890cf3e5  <= {(MAX_SUM_WDTH_L){1'b0}};
               If46a830ca08eeb2b8b3d8b2f996491e8  <=  0;
               Iec6e9640b0494777c013c97613855ce7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I13e6271176ef80d03f8878441893c467  <=  0;
               Ic10f396b52dda0dcfbf2a847cfed617c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idb5b4ae9bb42a053d9db8b8c71a0b9cc  <=  0;
               I94ebfb633f3272b8f40303ce768f0ade  <= {(MAX_SUM_WDTH_L){1'b0}};
               I96c6deed53888cfe0b1fcbe6832a1d61  <=  0;
               Ie975a6fd78adbad8b8a56bd6a3802e4f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibb40e3b624d2f19eeccfe071e540021a  <=  0;
               Ib852991e38422ba6de5e18a879ddc3f9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I93bd27a068e6fd416060bd5d919b3451  <=  0;
               Ife665c9aa6794cccffd04923f4359047  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iaf516c91fe1544bd0a6f671635eda05d  <=  0;
               I076cbc669ff4fb135ffc85910c888241  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6029a024d76e9357223c6fea077501c3  <=  0;
               I50245c953aab8c513b17b894afb36a6c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8dd3c6c27d8fea2b67906c78715c5854  <=  0;
               I33ac557ef59d79e8b1b359e499a00119  <= {(MAX_SUM_WDTH_L){1'b0}};
               I244ab0a87c282939527938b5d43c90e8  <=  0;
               I173fd30c1a5367b61e3fda352365f557  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8b9861dd9f6dbeaedffc07a3e088cf49  <=  0;
               Id6f5041043fa4fd352e74016c4e7de48  <= {(MAX_SUM_WDTH_L){1'b0}};
               I71c3dc98a45a807f146ec052c8a9fb82  <=  0;
               I6d863254c7f0b52f803b2af4b184f99d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iaa6c753b09c2244d22a8680d73670deb  <=  0;
               I1eeb9c94908cc9ddeb8e3904a145ec6e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id8e40a0bd35259f34ffc971eaa7f2fc5  <=  0;
               I6211e241282624fc50fb4ca1842ff9db  <= {(MAX_SUM_WDTH_L){1'b0}};
               I59df806ee758f4db794635ec24232ae9  <=  0;
               Iba09e22ece1eb1639d2bb940d3273fe0  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7bd8b1c89a39e4dccbde5c5e040c162f  <=  0;
               I2fe99e4fb8c660d83508bff50ab4929b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id3d37273d55ba1de64f97f6d11e704d7  <=  0;
               Ia73db0428763da3c0feffc94a8a8f4f1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4ff07696ccaf99e49d575694d3a2670e  <=  0;
               I6542fbca90e189048b15deaa3af5d836  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib89e0144bfc6be3be9a06a08e4f297ca  <=  0;
               Ieacf022fc976bf397946d6481468d6a4  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ife372091864d6ae9b770b69db66ff3ca  <=  0;
               I1cef7e6e0555e076b68bbc57de8f289f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie81b8b84cc2795e2e92168bfa496ece4  <=  0;
               Iadaaac832a1422494d4206edee770d63  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia6eb1062be96666c061e5fc1f830e1d3  <=  0;
               I905b0ec8983ba423798bbe8282728af8  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia0947c561ef360d78d0dae68baee6161  <=  0;
               Ic646b82fb6e3d0afb3a58c4e0d68f06c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3cd67e0abb8ff03aa1068dcb61aa3468  <=  0;
               Ie57f41c62e23092974664f967a27566d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic64779388389bf13a0e5240613caefc7  <=  0;
               I34524ca1dddbeadcc060954238175e7f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I767cd611a030d15fc5eebc6e1b9ea2dc  <=  0;
               Iaf2a93993f99814321951a6bffd8bdd4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I03e14765645af77dd39ed51320bf7a95  <=  0;
               I97e4f7a9a8a42be813c6e4128936df3f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I29e966dc25c12cd095c25c5e6fd6d872  <=  0;
               I682a67100f862bac0155a870cae0528c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie8b68c8c51e2e03a3797a2ec3f8a56ae  <=  0;
               Id5296b03b99bbf52d3ec04dddf3e84b1  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibbcfb7c284a2c99332d9261a4de199f1  <=  0;
               Ibb089d47014f9002f2ea6b431156d9af  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3e33a1f3e03bdb35d7c03f17f4ba4ebd  <=  0;
               I83496522139d35aa028dc9cb8a78d442  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0f81337862e31b6a4a6db462533d17f3  <=  0;
               Ifd4ca5a83fa0c09b043ad54d25971410  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5029faffc78b92bc6e76d08fc4cd822f  <=  0;
               I6efbc715be55b616551a7d4650a446dd  <= {(MAX_SUM_WDTH_L){1'b0}};
               I11262f431003b344ab224ab5488995c2  <=  0;
               I572bf74835f5acdf5a17de2063c293fc  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3f0fc144d868b4446b6d261b3ac80a67  <=  0;
               I5f8194ef67d22bcd38f415fe8d9a6ce7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I463736cac698d2366442abf5fba61580  <=  0;
               I3d3f2dff1f64ce14071e5f315bb8a57f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6cc14595c5c11f3ef8daa2a0b0634f73  <=  0;
               I8e3880fe0374bc068ed14eeff9f6d009  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia2345aaec32840b490d4b58c6ab3f115  <=  0;
               I51d8f49653c7468b2923390dc5932a2a  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifdca49a87cf807777f2e460bd3d3a4fb  <=  0;
               Ibeb380f8f935c8e061fe00734675662a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4fab81c713b53f66f545f4f614713462  <=  0;
               I641f4280286c9343b7ce001a8b43fa21  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1dd4557e3f4df4fa18a9198f9f36a98c  <=  0;
               I796970d7c73d8fbd7d25793d0dbf9872  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id2ac1ca1ab4cb5eaba4ebb9dcb31d857  <=  0;
               Ied0b1d10ae09c523d1cd1cd3e5b184c6  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id40872fc0d4f1e9ce25d366069af2f1a  <=  0;
               I7d0d39d94d929741158c39f69e8169e4  <= {(MAX_SUM_WDTH_L){1'b0}};
               If3b1c8b7c2296e5664f105adc761fd48  <=  0;
               I2349636f6ea8796c7b798aa555641a9e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idd694db68c0f91155fd81a106d596d8c  <=  0;
               Ia3739201eb91605fc115bf320d4c24f0  <= {(MAX_SUM_WDTH_L){1'b0}};
               I89473d1b100eb64c951e986819a4bc59  <=  0;
               Ic74cc511acc98510da011e126edaf3a3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4351f5987566977330a1e69b78d4e6aa  <=  0;
               I89b1312c0696711956ddcf787e37f3c9  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic067d44971ef80f6c63c6e187a583e3e  <=  0;
               Ib2ef1187c1743da2cd83eb9231a7ddf1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9d46fd2fca52ea2ecb6242801a4378a3  <=  0;
               I21710bdb6874ab83e2b2a2cffb026ab8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I916104565afa11bfd9b3ef53551ade1d  <=  0;
               I2ec8afd22c84596550412a5d2c7129af  <= {(MAX_SUM_WDTH_L){1'b0}};
               I48812dfaa796a851f23d230227be8969  <=  0;
               I57056cc2fd4bd1ea6e980cf90c22e871  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia2d3db44f16c9bf381145ce71ba2efd2  <=  0;
               I233becd31032d63e65371119edb2cf79  <= {(MAX_SUM_WDTH_L){1'b0}};
               I849110a991c42aefaead8d9500a18912  <=  0;
               I0142623400f5994f581a4797fd9d327c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic4988fc07458064e44f882807bd13c4b  <=  0;
               Id3e298c9f2709d8dc01c18626ea846e8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0fdd344f1ce42003661bb06c2c0d2fb5  <=  0;
               I1044e090bdf84a1bd30438137d6ed056  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib2ab217127041c49acfc86ef2eba3350  <=  0;
               Iff0f43c1fb40bdb3271a3a38d89f4d6d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5d6dfd14a38b207a97ba02a357965d5e  <=  0;
               Ibc71a0c3641097c144513810bc9a0a7c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I963472efe41928bdcd4c87ae5d6d9781  <=  0;
               I6ef3b025eb065f833efe6daaab699efb  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id8cde19539c6cdf7186230e34b96dc15  <=  0;
               If76152e9435e7300b19095a9b070e0f4  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia31ee8ac9735d3bd38298fd5d9812aa1  <=  0;
               I5fa63303ab85db9c8cd268528eb604ca  <= {(MAX_SUM_WDTH_L){1'b0}};
               I79bced0e80e2554a4e748644c5985896  <=  0;
               I69d6adcd3d35a24b393e97ed6a99c061  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id0216555323efdec39d0448568f59f23  <=  0;
               I8980eca0e5973840121576b6eaaab736  <= {(MAX_SUM_WDTH_L){1'b0}};
               I35c6735d2fa06f57341b6010f5bb825d  <=  0;
               Iadbb5c4f7b7c02e151d5118a7ede1f0b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id2e8b17327e8c85999d3d6b3dd31a164  <=  0;
               Ifff90bff22a3bcc33261004136d2e655  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iccd9ca809045617acea3364a6c86fde9  <=  0;
               I8d13628f322640414a4b556ee48d3bdd  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8ce27f01f84ea9babfca8074bb57417a  <=  0;
               If7d187cc56b1014b1582c5f5b94759f1  <= {(MAX_SUM_WDTH_L){1'b0}};
               If6bad1b3865cb4cec97a730043863b3d  <=  0;
               Ia01d5a33078abf4b2d6c625af01c25f6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0c88089ad1c5fc9928c091c1c677ca66  <=  0;
               I4c74240688b5635b5323ce3a8ac666fb  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ida2ed38c156200b9511c3b4515f42e5e  <=  0;
               I943e9afa0dc80fb50b5869cf34726823  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id322e4a2b0197e5b0f67a220134ca540  <=  0;
               I44d8779f30245bc7f1475e6feb762cec  <= {(MAX_SUM_WDTH_L){1'b0}};
               I935862d2f7c82e05768f55434167ba47  <=  0;
               I479e7456c445ad604ebc134872a0fbfa  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1c6dd243cd7d2b8d00eb59e2ae30331c  <=  0;
               I484f372e3a2e74e0791b06aa666b781e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8ab7b4e7f78fa63ec77224c7e5a31198  <=  0;
               I64b07241996c48963595f28e35a75be5  <= {(MAX_SUM_WDTH_L){1'b0}};
               If20d6cdf73bb1a925317f35de01b6f62  <=  0;
               Idf678798bf4e1cd316a49a2b413cb29f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8c2bc7a3c5c7e798a9dbd0199d37bfd5  <=  0;
               I35fd5e5e93f992ef5ff6b11f9d69609c  <= {(MAX_SUM_WDTH_L){1'b0}};
               If814b033c7e3229ba1475b305fe98307  <=  0;
               Ie72397edc1c597c0a8213b67a030a482  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6e69f6d33a933441458f5a46decc4e8d  <=  0;
               Iae50178e99a07cee0eea6f7cfdcedf1f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie2bb4ef41cf43cbea46b7a6d492bf03b  <=  0;
               Idd7082c7a65d7f8e0ea88142312a631e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I757b0e2104a4d9913cf6b3a13ad7d6d6  <=  0;
               I4b580dc4cfac9e9315d03b60e2a915d9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I46c7f4a6ef4b3ac3eb74b4ba2552fcdd  <=  0;
               I77cdc9841414221c3f6c3cf35397059f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I247479fee56f209f758feeb4770e50de  <=  0;
               Ie59619c3e78e616e1febd2db2fa940ae  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2ada4b104b94c163f3d9201808d21121  <=  0;
               I5bc8079a5896f59bc6137b59c4b7e750  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic7f0721d5160d4ce266b21c53aad0b4e  <=  0;
               I239bf978d991f702ad23bc6b4b8be1dc  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9af70dd16bd606c4b9588ce32ce9844d  <=  0;
               I450351fbb31246b49cfb2d622b9e90b4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I30c5fca5bab3bc9cf5c024c3302bbdbd  <=  0;
               Ia7c17a0979f3bbb9e9e821bf69a239b7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I09db79951c2115c2db0a3036bcb2b63f  <=  0;
               Ic22975c34b92a39bc8940076e80d3c0b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id76636b29db2c1a69d585b68731fc3b0  <=  0;
               Ia7be8cf38ecee4568a939cb2ef727619  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2ce42f5733f4d0cf15d1a7944fe0344f  <=  0;
               I3e475cb1733d494f5f7c4b26a07d5852  <= {(MAX_SUM_WDTH_L){1'b0}};
               I87e7191f5ec3f0847afbca81660a7608  <=  0;
               Ib2c0df16678f6aac19f7af4ad4e53ef8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0f8f4304c88efcc90c021be7764be01b  <=  0;
               I8bd2ef39eeb7089409db02e3806956ac  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie8b6b834bdde210d6f7a3e60fc78275d  <=  0;
               Ie3669e34cd19462f524932b3d232b546  <= {(MAX_SUM_WDTH_L){1'b0}};
               I591b99ab1b55e2eb4c10996efab5e0d0  <=  0;
               I1ecea23a4e56948365dcb04c5bf6d6d6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I27402f7d7892626f9b5ea1fc39987c23  <=  0;
               Iac222e9e39e300d7161ed05153cd9ca0  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie6e9475310530f511d38602f2c58a28f  <=  0;
               I292683f8453be58f65370a286c1a4505  <= {(MAX_SUM_WDTH_L){1'b0}};
               I30eeb2d396c381acb08253d886025fe1  <=  0;
               I1dff7459553fccefc94a6020cc248a49  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9a9a3b834bb25862cbe40375e20c2163  <=  0;
               I9acec7aa4b420b7c820028b669a8bfb4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1152ba49a018ec527bb8091c0cebd737  <=  0;
               I714b7d8b39c4135183b605dd97ff15d6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1cf3b72b3aa02961788688172c1ad2b2  <=  0;
               Ie5856c36d9a310f890ecc5220590fc3e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I09293a7f47ffb53331aad25a876d2562  <=  0;
               I062b1d8d3b6fe6d8e158ede1f0af9eed  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic00d9c70df8f473695a4aa76827ef690  <=  0;
               I0fbd5b5eef6da9adaf918390f6bdbc27  <= {(MAX_SUM_WDTH_L){1'b0}};
               I36132477ed96c4731e46d24e9ca1e9e8  <=  0;
               I73fb14b30841cf67e96ba329fdfa3e35  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2cb80c174e5ddbbaca6eabbfa7c669c7  <=  0;
               I6d6cfca51988c5ac32471fe8f4399bbc  <= {(MAX_SUM_WDTH_L){1'b0}};
               I359e17e055d03931cac7b41c77be575b  <=  0;
               Id7940e4951c96c3de9f45119043fbffd  <= {(MAX_SUM_WDTH_L){1'b0}};
               If466ac9d4d278b49b4aa91650b30ec2e  <=  0;
               Iea71361c5f846419eaa18ae4b9463ee8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I17d171b83e60410ce78a7e4fa9d17001  <=  0;
               Ib67ac5fdd6e068ee799965b51aa893ba  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id79a4b98545d81fef573054b93ae80d4  <=  0;
               I0bd84509dde112f3657bd5a12a8df72c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4e8f5e83e32143008d70a8edf17e2ff5  <=  0;
               I2caf86026460a024f752fa71b44f743f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I57cf1069290a2a5f30b75eb592752b88  <=  0;
               Id81d9c9ffa81c2653dea2e872ab2f71c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7447d4584dccf4dac9f0d359748ae327  <=  0;
               I0b4d1a08307d452870c3e762bd038568  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic4571481454a10eb7f8c0b58f9d35178  <=  0;
               Id75cc40233cc8648e21a750d882d5ed4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I00810b2849a3d3097e028efac18c0a06  <=  0;
               I3ea9815ba887e373a0a477654f136856  <= {(MAX_SUM_WDTH_L){1'b0}};
               I19be1cf97631f5bd782d8358fb55954b  <=  0;
               I8b26e270c3ca5563da39e7092ef830dc  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id7fe36cc9d5c1d7cc54ee1040e6578de  <=  0;
               Ib03f94d7e5ff830d5063cd514e7f7998  <= {(MAX_SUM_WDTH_L){1'b0}};
               If6984aadfa0583c3281a04ba48f3d765  <=  0;
               I00b05bb0b225b27562d6629725ac2126  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia7750161c32ac0507e1ff6a8fe896148  <=  0;
               I1f273682cac5644f1fcc30ffa20f8cd8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I97d6084735a682ba654fc70a9e07f27d  <=  0;
               I483725645504999df82a4d0660873c1d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3e9d85c0ca08314fe2da0fa6977942b7  <=  0;
               I689dc18b56442b8db01bd7ca4c44d615  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id28d0dd03217797390811bdd3564191b  <=  0;
               I805d665f394ff24f230bebfa6d252122  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0eb20560e7e211b67cfa8ca9e056c1da  <=  0;
               Icfba3f165f1cdf2e6070239100e9ac3d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id089d9523253f91c670099157325af05  <=  0;
               I93c51f71db0e3df7f6e2978fd93fbb54  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4db3f0e5ff2cc72e499ab5f1b9fd1d14  <=  0;
               Ib7410e44d23eea21613074695b64bd2b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I082972cc68873126a258e9db29e524f9  <=  0;
               I93cc273684a376d76a2e3468b3dc8bd7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3ba1cbc9ff352842d6d687b2218b6c0f  <=  0;
               Id133dc3fa65840136b1157fe97a1e962  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id8fbc7f9a403b07efd27c20d6d78e661  <=  0;
               Ib792104b6cf946d632f7591f2cd5e104  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0628944b437e239b25736381fa59901d  <=  0;
               Ia44bcc8308360d3e6fa351bc108df3fa  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icf6bf0aab709fb68c18e26f9fe7503b7  <=  0;
               Ib29a26c41a3ba089efd30c3256106a7c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I15947ee18296366e3e13cc9727ad2ebb  <=  0;
               I8999f385aaf15b67e4c12e56c7dba7cc  <= {(MAX_SUM_WDTH_L){1'b0}};
               I23b16e4f6f2fab529ae42009d38cee85  <=  0;
               I202980f6263e3b312c38061224992740  <= {(MAX_SUM_WDTH_L){1'b0}};
               I51e128a639866ca032029880ae59e874  <=  0;
               I1fd9ed3763ff0ce0a671360f83bc3613  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib14c75f869e8f09519517f3fcbdfaa7b  <=  0;
               I4b58194aa6a5b5c825f14bb926a0ae9f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9ceea65912b0a100eaa0afb42e84e5bd  <=  0;
               I706daad77f6a6eddf5576c238fa4714d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id93be78cd06b38e1d7ec35ee66f878c3  <=  0;
               Ibceceead1cdcf8805e9a9f93b3b783ca  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia61e18c0042f8ec7abb670e7f0648b45  <=  0;
               Ia5956c899daaaa0b2b0c16f524feaf98  <= {(MAX_SUM_WDTH_L){1'b0}};
               I117b1ef192f2b24c6764c2d96864cc5f  <=  0;
               I7f353333180ccbf6a271c9745430b199  <= {(MAX_SUM_WDTH_L){1'b0}};
               If5224b5f45318dac2a64dcc72c6afad1  <=  0;
               I958f0106e3ffe429d0450f4b6e9ada3d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I41710bb2545ba34f65e6d9a24086185b  <=  0;
               Idf02454b4aacb6ff03288bb19a4771b1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I15a9f9397a5d23e6885ac887723a8a19  <=  0;
               I42f39cecfe5c3d77b3fffb624cdb2c0b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I46f40fec14e2e6d5060c97f0a0d86696  <=  0;
               Id7b0871cafd2630ba4dfc3e058613908  <= {(MAX_SUM_WDTH_L){1'b0}};
               I06e512c9097f76687d65c87f99c74764  <=  0;
               I18c1c4d71799c5da8172f6cc63d2d37f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I17759c97920685cd28c898441838531b  <=  0;
               I7d53f3ce487b0a2446d5205868c29175  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie7da1180f2c4eb8153421db4c6317a50  <=  0;
               I37fb9120bfe27a0e7449583dda735479  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie6fe42c4fa7e64067960cab4edee83d5  <=  0;
               Ie7e15e6743a750cbf1b272da694b47dd  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic064e5425fd7a36be5860a40bc765994  <=  0;
               I66a1e62b25bce18e36d78c382b40b1df  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifc8326ba561071589aec67a7de4276fb  <=  0;
               I9b81ec12daf51cb61f7dc0b9ad01cc1d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibc55f69c8c895e9fad768b4b1a4a7a20  <=  0;
               I9d76cb6c99a69086774f7fd471dadf53  <= {(MAX_SUM_WDTH_L){1'b0}};
               I50b89d077d160ee7d56376ae0abd9c6a  <=  0;
               I4c59798356c8e05f8b2cdb4e202fc4bb  <= {(MAX_SUM_WDTH_L){1'b0}};
               I59a2c5b8dc1924b8503c24efa60c0c4a  <=  0;
               I395b43b11730131a5f4331b2ce82717d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I57a7c62f6cdf0fa0bd65df83a4904e36  <=  0;
               Ib3f07793c2e2cf7b6ac988be01a55829  <= {(MAX_SUM_WDTH_L){1'b0}};
               I733e71d48b2ae728b9d7b6a86261a156  <=  0;
               I05ad19dc723fe482f93cb524c8c86cf6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I20386e26c247b478dd7f2c89e73a1016  <=  0;
               I1db8d47c1852578aa6325919279419b1  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iaa6dcd47c9356b0b3b93d83f87c7fa05  <=  0;
               I98ec1bdbb599febfcdc06dbf807ab781  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8913043709d09e66411b5e70b0e3c969  <=  0;
               I86f73b27c90bbd800b521fb8953d5506  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifdcd9ff3c567f73e0366261dd09dee05  <=  0;
               Id117870de7302febd51da982ab8b524e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I95af25eeba42e7fb3dc0dff9b702f61e  <=  0;
               I6cff1d82f4c1bf7789e39b964dd9e6fe  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idf7fd041b837ee19551784f305c4efa1  <=  0;
               I5d9786c9b4566669e7981654c3c10da7  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ida9601d0e04fcfa1e448b681c4aa6bdc  <=  0;
               I83dd9071e7e35d7165d556a67d2d1658  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibf6735fa3cd381ba501ab67979729a08  <=  0;
               Id62c5db9d4a4e5eb91ca4b6876d36a9d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic78e2d18e11538916e6726418f181e48  <=  0;
               Ibeb5414f37bbb8176c1a9ac51957dba0  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4b62c23b8d6b70c44af359b951424df1  <=  0;
               If40561e9d6ab97e7dc2c6eca6d0725d8  <= {(MAX_SUM_WDTH_L){1'b0}};
               If6467cc6d4b393b76586f5b65ace1435  <=  0;
               I630618151200231dda94b3fb59a24829  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1e79f24aac8988678a3ac91e9dfa493c  <=  0;
               I45948c2ccae2bd2c2fcfe9c75787e2b4  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie3e87c23a6fbd77afb7a98ba764d937c  <=  0;
               I73048e349b470dbb16b2b3e69aebcb3f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6406707a5545040df609c67f677e983d  <=  0;
               Ic3a706eeb522f64147d4946983a9fcb4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6aacacd072438b5172d5bd0be77c9ff8  <=  0;
               Id8934e8818877e81d701105823366043  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifea8a5d86f6681180539911cf637e785  <=  0;
               Id5fd5653bfa014fa0e956ef4b1d83291  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8101cabc2e8401f77a50d561a53b385f  <=  0;
               I41821f6b5a613fde6539e41a6a0c7b65  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9574b260963de729540209c0138de41c  <=  0;
               Ie8d437ed136f7f5971638d1f62ffdf15  <= {(MAX_SUM_WDTH_L){1'b0}};
               I791728546a36e98c0d5c4eb1063082b3  <=  0;
               Iaf46eedc430b55905d73486ac0752c8f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I338183bc2bdb39e2a3820a768d78ebdc  <=  0;
               I32671ef3896bd0b586f13c092dd04b9e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4197bb0d6d0465aeb6fd7f0a8189a368  <=  0;
               Ie8bfdf207d647c9f161bdf265a8472b4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8f0d7e1f97b611f6c4a231338aaba68e  <=  0;
               Id44fe933294cafff88d133a0ddc1a832  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie50a86c3b69d3884c72948133083e099  <=  0;
               I20c1f8e56a14db0665160ecbb277fb1a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2cf91b227a82701d912cf9e9e1040ddc  <=  0;
               I7627f96e870f6a3e8abd7ac494bc178c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0f50e2edf3586292da17ce7214d37038  <=  0;
               Ia2d3997dce108f85ed64e88780e99efa  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id7666dd5135e45a1e42f13ffbb8558ed  <=  0;
               I6a25dc88186816258f1237123ee4968f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3dbcf0199e35f410c38ab3d9e2cac2ef  <=  0;
               Ia9d61848b5384a8cc63321201174f3d3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I06c6db30fc7e63facd144d0166702e6a  <=  0;
               I53ed79856aae53b180f28b47822e89b6  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id20d5070afe5748b50833f0593777c49  <=  0;
               I76503bcb779e039edc9acfc03a2d1ee6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3d041f7cf6c679d8d9677445eac96640  <=  0;
               I18ae85d6725cf0ab3b69bedeef651425  <= {(MAX_SUM_WDTH_L){1'b0}};
               I51d27603f0a87b78857b8e064182d925  <=  0;
               Iaa3bbfc6704e70a55b8e1083c326820f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9b6d48e71d050b9b0b5c5e7407288103  <=  0;
               I8c1c3ee4b57d56ab362672dfeb4e0ae9  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id05706fe9e0fc4776e0446aacd4c118d  <=  0;
               Ic8e0765b1cf95f2578a7ec656d027f6e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2ec61e0e1b707857ca39f532bf970e03  <=  0;
               I39eaefaae486119c8741c5e9b7f85bd3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibd1b4a1010823cc9e4a78a0fcefd7d01  <=  0;
               I6ac8d8000e434fcca222525ac00f9849  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6da2861072f65e35d46d224b982eda7a  <=  0;
               I114cfd3fe8f5db92b879e0dce592af3b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I860c7e185d38d907c4ed20a64d238dd6  <=  0;
               I8db1c7f6b5c7c04f71e7fcc18f7b9941  <= {(MAX_SUM_WDTH_L){1'b0}};
               I76e06fe466c43e4aef0ef860f0274fa8  <=  0;
               I89e516738a408ccbd495e4f5aeeb38a6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3c00d8a5dd8c99ee527ad4180e469ab7  <=  0;
               I0c02b9318bc4f50969f8d486e587a627  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iba2018bad14888e510fc7f4a4e040ed5  <=  0;
               I79224b17e2d1f87175f3118287351e0e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2e3d469ef08219887c92189ad3759da9  <=  0;
               I41ee2f859df1db26618ab9c2c0a57be5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I74628364cf049f0e6de34bd1f9853985  <=  0;
               I15a667ea371ed0fd464f42fb9ef61766  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifec818042c24c8eb96832c782f09ab04  <=  0;
               I25c2d3dd7fedd28f0be0e3d8dccddff8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0aa52a892c8969087bf3f158aae7078a  <=  0;
               If22b31d70158d864ca6b0201ffc2b7c3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I31b799a3279d7d66b53f4be544498602  <=  0;
               I7950b8505327240095538f60d81834d1  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie8e004bf6e301a4ed9d9dcca91b2dc85  <=  0;
               Ib75297152c09323c7a6f674c93edc01f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9995a84609ef3fe477c73f136515ffe9  <=  0;
               Ie813deeac800a6b251209a1c8e2adb12  <= {(MAX_SUM_WDTH_L){1'b0}};
               I54e519ab156fdf2054472d4684de064a  <=  0;
               Iada283b3152a5316b6c7077292ac0a29  <= {(MAX_SUM_WDTH_L){1'b0}};
               I527950bde49a5c46e818225e41bec4f9  <=  0;
               Ic14e12a907c5d6b7ad2615905a64886d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ieb876e18857117935ca3aecb6a525b1f  <=  0;
               Ife78b0889c9c7129a3000cca66ae4aa2  <= {(MAX_SUM_WDTH_L){1'b0}};
               If22f8fa601e72589b3a5779f23ca7454  <=  0;
               Id926d49513e089a52b17978a9ab84372  <= {(MAX_SUM_WDTH_L){1'b0}};
               If222f8f81e40570854a512fe828f9ea9  <=  0;
               I4dfbf2a2c01ce39fea9b756f9b106fc2  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6bea78584853c37d7c4993a45668542a  <=  0;
               Iad7cce628396ce9ffac3ba9dde7ac494  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id7cd91008312189123519e44cfb2e141  <=  0;
               Ib71f9f92515c200bd16591c656d69ee7  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id3c95ac844fe01a85e6251683bb3f9cb  <=  0;
               I8e39b301e04135b8ab88d54e7c1e22f7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I49b96dfb05812ec7b0632bc722d417df  <=  0;
               Idadba73fb37b81563818e82af3d89a58  <= {(MAX_SUM_WDTH_L){1'b0}};
               I89b8ac7adba1c7fe4f04e408857c92bc  <=  0;
               Ic19accaf42ef2b61fb52ab3621622ef2  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic1a67160ca63763ce6b850bed5371d32  <=  0;
               I94f508ac67f07b73b3ff1d5aa5955eea  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iaa1ed0cec8df6dec4fb0ef9c57c98d19  <=  0;
               Ieb8588293562c9c25897044b9e5ed6a4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I76465e13c5a9ac236635e663e543487c  <=  0;
               I671d71d9ca760cc759b96bbacd361f90  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iff18998e317563a12db412950315b397  <=  0;
               I3f793de7fcfd045af3970e4ec219128b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I279642da9295f410b7482eaedfbcde75  <=  0;
               Id49f950b3679093b10f8b64ae89c5558  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iecceba6850d58cd1500bb5129abc8035  <=  0;
               Ib70c7567e552969a2757c1f48a2468ef  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6ede97dfb1484ba6fe621c7034e22c0b  <=  0;
               I6dbd0c3ac9f2b3887d87e316b8b40b55  <= {(MAX_SUM_WDTH_L){1'b0}};
               I57bf6d033eb5643e96bcdefcfeb76a46  <=  0;
               I8c309d7fe6aaa8c996e39b8f3dfafef6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5ba33277f07eadbc27835afa96bdc535  <=  0;
               Iefdfd7b1924f8b6049b02576f9948027  <= {(MAX_SUM_WDTH_L){1'b0}};
               I256096a960771679c9a7a391448aa711  <=  0;
               I2c14ee79492962576e12ff1698ac0fe1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I220f38bf301ec4abcd1e07727fc5bae8  <=  0;
               I56e90395afb09c7d775111d19856da1d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id6cabb7608d470ad7dec1951618efa8c  <=  0;
               I90f0c524f6b98c28d18db952ac40c83e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I30ac677d67ab06a6f5759da2717ef6e2  <=  0;
               Id50649fc4e9de24fdd9f06499a733b87  <= {(MAX_SUM_WDTH_L){1'b0}};
               If0881734b6b8bb6e3e22823408203887  <=  0;
               Ifc988e99b4c4c1ba2d5cf3a76695900d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I29502a6df7b40a59cb84f6c1a0d30fbe  <=  0;
               I53c579c64f0d911fe3fbc43dc3e981de  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ied5d76051c9302e2594e5f1c34dbe8a9  <=  0;
               Id729d27d6424495fdb4deb2ffc038f01  <= {(MAX_SUM_WDTH_L){1'b0}};
               If6c801f61074108c3342f1c3d0b4a39d  <=  0;
               I8816c4edb8c7f5fd6e7a3c81013116ce  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3f15fe479ccd6715b63db728ffa8b49f  <=  0;
               I88ba486c5bca54f6c120a654b81e0a90  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id7e322ddf8565bb59e6377bfc7b3ab36  <=  0;
               Ie1ba6d92c19ebbc5c994d9da3881f6c9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5a325c188a650a75ab298719c0287618  <=  0;
               I023278cb7d70d4608259e10c89e97117  <= {(MAX_SUM_WDTH_L){1'b0}};
               I763f7f930d12bef17e0aa5ed0d6abf96  <=  0;
               Ib8c744194310bd59e983e392b828e9b4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0e34522d1f95f50998246232512bb60c  <=  0;
               Iaa2aba39e0454008fbeff8f9aa87a481  <= {(MAX_SUM_WDTH_L){1'b0}};
               I45b69f889fd15cce35f6812afe0f4894  <=  0;
               I61a43aad15d7a9943f74617f434af306  <= {(MAX_SUM_WDTH_L){1'b0}};
               If4db281fdcf771156956dfa30e36b29c  <=  0;
               Ibd8114af3027bd3364395e7b94484272  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib312a09daf5e5c38dcd59128256a3ebc  <=  0;
               I49167fd9caea095581855b45b1f85d49  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iaf3e2d448016a50829b4b0ea6f144b27  <=  0;
               Ic502f151ee9ee01786e216d90a29403b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iddbd5820346c3ea47bea79b2ee1ab7e5  <=  0;
               I25f89c7f7f11c7e2811913d6254dbc8c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1b024f329d24692f8d143aeeacfaf555  <=  0;
               I3f939889c013f740cc63c981d2ff85b2  <= {(MAX_SUM_WDTH_L){1'b0}};
               I83f200ddde413f07bd296b8602aacdc7  <=  0;
               Ib0d2fc4f353a82d37bec9aa19a80475e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib4cec30021700f9f02847c2f1e0fc425  <=  0;
               I2f19b77e5bb1b22b3cf5b1ace31ee6af  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3cddf5a4ce875cb4e0c2fce7e36e5200  <=  0;
               I283f82fd4a9700daca6ff1d16f747a09  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9c5d93dc3faea27b0f38898609b41545  <=  0;
               I8dc5483fb01a06ad8650e5fd4df30f49  <= {(MAX_SUM_WDTH_L){1'b0}};
               I426a2f3c939a72ecff6a6314a19d52cb  <=  0;
               I7e3f6b4bff19a0644c12fa4ef3667d84  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5919e3d3ea27d29a8093c52a6645959e  <=  0;
               Idf2371d30bec7ad5dea346a4a48a6e75  <= {(MAX_SUM_WDTH_L){1'b0}};
               I68c4ab26cc7c41ea3f9b8afec502bc42  <=  0;
               Ifd5a3069363cfc42e5a436856eeee708  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id4ea7f8c016571cc5a0af8327e2f95b9  <=  0;
               I1a4e12577ac5e87d40bdcb54fe55818b  <= {(MAX_SUM_WDTH_L){1'b0}};
               If6b109772fc17d898d70f75f538a0fdf  <=  0;
               I1f1b6c20910c4f14999da6c9fdb4c349  <= {(MAX_SUM_WDTH_L){1'b0}};
               I930235d80caaa415247c7fb380b3a134  <=  0;
               I1b0a200eea98f075f059d2a26b00f833  <= {(MAX_SUM_WDTH_L){1'b0}};
               I324eeb4bf0e552118536fbd641189af1  <=  0;
               Ie0dded072843efc1613cfe7136af37da  <= {(MAX_SUM_WDTH_L){1'b0}};
               I839160e07222b1f9f293efe22d68c168  <=  0;
               Ia6d6a867ebe63a8926d9affa4c15e376  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5244962685ce36dd805a7dc774c05d31  <=  0;
               Iddfc447b0c96056ae6e6434799ea00e9  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib92300e3d61e8a2bcaf0b2f40d4cb18f  <=  0;
               I36d03daaaaa37229d462f4bf5e521f73  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id76c8bf8796c329353836a52e1dd74c3  <=  0;
               I91e49319831eeee5dc75eac77ed8f8a3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibb163802022194494881194dc6b49c2d  <=  0;
               I4e9f03752b041491ae2bc40fbd2b8d43  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iedb3b8bfd024408f08a2b377956239af  <=  0;
               I9a71e50dac7ad707a4b0946ebc1fe6d4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6cfe7ce048413c7c959a0eefe967885b  <=  0;
               I8220d15825d6bac07d773ff0db2f9795  <= {(MAX_SUM_WDTH_L){1'b0}};
               I664a362c93dd438aec485063a6f0c7de  <=  0;
               I6b2dc98acc78a1151dd6670ed981d839  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9252e19b54173ae2a9d0815dfc46eec2  <=  0;
               Ie371be4323965591a5786063ba028ce1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2ea93b2142eee9f44c8e7bf892bf02ab  <=  0;
               Ic4985251ed9f9120d2232ec96949831b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6772834728b2e641c6e3c14cda255ad6  <=  0;
               I6015d64c067415fe216d90a5be409e33  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id6a64c33b3beb88abcadc06af18e1858  <=  0;
               If6f304fe091216273270713c6b6e8a6d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib89f2aee80d36f4e473d1a1046e836dd  <=  0;
               I779ee6daefe3c5c96548dc5e0ba83bd3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I78aeec1644701502f6f71c64341274ab  <=  0;
               Ieef21b505cc215387f8930888062b767  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9a09fda6e73783a7c9a4582fec8121b4  <=  0;
               Icbabacaecbbac74901402e5e5874328b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9db6919efaef0952b84eaf8e71f77777  <=  0;
               I6ec13a161f7f1a0f57e9ba4998474954  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5a4646a8adf0ed43a905fd4ee84d85bd  <=  0;
               I71f9823e92c51be2e9a050d01e63902d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1e3444ee88dc52881397d266f469b45c  <=  0;
               Ia0037030d79400734732f061fd81edf6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3c42e969e5e4b99f1f2eaa01419d4ed9  <=  0;
               Id796584e3e7af67536a27f7299b71916  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9210d06734058f76e7a5a470dbe6e74b  <=  0;
               Iec938bc1bbad930fade05d74c10989a3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2b35c8fa7c947b3e7691cdcab0c5a7a7  <=  0;
               I2a7a7c5eabd1623c1c3d4bd93bf18617  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id58d1af007bb5858499af71a43e6574f  <=  0;
               I71cfc7fd85636c5554b9fe9f9ba8e3aa  <= {(MAX_SUM_WDTH_L){1'b0}};
               I12e92aa9c9ca2135f7ba879d82ad615b  <=  0;
               I4c8ae97548bc3dbf3e3621f80c3e0835  <= {(MAX_SUM_WDTH_L){1'b0}};
               If32ea54eb47d27e35a81aa4b9e1f7713  <=  0;
               Iaa93c760705c984a0eea90d41a6c049b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib1ddab09d1a726176414e4a877b66e3f  <=  0;
               I2acc73851f8a803e69c0f1865e00f46e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id3838f634ce2d90a19622185391ba868  <=  0;
               I928333e9cc75d49fa6f7094e49631123  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia3f429c43f23f4f057abed98cfa94748  <=  0;
               Idf02dd4b7e8a6958913e6180fec1feee  <= {(MAX_SUM_WDTH_L){1'b0}};
               I62b423a6061215d16871bfdf9a9cdbd2  <=  0;
               Ib30cc7931858974728d92eb68890449f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I17f82f6daa8a92f1da5a1952a558ad7e  <=  0;
               Ia504dbcee6e5894fed83371bf70b2d44  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie0e9f7c1d69d8930f8452d3618512877  <=  0;
               I32b4e50b8acefe1c108d777da565f4ed  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id9de214d84792861772ef396b5b9208f  <=  0;
               If9fd1d8c0c13042a6f2d258478b63925  <= {(MAX_SUM_WDTH_L){1'b0}};
               I027f018e60dda98666458cb69a6e4be2  <=  0;
               Iccb437017198e4421ab51d74aed779f0  <= {(MAX_SUM_WDTH_L){1'b0}};
               I996821515569c215f3f688d91dee8abe  <=  0;
               Id10bf2bf52a8f1be9eeafcefd6dd5dcb  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6f617bfa2700fb385d425f6b4581f594  <=  0;
               Ie590c921147b7252d2605f7712dfe437  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id5f8b6b344dc8e629f13e5d157f510cb  <=  0;
               I178ed883c28bbf3e1ab05cb95f62b343  <= {(MAX_SUM_WDTH_L){1'b0}};
               I579a5dc98f16e0c5d52fc7958586a8d5  <=  0;
               I01971a175615a422d264805252f91f3b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0f2769698735ab28df30370c3c8b56cc  <=  0;
               Ie770c4567f35b40c46ccbda059e6d3a8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9fbc79fd7be52757770dce6e04749b4f  <=  0;
               I25975702f0b9c0baf586fe471676dfea  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idfe33235c2f93ac311da89ba63e0f1c5  <=  0;
               Id2ef737d910326394b68eaa0833bfccb  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic46d706f6be34cb4133a4128567837d3  <=  0;
               I577cd1f9ad512ec10f5008165f2e4a74  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibb3c635f2e62a63c9bdb150b3cda7155  <=  0;
               I1de8f87eb39276e073f5804b1df3b67a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7bdfb2d2b7dd18fc7c0d43b708fb1e35  <=  0;
               I7f8e7928e6caeac14f787d7e0b6a47df  <= {(MAX_SUM_WDTH_L){1'b0}};
               I42a1cd616514a1c7384d07095e6b2d70  <=  0;
               Ia7048aa3f949b0b2e54ab900efe01131  <= {(MAX_SUM_WDTH_L){1'b0}};
               I19a91106f189ef43ee50edab49d297c1  <=  0;
               I1fcbb73d165eab038c745fac370fd68f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I90088e4928092e62e193039faf154240  <=  0;
               Ia822cd52015d599bc45ae7338b4e88e1  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic0fed8f997e03bcca119270589f8bf0a  <=  0;
               I56b85e2d5a7259eb50fa983b92d8b160  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3ba811abe28766d976a2afd02c22fc76  <=  0;
               I1d23632f8e8f66a30b4ef6c76aae3ece  <= {(MAX_SUM_WDTH_L){1'b0}};
               I66463d17d0fcb691e727568e4d55ae43  <=  0;
               Ib578de11f0407cfeb0dac68bd5fbf7a0  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icf73bfd92fe6265b8e7d9b2439573a96  <=  0;
               I08879fb80c58de5fb2bf547ce013c67f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7c3f7076072ee81960c8b0187648eb41  <=  0;
               I8f7c4c602b7de5d9a401d3933a7e50a8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I68ccb34c409f89f1a2872d64f85e3245  <=  0;
               I2ab4cc1ef6b743cda8765a22e28fd7a7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I069661eba4d8f68a4e5c78e99e9355e8  <=  0;
               Idc58a89f7d8ee884b198b6e4752ec58f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6cc756f9cb1020c8045872d628b771f8  <=  0;
               If9c0f4c64c7648e509077df16c14b7a1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I95494fb67de54f6055f54c7568106488  <=  0;
               I8cc434418203702ad5a21eb4f0340dc5  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibbfab9efcd61f23b09e371554c0778b0  <=  0;
               Iee9d96f800fc848f3c4b6b6901a72623  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibb2a246712268d6d8a0ad0354b8e611f  <=  0;
               I989036e56c9c7386279e83ae83ad4f7d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie9f5d2f06f60d7f436118f2c92695107  <=  0;
               Icf23ca0439c76198fe647a0b785d9503  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0ee25f335a84b7a190ccd690fccc1fce  <=  0;
               I406bddf2c4a4b6e6aedb86d72f14994f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ica83129589b16c7392387bcddd9e81e9  <=  0;
               I5331e97930599788b1df06992c5e4a5c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I91fc1c1758eb8c136744c1ef47785b49  <=  0;
               I98577e71126ac9bdbe4359101d4d48d7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2bede76feb8d499cef693a3cc0bb95f4  <=  0;
               I696f551b6f96d0f7d27eb685bd374229  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia0d9b7bd503ddeeefe9d0646c1f4e6d8  <=  0;
               I1aa256ab19406597846ff353b65224cb  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2af1f93bd1d85a66028ef0add7a69962  <=  0;
               I00f1b24291a0e8496e13fe076e377cb8  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icc568348313201d6814f92694d7db06f  <=  0;
               Ie6f40dc356120aeb6cfa7a3fb5fae8cc  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iba815b719f813a245efb2627660634ff  <=  0;
               I67e23e6286edc4e01a7ebdace62ce56d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id67d39730eb990c4b125cfa772e27e3a  <=  0;
               Id2c7c6d20146edcca65120c025e25a0a  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib09008d80ae9d6708371c0c40f157656  <=  0;
               Ida1e2d8b0e45e14c4c669c8b9d6947f5  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id61b17db82e540f939ed8a4c3b596278  <=  0;
               I1fd443d00410d0577eef9f1f26e64700  <= {(MAX_SUM_WDTH_L){1'b0}};
               I24868694c2523bb657da19c2e84ec8ef  <=  0;
               I9ea760f08ba7b84fcaad929a3669450d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9dcf88e53c655bce8190c5e85f5ca777  <=  0;
               Ia522420603dbde92a49da297554ede5e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib881ec4b6a6de42dfcb2be830ca39ac8  <=  0;
               I9be575cacaafcc13a0306545be56a04d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifd2ece02d5ffb0a50d8b151a8fa8e703  <=  0;
               Ieb9a03ad2c7c7df356477e8b4224ebd9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7da3a787760c42ef510ece8234c020a8  <=  0;
               If7f263cb2fb7fd35682d44c42639bab6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2204fa0d852e56e843393b3959f3df72  <=  0;
               I5046227e18f800785f8ddfb4a89b1bea  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iaee3ca649d20dd29363781e8dcae17c0  <=  0;
               I73feb8438775bf3faffed6895b6a4638  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id8bb7c6409e383793af592892caf23e4  <=  0;
               I6a423d4e11a97d84120a475db8fabca1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I96c6b861bfaad7c411db93f1318d6b87  <=  0;
               I2098616787bd728bc4af6be5ee094bae  <= {(MAX_SUM_WDTH_L){1'b0}};
               I76eb400ed4d1502f7f1864d9556948ad  <=  0;
               Id9ef21a12edf48e574256ea34fcde992  <= {(MAX_SUM_WDTH_L){1'b0}};
               I02155a5c26345ff00d18cec6e2f01592  <=  0;
               I31ab57596896201ff52990b0641b9511  <= {(MAX_SUM_WDTH_L){1'b0}};
               I91e6dcd9fa2efd055125878ab38de3fd  <=  0;
               Ib3dd33a163b0c8153edb4fcc90a453f2  <= {(MAX_SUM_WDTH_L){1'b0}};
               If561e078b234a0be8c0b8ade8f5ec0f1  <=  0;
               I28496a34b2ee033767fd64f631426b23  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0ef01533d6494ce8f092d54c5fb0865e  <=  0;
               I0a4ef7fac369df46d1a4b094d7687645  <= {(MAX_SUM_WDTH_L){1'b0}};
               I782b73148fd7ed7f9d734baf42b8b5d0  <=  0;
               Ie7944f3e2adfac325808f8711c0eedcd  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2099d6f614a5f7432f6331b1bf56c31c  <=  0;
               I58cecb5376f675339028440f0671b0b7  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia8c9228b5d23c91ac06450ab1296dc65  <=  0;
               I62f85c1602819e586d9656ba42d263c3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4b76ea8b5d4ed8ccd8ec532889dd6d4b  <=  0;
               I79585885950084095d2ce4a31aa73e4c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifff6d20dcf891c78ad12a304ca757c95  <=  0;
               Ic3af09106eada35f1d786ed60e314ea5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0dbefebca7ff055a6e9dce2a2c37bd69  <=  0;
               I81e374d671edb31d060875cdfdcd61c7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8aadd755861e90ac12047f259091ad85  <=  0;
               I1e22ea5ecaf87499b7106246a824a547  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia7d21a17d62e7bfb00b83b244201e941  <=  0;
               I0e46eb0f32c91384b07c7b1ba84caf98  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6c63fab8059cc3f0c02b0dff5a8cacf9  <=  0;
               I562b5f77aedd91f0cb3df00387c7956a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8744fea2c7de33b5308dc9a2828647d4  <=  0;
               Id819e47f502c18dca8d1e804d346c1ea  <= {(MAX_SUM_WDTH_L){1'b0}};
               I04c99b4d0c54b23a72b698753510a4f3  <=  0;
               Ie0586f4b015fd32777d24c2d9856b27f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5de86a27849e73b21e4c40e9e8515033  <=  0;
               Ic28248b41552d2537d0478c23e33e0f3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I185257f76b2886cd845e50a01ef5b05b  <=  0;
               I3463cbe0d16b14aa670fda6a0d34e255  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1a2c7b5505f4124f945a28565eed6013  <=  0;
               I0aac7a09d9253385d34e87bfbb216a79  <= {(MAX_SUM_WDTH_L){1'b0}};
               I771d417f6226b04ef016d0943bbc4584  <=  0;
               I305967a657db8531d1ae309fa3e3b98f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Icb0a73f2dd46e2195d5efd34fba3a985  <=  0;
               I0524108ee49eec5fa7861bed35e4ea3c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia992f7eacefc028526ab4f105e244e02  <=  0;
               Iced1e0b874918a1c66e28752e340a51b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I85454620b6568bb7fde468a2e9a5fb42  <=  0;
               I670e910f74fafccaa9f1a8279fd6ebb6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I87557ef641a7b209d4d210498bb15271  <=  0;
               I02fe6b32b2405fb94afd5d7abbaf0195  <= {(MAX_SUM_WDTH_L){1'b0}};
               I28d1125b647b953f2a19ecd6edd8e450  <=  0;
               I5f5304e4b132f816c87248d3ca954164  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4a8aa3010248f0bdd3e31822bf2fe0a1  <=  0;
               I0ecebe47e1a9ede33c3995945a6ee760  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie1966fd5b564dd6eccfc458e9c6aca2a  <=  0;
               If425109071b5310e097d2174625b6383  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8ad51753f106d0a30cc79bd08e799348  <=  0;
               Ic0f324c7ba05a7cfae9d70b62e30f94b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1c3bf915a6b62d22d04b8c8d92a72a73  <=  0;
               I35631cbe926290974c90ddeb9b07f231  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie557629e9d52e5fa7435b4fb19e5276f  <=  0;
               Iceae425f37f3b1194a2ef5cd46d1b6eb  <= {(MAX_SUM_WDTH_L){1'b0}};
               I38fc977bb1d52cbc5e02a6733f6a8190  <=  0;
               I4faa2187d970078870078c3eff180b4a  <= {(MAX_SUM_WDTH_L){1'b0}};
               If84914aaabb020baad2b222f27c9ad38  <=  0;
               Iec2860f518edf688a9b1b2736ae00835  <= {(MAX_SUM_WDTH_L){1'b0}};
               I54c457a658721fa7de175432b340532e  <=  0;
               I20e7b48527e4456874d59e50c723c6a5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9036f6cf74a2aecd827c7239da13db70  <=  0;
               Idd60af0dbb02680e11c1b1734f23b895  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8825e2665dcee58925a5106a9cbce9ca  <=  0;
               I79cfbb5d5e920bc8cece60565ee0c5c2  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic3311c2f88a7ae151999b2de86d82dfc  <=  0;
               Id765a3f659dcdf01cfe23cafdf066f92  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3ef7eddb92284b28f97feea52f489aff  <=  0;
               If370aaa56b4ba3eee873c99a86577c3d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I68728d0cbb3a84370006277186a0829d  <=  0;
               I4508376202467dc1bebc69757bd5f95a  <= {(MAX_SUM_WDTH_L){1'b0}};
               If5bdbdfa73406a6a9d426920f51fbc73  <=  0;
               Ibf115f80ad72df8599073c05ac58e028  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibd3179c01665a17f9c232196648de8d5  <=  0;
               I27960a9d3923d053d466955c660a91ca  <= {(MAX_SUM_WDTH_L){1'b0}};
               I42c2c03a158ed79ea91ea6b9f9a6f243  <=  0;
               I7c52711e3b71823dd47861341d22adc3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iec064c18b262b95bd6412b1e50e4b5ef  <=  0;
               I547ea6a130740e4b0bb85f6c9d3a6549  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0470f0fd133851c1241c654abc19992a  <=  0;
               I0ec19c18ef7da4793427a00a652a9a35  <= {(MAX_SUM_WDTH_L){1'b0}};
               I550661edfa7a7b440d43c0840aeed8fe  <=  0;
               I640d147f241267ccc89f9ab132d724f8  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2f01145e1b41f2f7103c5247bb548a6b  <=  0;
               I3507152877484394769c12879ce0aed0  <= {(MAX_SUM_WDTH_L){1'b0}};
               I34d143e9a6f936b83863a5ebdf8afc43  <=  0;
               I382f86490f568ead2dcf51e8bc6989f8  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id2f831bc219ca3f43c5c4d69f6724e64  <=  0;
               I953178c54a672474dda2f48c70ec21a7  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib708fd61ab7016190a2a7156439201cf  <=  0;
               I13b43982093e885ae7bb04a2b61e4eaa  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6a2e574a2d27e40faff379b6c26ae51b  <=  0;
               I3d7491ac28a4adafbc138d17f08c9111  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4be2286baca2745e981a0d153c0f5c42  <=  0;
               I3e0ca15752add87cc01981e7d89d53f2  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib9643265dc8c283d7b0c7afdb19101fd  <=  0;
               Id1b152deea3ee894ed5a4c6ff10a6fda  <= {(MAX_SUM_WDTH_L){1'b0}};
               I78d7637bbd13c620434d3619e615114c  <=  0;
               I7df9cc0e3ad69985fe9a3c8f2dec1de3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I358ee555d9955cdee436375ff898f4d6  <=  0;
               I52910c0c2d26095c965d32b85e850d92  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic3961c918c81b14d964e96892b95f00b  <=  0;
               I93fd4b4f7d01ec59834f3054fc2eddfd  <= {(MAX_SUM_WDTH_L){1'b0}};
               I580e98d4bec3eeeb1642baa425a96099  <=  0;
               I481b6feb1f1ced501a157b06a4782e05  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4cec0a54301908b3f58166a9b0ef1eb5  <=  0;
               Ie99b8f3190ee307e743255156b7f7f90  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib7f7c88d83d207bac3daba4658342879  <=  0;
               Iac858597facbc0025a4760eac49531fe  <= {(MAX_SUM_WDTH_L){1'b0}};
               I371401ca0c589a1b8fa816beed36ab0c  <=  0;
               I18c2833554a5b358578e7b6901c91c0c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I81f561f223b916600ebc572c05dedde5  <=  0;
               I0cc6945a47b3ffadd1e52e3f71c9728d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7ee36d73f8c69e5e017f4616094d992f  <=  0;
               If2807866c5d481cd31c69b67ec537a4f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I706d7d2238c5882491d479df0cc40c3e  <=  0;
               Ib24d495a86e15d9c8b2c8d360445e511  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie28bec241cb36d75c1f2ad846dc5c7d6  <=  0;
               Iad2cdac80bc26a0c50335c6467921c94  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9fe8aa4f9f74c1f004e5bb536e902ea2  <=  0;
               I18c93f107d0520171864b789ae9707b9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I444003b27464f275311d07ae7d4fe016  <=  0;
               Ifd40aae90a89d2420e43fe4ee533a1a2  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibbe636e1e98bbd4cd97dca56d769d269  <=  0;
               If46a176f32240b03ae959e9ad889fc2c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib195ccbfb4411bd3aaece336a5aed65b  <=  0;
               I5e7b386298be05835cd24554966cdedc  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ieafb75c62922cdb3acd95a9614a86efc  <=  0;
               I5258d2bd4ae07dcfe7e022b046800856  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5d7018ab259e054ecb48a238f3c03208  <=  0;
               I14da6601ba08fd3e9a2bcdd20bb43536  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iedabb09ffcf910c4dbed2f142dc96df0  <=  0;
               I76bbfed1a115c2f503531682cd171185  <= {(MAX_SUM_WDTH_L){1'b0}};
               I07b84cae4f002659d68f5c1746416e70  <=  0;
               I64f37f25618c6bf5b35e863e3be05a3e  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iba31516a82e9d2a5ad1a1c89dfb6af70  <=  0;
               Iba3b847497a7572624a3a1f172b47d3e  <= {(MAX_SUM_WDTH_L){1'b0}};
               If5c42feaf3d586e1f2285b0f3e3a2d39  <=  0;
               Ic9885fd472d244d4810bc9ff0971dc65  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3f15f6722f339c32bf1dfa41b5b24648  <=  0;
               I5753bb74c9d925b91c0173bcc320af36  <= {(MAX_SUM_WDTH_L){1'b0}};
               I74d5d4a25b6ceba088652dbad9c35bae  <=  0;
               I66cf73ce0a93f90287df52adb628716d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1e3e7019425109b26d4ebc7522074e33  <=  0;
               I84a477263ea86f2014d28e9ec928fa1b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4f0d4baa740b2f9bea59f4653cc9e8fc  <=  0;
               Idda9e2f9a5e24406700b04e6035dafc7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2df393a2d764f120433f310797abb2c3  <=  0;
               I694ec5f3a1e7cfc02c1af8369064967c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib9a2e4c37430ad33531f318a313d4646  <=  0;
               Id0c6285ee3789c104e483a5626b5827d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ide344589b18aa0332a7114424956b65b  <=  0;
               If9bc7b1498733ed921b51cb613c2cf53  <= {(MAX_SUM_WDTH_L){1'b0}};
               I789b8e58762f722bc0e86e17c2655965  <=  0;
               Ieeda4b6b301d662ab9be9f6b979bb1f1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I243898aa7700f57974ea2834df469f48  <=  0;
               Icad98c93196218a7dbd25af042b4a32d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic65d6b89fc082438b9956504f30a5483  <=  0;
               I408e198b0eeade8b94c27ab7e04a8776  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibdcf7926e0b7412e4a56d2ae15a4e892  <=  0;
               I24b90526a93dc177a5d23b61d20f8797  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie552917ecc454608adca6dbc4d9153ad  <=  0;
               I4da324410e88d8c9738949c287e7bff9  <= {(MAX_SUM_WDTH_L){1'b0}};
               If3b234f8485412e76e5cc497b7c3a6f7  <=  0;
               Ie24b89ee61bddac2f2bbf1b8b5dd437f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I67c58e4de1a3413b77529f5374201308  <=  0;
               I27b99df87eefd6fcd484ec321bb73dc7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9ad9a905418216c83643eae11965f330  <=  0;
               Iaac7f8ca30f4e74e1ae5016a222673d7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2f3232289260297dfb0cb36e42e459be  <=  0;
               Id3076c8e12f28723096148d8cf91a13d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I58525519bd3b6773ec9ebabdf2764f69  <=  0;
               Ib2e36c2d0a51f5b953b9f368f11bb295  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0e369759d6a2e5df5cd4fe6765ef8436  <=  0;
               I9ef5138c78fee50aeb2568def8bc62a0  <= {(MAX_SUM_WDTH_L){1'b0}};
               If155fcdeb6ebdce7305bf57a5e8fc426  <=  0;
               Ic1cac944a0ed80e5b6e3821e8451045d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I53e38457ad9a8a8244c9a2dd06034f60  <=  0;
               I915f18e8333d52f6ec4162fe35317d17  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0cdf5ba9765cb28f2718129218794ec3  <=  0;
               Idbcf9e41a431a42028cc99d6be0c46da  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic8e633425dff5441ceaa669bdd924077  <=  0;
               Ic46dd35355bcd4470886fbd416b3c75c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie7efb37f21bcddfe6cb7969533bbaca7  <=  0;
               I0765c8beae32257c6c37dabd94cbab7c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie5a9f440574d20f6047c0ce556bc8477  <=  0;
               Ibc002286423e5ddf50b8ea25ea1b3377  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8fb0748ba8138a9188a557fcf752a055  <=  0;
               I714b85ebaccb1e11d16d53cf6bcf65b9  <= {(MAX_SUM_WDTH_L){1'b0}};
               If6261c7d9d9c1b95edf08322eac2332e  <=  0;
               I864ca16e4e93b435a94fb012d995c7e5  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib9f5522d41ddd9087096bb10ce7f5e23  <=  0;
               I227ef7de18494a9f62b2e8cf37687840  <= {(MAX_SUM_WDTH_L){1'b0}};
               I686a59acf3c8d19e90c2060b7db4be8f  <=  0;
               I535a78cff546aed9fbd1d79827d56fe6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I73ba52dc87f86c76035540575994a224  <=  0;
               I90cf52bd1332ea1b955e8c193b670218  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5947a59182e394e4b2f84b68ffd7bccc  <=  0;
               If7dc2cec6ded3b32d42281d08e871513  <= {(MAX_SUM_WDTH_L){1'b0}};
               I006c14dc1c5be7dd3c5e1e5dcce08c21  <=  0;
               Iee43875ccb00a79e67acbd3e12cb516d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iee841700cb259de93cbbfb47e828e1f4  <=  0;
               I7aaad9fdd239670e028a896695c01216  <= {(MAX_SUM_WDTH_L){1'b0}};
               I71e36dabaef7951e59fc8b08da50003d  <=  0;
               I4a992ed2550a3c5b346158ffe18c255d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I323df8d18a73cd3947512f8a2c41b323  <=  0;
               Ib2eb28843cf201e8c6f8900b7029d42d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I30604b84bad8b4bba6d340cf020ca901  <=  0;
               Ic9a5b2c8aee24c3fbc7e92b8fdaed5dc  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib436620d6352c9ad5fa1d1fb5083de7a  <=  0;
               I6996efa8115f38da03518dcb7dd42a4d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0722db2c7497d82a0ee09a109f698250  <=  0;
               I1c4bf7954b4bd5f4e9c176a3ae1fc28a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I34fe1fee7604351d37636552ecb32d8d  <=  0;
               I55d0fd8eda9c128cacdebab55a8dda5b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie9ca773a78e9592fc49a7c590a3afee1  <=  0;
               I02fcd92b426929f24b9a8c063a56c0ed  <= {(MAX_SUM_WDTH_L){1'b0}};
               I023b8de48fefb0b45bed81ada503d779  <=  0;
               I3202a0ce45afe072eb955cd6e0789cd6  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id0ac1f9bcd5fa52b3b0536f0c831d504  <=  0;
               I06c82466a2ca646abb62bcaad3d63748  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic5c3ce39ad2fd88b6a26e639e390155d  <=  0;
               I23af695cf96a03638f0c1ef719d8d530  <= {(MAX_SUM_WDTH_L){1'b0}};
               I80a34c662ed81f7d38d3055d470a1d1d  <=  0;
               Ie20b7fc4110631c1da7de4c7f38e2581  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0552127e741bcac86d4ef3994bf8830a  <=  0;
               Ic6983ef65e0de21992fa0b90ddbdce9d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idef88c7c7169dae7b6d14e0edb17f47d  <=  0;
               Ie7c2317cef621a89ad24c8b5bc79a39c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6f2e27ee85aad612520efe0e53f05aac  <=  0;
               Ic58955d8604cb1a6a20a199372d44774  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia9afdb2578f40035f59aabad30a7e156  <=  0;
               I8198473d2a666821cdf398dcf1b0fdc1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3c07ba2d2d09f45d52fbfe66bc54975f  <=  0;
               Ic60bdcbc8a55bc760e52c37aa3030001  <= {(MAX_SUM_WDTH_L){1'b0}};
               I77a2d8cfbb2e6f050545e2865b514205  <=  0;
               I987cca9a9fcbe4b617a7e524476431be  <= {(MAX_SUM_WDTH_L){1'b0}};
               If126c59dab3d743d2451279fc184182d  <=  0;
               I765c7209f3c7173362057fdb60aab732  <= {(MAX_SUM_WDTH_L){1'b0}};
               If745dbf2f0d756857eff51da036067fe  <=  0;
               I2c117c8ea4060a5094453cc6140c9bb6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I22231ac2204ad703262885231f7451e8  <=  0;
               I56a6be4115d52bd49fc003b164fbcdb0  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4e1e119c87f56b39ec6ddab9b160430d  <=  0;
               Ib834a7e4f3a491e351e2e49d809d2448  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9d9cc96988bd0af2b2c8682af3779794  <=  0;
               Ifdcb28209b39b8d99c2eb00a72921a75  <= {(MAX_SUM_WDTH_L){1'b0}};
               I027210d36e2ae38a39746ac6fde3129a  <=  0;
               Id721a94e50637fa39c5bf6124ecfae6f  <= {(MAX_SUM_WDTH_L){1'b0}};
               I28e32abf786d964b95d72bc17425a90f  <=  0;
               I72ee7b62c165dc693cc6b5185970f7f5  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id29266756e91fa3c40480f9cf22f1671  <=  0;
               I564ae36637e0cd6a8a06289e95823572  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iad31d6f7d366c849222593883210e817  <=  0;
               I085e99650c86078bf02f1b2aed141add  <= {(MAX_SUM_WDTH_L){1'b0}};
               I495d2cfe02637adf0bde6dd48201cedc  <=  0;
               Ie4e63cba44dee9885eeae32cc844c3f5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I544225b6c571710d59f804f082f475c8  <=  0;
               Ic054b062712da78ddd4a148bafeb1a0d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6f7ff2aeffdfe5bd4090ecd655ff5aa2  <=  0;
               I81b01fc018ad1c79ec03a123763e95d9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1783da96203ac6a00cd2e8f2dfe1ac34  <=  0;
               I1d38ff144c3dcfe4c04778e50a044d5e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I00ae9e980c05d6d55570d92582a80410  <=  0;
               I2e31a90886f87907d19d0c034caeee9c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I86282458466a079a1063e068011d58eb  <=  0;
               I7c48130cd79566b1f1e30b7c709ee5cb  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7dcde2729bcd8e63b86dcac06325887b  <=  0;
               I3868c6ed60d1f0ef9d3ad98e91931acf  <= {(MAX_SUM_WDTH_L){1'b0}};
               I31ca3f6f5d61b73718bbd9c19f7fd53b  <=  0;
               I7fa57873a108e5894f837bdf45979b8d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie01688869a15f6b506bc3fbdea78b6b0  <=  0;
               I59d4025a86d065a84741dafb86b50cbd  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iff748fa3440e5d0f80969f64b10eca98  <=  0;
               Ib28a3fb3dcdea36c883c88b017fefa56  <= {(MAX_SUM_WDTH_L){1'b0}};
               I85018196561b6ef22994dfff7e3a8b80  <=  0;
               I91e4dca55e1a5d1d8ddee5c3bd1048bc  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifff25101d23e8e0ac43d5f0507a34217  <=  0;
               I55dd62b8ff91323075533e896207c1e5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I261ed926e2e82b283ac24970f546a5fe  <=  0;
               Ia30ca84355bb976cd045e969b2862856  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ibf081c14165822b88553a913ba320016  <=  0;
               Ifa1359651fd7e160301261bdbb81b02c  <= {(MAX_SUM_WDTH_L){1'b0}};
               I595bd58339ea7427b88385a62835aab6  <=  0;
               I0b465f693268f6f56f52d41165bf66ef  <= {(MAX_SUM_WDTH_L){1'b0}};
               I41b82d4c805471097a0dd4f85615f990  <=  0;
               I3deffa3a53b31688f28dfbfa66571d0c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie07ed8367e7b83324c539bddcb3b1dfd  <=  0;
               Id40c9857a5bb6c8cdc616fe68d8dc39d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I67ba6804ea940c34c7c588832272581e  <=  0;
               I26754124b13858a3b925cddca5cd8c5b  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifb2d4794b0630c3cdecb6cd2d2b1b384  <=  0;
               I2ebc1a7d32a5457de4d35b6bb25507d1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I9c6dda8e9e0d7e69032a1fb40684c87c  <=  0;
               I77bf5b03fa300d1dbf8df5ca4acbed14  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie7d857b468dedb6b7a73fe918332ff1d  <=  0;
               I6c1c1e404f92fc80495e8e5d187934a6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I34662a12c505be8abbe01cb690d117d5  <=  0;
               I126a2b15cdc34d88d17ebacb3681625f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idc13433074453a726e7a35789d7d27d2  <=  0;
               I9c5ec8e21febe3ebe00c53ac8b21d1f1  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id16d40761b18218d4270c00db6d4eca2  <=  0;
               If27eaa7cc4d1b5d2b7a962b48f0919df  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifac93c987a8fb9726d85b77a2e4c8bba  <=  0;
               Ic15f443512d68537f9764a3ba88334f6  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id742302a78483bbb2852b002262ed33d  <=  0;
               I47b266262fb5a98f66706f460f1248e6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I2f87df8d48fe83aa0ce493d69aaa3d88  <=  0;
               Id301f31702270a4f8e9964e3a75e3d62  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic4bb880cb9f8d5a6d1cbbdf7cd205470  <=  0;
               I097ba3ae5a0232ae6aa35478635640b3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I369ea36c9da8f4c9b93ee70f8d4c149f  <=  0;
               I3b65eb49005aee57f61279c5a172d158  <= {(MAX_SUM_WDTH_L){1'b0}};
               I17f6c250d2d07a58ddde6d232a1ab5de  <=  0;
               I8573059885be4373531275502affd59d  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iba5b23512434eb51ec8679a798273551  <=  0;
               I627f9d9ac0c07ded7306fd14773fbee4  <= {(MAX_SUM_WDTH_L){1'b0}};
               I91a06282a09b01980f2e7be4ecd3a982  <=  0;
               Ib559f45098803b21622fa96ade885abc  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1b928fa95275de94960b3e2b4d67338b  <=  0;
               I10e294379879538ecbf65fd423e7355d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6488c30acdb3b47d4d4ee7b5947abdfe  <=  0;
               Ice861034cd3b2f3847f325dbc9f52d08  <= {(MAX_SUM_WDTH_L){1'b0}};
               I29a436013f98b750df592eb7d26d0d1e  <=  0;
               If201eea7e0023bb17fe41dbb4b5ec076  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6fb12e6f50ffa6e94c9d43a22681702c  <=  0;
               Ib15f9bf401d734008d6a2b9a00c572d1  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib3f42f17505d5c091c8c924bbc26d117  <=  0;
               I581f4e137ec21e639eec32a1675f4750  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia4c22a118187d5b2dd154a4371dc06d1  <=  0;
               Ib7ff7b93c88fc8d9bcd915f0c678acff  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1a87822c50f6a0ac5a5e96021ad49fb3  <=  0;
               I34dc9dff97e78a2d711f75675944b0d1  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6addbc7c163ce97b3482277e76c5feaa  <=  0;
               I8bc35065fe56bb75e6595937aaf9ef2a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I124c4374f19808abbdc401a3b85aec67  <=  0;
               I1822ab8ed690d872380ef820dc4282fe  <= {(MAX_SUM_WDTH_L){1'b0}};
               I162653d33938a4553978b08df208228b  <=  0;
               I1a1965726584c6c91a7e20de63f0fce3  <= {(MAX_SUM_WDTH_L){1'b0}};
               I291a3bbec5669b8958c0ded154af1f89  <=  0;
               I08c5dcac6674c1671b85d07a55a005b0  <= {(MAX_SUM_WDTH_L){1'b0}};
               I53a1d11cce6e036ba3a23dcc29d1cc3e  <=  0;
               I40d67287bf525ab2696c30755d6babd5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I5fda5f3c582bb88cb7de87298d15194a  <=  0;
               I60dc8e5b6204e3a5fa32e79c5cceae94  <= {(MAX_SUM_WDTH_L){1'b0}};
               Id3933d661bcebbc3584c9e437c96c89d  <=  0;
               I0074b447046d75787aa872d8167171aa  <= {(MAX_SUM_WDTH_L){1'b0}};
               I0d38a30070a5ae3e879c357c3dde88ea  <=  0;
               I384965816ec3b915b9b623ad68fcc4c9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I928993ece796543b23fb83df8c250845  <=  0;
               Ic0e2656bee7174384f7f952dbb9da619  <= {(MAX_SUM_WDTH_L){1'b0}};
               I226f8490438d72f58c43377c8e60fc34  <=  0;
               I4cc3b0546ddc14d78da59e4981a77b58  <= {(MAX_SUM_WDTH_L){1'b0}};
               Idaefaba16ce80e24f16df683cc83d759  <=  0;
               I7b680caf7d0d94114fae1d96ba374e68  <= {(MAX_SUM_WDTH_L){1'b0}};
               If1da75cd8208f606c1b121f441685cbb  <=  0;
               I7f8986a922c03b6afb5786cd2e1d5288  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib63f66960a3981879aad950588ea14be  <=  0;
               Ie7814643e3833736c0f54b39f91fe792  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia2c2ecedc809186e3f9224a9aa4bf385  <=  0;
               Id1f0c95b85ee041818da4fd9b5466c7d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1fc189d6e8a90cc0033c6e690916de83  <=  0;
               Iefa8421c0c908de69fccffbe22f40911  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7fa18d2c7159b9fda8957384ebca5700  <=  0;
               I4319bf1bbb31debc7f58157b75025134  <= {(MAX_SUM_WDTH_L){1'b0}};
               I7ea0274f5b34aac64a17fa9171201a5a  <=  0;
               I4a349021efeeda16b646979a959bff6e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8d26db6f54d068f798e2951701aebed1  <=  0;
               Iaae0c136077ecc36fc382a76abd550e7  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8fb8a6e1ab4647e8e1dda4da8b3ef3c6  <=  0;
               I4a442564148493664046e7b38cc6cfe4  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie4821dad77dec0567d64f7c1de7710af  <=  0;
               I12cc5eec3de8ceb3ca084194d430d9a5  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ic4d741a90fcc86f31eb3567d028eb27f  <=  0;
               I56db71b7df11c35080cbaee80c389c59  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1d2641b8888a0f7b4b78cae16779da75  <=  0;
               Ifd1431230378775456efa4bdd5bfc397  <= {(MAX_SUM_WDTH_L){1'b0}};
               I48badf0536ab133751d4be1e0450fd81  <=  0;
               I6f0cef6d870e38e5ba192463a3920818  <= {(MAX_SUM_WDTH_L){1'b0}};
               I043ba9e5157ad18a4e466df0540b79ba  <=  0;
               I3ee87c05f23571b687611fdce84a1b91  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib9760b69084b2d4a3a93126e5da0f20b  <=  0;
               Ide521f7523b897bb6fb747202f730ac5  <= {(MAX_SUM_WDTH_L){1'b0}};
               I4978a011cb09d68ac2850e1f515d7e88  <=  0;
               I314b64e5fbbc14807fd7fe3c7bca101f  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib09ea18232dfca23f3f139438e6cb800  <=  0;
               Id5ad2e12b160bc6a9f96f2524f849c8e  <= {(MAX_SUM_WDTH_L){1'b0}};
               If29c61ebd2b452efe995c212a76a77a0  <=  0;
               I2b2bf6d4e879b8f53b02f94f1e964344  <= {(MAX_SUM_WDTH_L){1'b0}};
               I60fa2e2b5dd8b0a99612d2f2f6c5c740  <=  0;
               Ic60cb038b4b90d8035059b1e06f8d765  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ifc9b6cc64f5bf8bc685911bb28884a0e  <=  0;
               I707e2d6d9807076bfc91417fb9e198e6  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1aeaa36994ba29298931735d5a1237e0  <=  0;
               I49f5797b92e17562e6dfde42c20c7a37  <= {(MAX_SUM_WDTH_L){1'b0}};
               I415ed6a9802acf39be10b220ddb3ff66  <=  0;
               I0a9f0274dc61d574c40e0e2048fb0b9e  <= {(MAX_SUM_WDTH_L){1'b0}};
               I1c06321ed28c991ad2aa8a3725769dee  <=  0;
               I53ae3de5769255a9e69a2ae690d44ba9  <= {(MAX_SUM_WDTH_L){1'b0}};
               I198d5b5bf8f39f9bd6b2f4c993fd58ca  <=  0;
               I1390f0ff082dbff11a64cdfcbe1b681d  <= {(MAX_SUM_WDTH_L){1'b0}};
               I3bf64d0a85c83de954a286e6afa8f727  <=  0;
               Id2f8816659d3881ee1b1d14668a53a08  <= {(MAX_SUM_WDTH_L){1'b0}};
               I897c7fc822d490f69b531a8f749815f4  <=  0;
               I286bacc5a8a77b89cb99dbb00962555b  <= {(MAX_SUM_WDTH_L){1'b0}};
               I6c7cb10db83156b49d46fab38d0f9fc5  <=  0;
               Icda8e8a6ba7607752ed282114a542b67  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ie47af3b071351ec683abe28b7fe2b642  <=  0;
               I2da4a59f9a6bd71af95790a75b172df0  <= {(MAX_SUM_WDTH_L){1'b0}};
               If2dd4df3af6446c05da4afdaa7e92cab  <=  0;
               I1bcf01b7fde13919f5d7c4df4483e61c  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iabf085ea078abe8748810e81a6d03cac  <=  0;
               Id5f000c37734979d057f7887739a5615  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ia2ae348906a599a4d327ff1419315afb  <=  0;
               Ibccd7142ba951dadbeca13178458bb3a  <= {(MAX_SUM_WDTH_L){1'b0}};
               I18df34aea04ea7dc99fc918892bf8f0e  <=  0;
               Ic1fe6b93bc8d517686ba430d3d1fe7ab  <= {(MAX_SUM_WDTH_L){1'b0}};
               I910749abcd809e1c730f27fb5e1ddab1  <=  0;
               Ib1c8d1d733e91f052f6d6824e734b1e3  <= {(MAX_SUM_WDTH_L){1'b0}};
               Iae95ea2f32f53a5060c0199c8196d681  <=  0;
               I08348d0a177e264af1a4769422878a06  <= {(MAX_SUM_WDTH_L){1'b0}};
               I8c3d927ec93e73c5bca489a2f2b43f55  <=  0;
               I2d2c2997dcc5167fc6ddc1e90f0ebc49  <= {(MAX_SUM_WDTH_L){1'b0}};
               Ib41ff881898782965734bb0cc333be79  <=  0;
       end else begin
            // Id66554a95b5375bec1ec7c8e6bbfea7d and I8fee031b61092657fa6474c0ef478763 I55f195813a158d82e2934cfac569575d I12de3a4dab98ef8a7d67aace8150b540 Ied2b5c0139cec8ad2873829dc1117d50 I51037a4a37730f52c8732586d3aaa316 I05531b19bb846b18c09f979eeb429ad3
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f == I40a85f3ef46def30cd7707afd2c7fa44 ) begin
                    I18d11d94a39d5d7687736d266d3e1902  <= Ifeb14203f4daf31c7701a6a742be57cc;
                    Ib64114b4af6a37b3d52bd38cb83459ee  <=  0;
                end else begin
                    I18d11d94a39d5d7687736d266d3e1902  <=  ~Ifeb14203f4daf31c7701a6a742be57cc + 1;
                    Ib64114b4af6a37b3d52bd38cb83459ee  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f == Ib8963a4ab143aba7fadc61d89f937f4e ) begin
                    I6b9ffa985ece553b83f7227e7a85141b  <= Ib581c19864deecf01268595049268b19;
                    I06ed412c4554e98837146a5c7a6c4789  <=  0;
                end else begin
                    I6b9ffa985ece553b83f7227e7a85141b  <=  ~Ib581c19864deecf01268595049268b19 + 1;
                    I06ed412c4554e98837146a5c7a6c4789  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f == I9565de7442acee8455d1c4f8ab43ab07 ) begin
                    I49fdba80df1c667dd264e5105a530332  <= I661d84af541e30828bcbd962d72baba3;
                    Iefa11849e46b6ccd923e622fdb878315  <=  0;
                end else begin
                    I49fdba80df1c667dd264e5105a530332  <=  ~I661d84af541e30828bcbd962d72baba3 + 1;
                    Iefa11849e46b6ccd923e622fdb878315  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f == I26b11eb80b9a1752998f7ab1379e4124 ) begin
                    Ibf4fc04c9e0aa536a8e4b8a6192d8498  <= I1c6928cccb4bf7ea7dfd74e425b9624d;
                    Ia4245ce0efa56b1234283f4969246280  <=  0;
                end else begin
                    Ibf4fc04c9e0aa536a8e4b8a6192d8498  <=  ~I1c6928cccb4bf7ea7dfd74e425b9624d + 1;
                    Ia4245ce0efa56b1234283f4969246280  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f == Ibb068f313ff784191769e8da44f023e1 ) begin
                    I899abb7dcba235ff2afb410a87e16973  <= I6eabc5c074fb1e2183a5f1ecee87a518;
                    I671b766473f67c92b75716e2bd9a9596  <=  0;
                end else begin
                    I899abb7dcba235ff2afb410a87e16973  <=  ~I6eabc5c074fb1e2183a5f1ecee87a518 + 1;
                    I671b766473f67c92b75716e2bd9a9596  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f == I2348d423bff186f1841ecaaf44f4f2c6 ) begin
                    Iab322f0da75316ca9937802a327dd537  <= I0107769bbd7c239685b4818731334437;
                    I24b5cce7252356b606027b301ac6bf48  <=  0;
                end else begin
                    Iab322f0da75316ca9937802a327dd537  <=  ~I0107769bbd7c239685b4818731334437 + 1;
                    I24b5cce7252356b606027b301ac6bf48  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f == I3b28138cac28625778c34d4bb1a4aa55 ) begin
                    Iba0a4530bce787d70253a92c123f589e  <= If723180430080198d18a08d6775ab208;
                    I2f0d19d012f0bd45308356fce1a50049  <=  0;
                end else begin
                    Iba0a4530bce787d70253a92c123f589e  <=  ~If723180430080198d18a08d6775ab208 + 1;
                    I2f0d19d012f0bd45308356fce1a50049  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0973b6e90e7678addcb064fded7ce0f == I8928563d2510725797f96917767f9bae ) begin
                    I4475d6a1e59d35444a6a2d9647c6761a  <= I44abc734d6acf92a8e8209186d7a1676;
                    I939c483ddfc18ee8dca73a1c98e6ec4d  <=  0;
                end else begin
                    I4475d6a1e59d35444a6a2d9647c6761a  <=  ~I44abc734d6acf92a8e8209186d7a1676 + 1;
                    I939c483ddfc18ee8dca73a1c98e6ec4d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iee06707670e19a82d911c1750bcfc811 == I989726d5ee5f23a016e85b0945573f05 ) begin
                    I217e2e1eb3404ba9ff06d284a18256b6  <= I72aa55988d58c664f3291b5786fc8ceb;
                    Ife63de208f77b322e1c885e78790f997  <=  0;
                end else begin
                    I217e2e1eb3404ba9ff06d284a18256b6  <=  ~I72aa55988d58c664f3291b5786fc8ceb + 1;
                    Ife63de208f77b322e1c885e78790f997  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iee06707670e19a82d911c1750bcfc811 == If88711683bd32856ce45937b841581e3 ) begin
                    I2003418e663144ee49f1ed044f6a0062  <= Ie69528583db8155917ab3d32a446de04;
                    Ia065f925c78015a3736219a5c7129439  <=  0;
                end else begin
                    I2003418e663144ee49f1ed044f6a0062  <=  ~Ie69528583db8155917ab3d32a446de04 + 1;
                    Ia065f925c78015a3736219a5c7129439  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iee06707670e19a82d911c1750bcfc811 == I015cf78df7e3417d5296eb0ad3019674 ) begin
                    I4496255218b6d0f5374328803aeeb412  <= Ib22b47d95b72871e74069fe80a191680;
                    Ie02e0e9e2627b178d6c54ea743b3993b  <=  0;
                end else begin
                    I4496255218b6d0f5374328803aeeb412  <=  ~Ib22b47d95b72871e74069fe80a191680 + 1;
                    Ie02e0e9e2627b178d6c54ea743b3993b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iee06707670e19a82d911c1750bcfc811 == I31908b38609b532f9f142a97e0442e55 ) begin
                    Iecbb3f290db6dad3393b592ca946fa13  <= Id9451e945bd26b8dcb4cb83ab4ade73b;
                    Ib1e432e0b2d7979227d2cc591ed8e383  <=  0;
                end else begin
                    Iecbb3f290db6dad3393b592ca946fa13  <=  ~Id9451e945bd26b8dcb4cb83ab4ade73b + 1;
                    Ib1e432e0b2d7979227d2cc591ed8e383  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iee06707670e19a82d911c1750bcfc811 == Ib98eadb333ebca2f58c40b8f93d87250 ) begin
                    I9f88e23f2a17035b31840356a5d0bfde  <= Iba4627d3d3ef91f168068ed128c04113;
                    Ib05aef46725afee38240d81738c673f1  <=  0;
                end else begin
                    I9f88e23f2a17035b31840356a5d0bfde  <=  ~Iba4627d3d3ef91f168068ed128c04113 + 1;
                    Ib05aef46725afee38240d81738c673f1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iee06707670e19a82d911c1750bcfc811 == I4a0f0579aa9b7af7b516780074ca6560 ) begin
                    I3fd4a13843fc09ca68b827a8b09e6c49  <= I39bef4d462b0a3f88ce1485a58d66da0;
                    Ie7bea07eac0dc36dbce430e6dd088b5e  <=  0;
                end else begin
                    I3fd4a13843fc09ca68b827a8b09e6c49  <=  ~I39bef4d462b0a3f88ce1485a58d66da0 + 1;
                    Ie7bea07eac0dc36dbce430e6dd088b5e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iee06707670e19a82d911c1750bcfc811 == Iaebca9b574d490aeab28fbbfb1e8fd9a ) begin
                    I1530e79da3803bb87787397f19822dbb  <= Ib95e457d5ae9fc89e197c249414abbcd;
                    I3f42e9b5ae0fc5c9315670cad33374ce  <=  0;
                end else begin
                    I1530e79da3803bb87787397f19822dbb  <=  ~Ib95e457d5ae9fc89e197c249414abbcd + 1;
                    I3f42e9b5ae0fc5c9315670cad33374ce  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iee06707670e19a82d911c1750bcfc811 == I3ad613d80a126f03fb9125fe6da1bc8d ) begin
                    I613821692bb99a8a6739d3c3ab7211ac  <= I2be28be47a38e9ca9d3b9167327d3d59;
                    Ie6f54d5d349ba8e19295a9ce17ba3f35  <=  0;
                end else begin
                    I613821692bb99a8a6739d3c3ab7211ac  <=  ~I2be28be47a38e9ca9d3b9167327d3d59 + 1;
                    Ie6f54d5d349ba8e19295a9ce17ba3f35  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd == Ic116b21b5744ec42a9f41eff3ddd1707 ) begin
                    I5ac600834d567934bd2f0b14a3c38ab9  <= I2ee6154b613d0d86c2354604e93a9a57;
                    Iab7ce2d8e89a5862f98bd812751d1d17  <=  0;
                end else begin
                    I5ac600834d567934bd2f0b14a3c38ab9  <=  ~I2ee6154b613d0d86c2354604e93a9a57 + 1;
                    Iab7ce2d8e89a5862f98bd812751d1d17  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd == Id9f7e6885737ee2d3128081915a685b0 ) begin
                    I84fe1a1ecad408b16557957b01cc94b9  <= Ia7479d4940b575cf918cb8421f041e44;
                    I8a4157cd8206e66109f979bd9bde53b6  <=  0;
                end else begin
                    I84fe1a1ecad408b16557957b01cc94b9  <=  ~Ia7479d4940b575cf918cb8421f041e44 + 1;
                    I8a4157cd8206e66109f979bd9bde53b6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd == Iad36872fbd9ac694d47cc0491f3d021e ) begin
                    I7d03cdddc264c89446cd80405c34d69a  <= I3c5b1cddd608ad869e0182ad68bd0494;
                    I5f0937deee06e2177807a6d0fbc2e2b0  <=  0;
                end else begin
                    I7d03cdddc264c89446cd80405c34d69a  <=  ~I3c5b1cddd608ad869e0182ad68bd0494 + 1;
                    I5f0937deee06e2177807a6d0fbc2e2b0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd == I0794dcad0f96cf58fda60c561a1144fe ) begin
                    I5cf7e3cb90e84c3ac6a66fb6dde220af  <= Ic4425ae997c479e05e12347a803213dd;
                    I598fa274e3ada377f2e7a43d7dfd9231  <=  0;
                end else begin
                    I5cf7e3cb90e84c3ac6a66fb6dde220af  <=  ~Ic4425ae997c479e05e12347a803213dd + 1;
                    I598fa274e3ada377f2e7a43d7dfd9231  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd == I8b4cdd738b1ed431764d4a51be668460 ) begin
                    I602c2e5bfa93cb3c87af70dd69b0375d  <= I3a0518d0d382758ae579acd7e6cd634a;
                    I4a3da449219c7068a0bfd3a192d2ead1  <=  0;
                end else begin
                    I602c2e5bfa93cb3c87af70dd69b0375d  <=  ~I3a0518d0d382758ae579acd7e6cd634a + 1;
                    I4a3da449219c7068a0bfd3a192d2ead1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd == I79e67c70ee26ab7623355ec5042dcb28 ) begin
                    Id50fe525d660f0bb0ac3bbe6e68758f1  <= Ifd28c1cd286b7a483891bdd094b70db1;
                    Ia7a0522cea2126afdae3fb9f123d51fb  <=  0;
                end else begin
                    Id50fe525d660f0bb0ac3bbe6e68758f1  <=  ~Ifd28c1cd286b7a483891bdd094b70db1 + 1;
                    Ia7a0522cea2126afdae3fb9f123d51fb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd == Ie0a573c73ca9198012dc8ff4f8373973 ) begin
                    I6a68067b177340dbea2c53f7d8bd5f14  <= Iadf7734be049c645819d9d023b58c4dc;
                    I5d901ed468b60a31e199d12612a0b396  <=  0;
                end else begin
                    I6a68067b177340dbea2c53f7d8bd5f14  <=  ~Iadf7734be049c645819d9d023b58c4dc + 1;
                    I5d901ed468b60a31e199d12612a0b396  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id8d5df9e869aaeb107a41a6bca3b89bd == I6a4cd5680e34df5ccfea4a7eb72113ec ) begin
                    I9efdcdeee8883d30159881f8831a2c03  <= I5f23af0d0853ea6de084ccf77702b78d;
                    Iceced38b8b522d1679ed4e1cad38c282  <=  0;
                end else begin
                    I9efdcdeee8883d30159881f8831a2c03  <=  ~I5f23af0d0853ea6de084ccf77702b78d + 1;
                    Iceced38b8b522d1679ed4e1cad38c282  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I507f8602a99a1096e4c293ba3c235bbb == I9885460698fe454e65fea4a6022e5df0 ) begin
                    I46290d63552b8cac8d22358cb38c5887  <= Ic5c99c42e9ebe5dded369ac78a1bedb5;
                    I7d3d6075ca3828a533b52dc3cac3a652  <=  0;
                end else begin
                    I46290d63552b8cac8d22358cb38c5887  <=  ~Ic5c99c42e9ebe5dded369ac78a1bedb5 + 1;
                    I7d3d6075ca3828a533b52dc3cac3a652  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I507f8602a99a1096e4c293ba3c235bbb == Iee7e507956faf7cd903ac2dd636b7819 ) begin
                    I6435c7b1b3bfc5dae42cb1b3b03aefc5  <= I4f2498bec0e96802b82f0419d97c527f;
                    I0869d337e6cce62a05b29c5baa4ed436  <=  0;
                end else begin
                    I6435c7b1b3bfc5dae42cb1b3b03aefc5  <=  ~I4f2498bec0e96802b82f0419d97c527f + 1;
                    I0869d337e6cce62a05b29c5baa4ed436  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I507f8602a99a1096e4c293ba3c235bbb == Icece56258c1ffa7a0257d68ef9ff5ee7 ) begin
                    I63b2f1c2148e595a40bb41968e4b9a65  <= Icaf86e0abee612aa972388c0b6f90763;
                    I36ae963a57878d2c5b647910e003dea0  <=  0;
                end else begin
                    I63b2f1c2148e595a40bb41968e4b9a65  <=  ~Icaf86e0abee612aa972388c0b6f90763 + 1;
                    I36ae963a57878d2c5b647910e003dea0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I507f8602a99a1096e4c293ba3c235bbb == I6c15ea618986f2043f402959ac23fb1b ) begin
                    Iafb6296c59c2dd241c880c6d57352617  <= I478c4f13c05651605a2045bb5fd6b60d;
                    I5851ca9a7e932378c2bdf2c118b498dd  <=  0;
                end else begin
                    Iafb6296c59c2dd241c880c6d57352617  <=  ~I478c4f13c05651605a2045bb5fd6b60d + 1;
                    I5851ca9a7e932378c2bdf2c118b498dd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I507f8602a99a1096e4c293ba3c235bbb == Ic45cade04982e60abe32a359999a778d ) begin
                    I0b982beca6221db7b3ec2afb3833a60e  <= Ide67911b52687d67ef0c25f2aadf14c5;
                    Ia5597b68eb3f1c1d371cda63fa1fe034  <=  0;
                end else begin
                    I0b982beca6221db7b3ec2afb3833a60e  <=  ~Ide67911b52687d67ef0c25f2aadf14c5 + 1;
                    Ia5597b68eb3f1c1d371cda63fa1fe034  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I507f8602a99a1096e4c293ba3c235bbb == I670dbb51097dde1f56eeb7e25ac50369 ) begin
                    Iece8968796771c1ef094808823da8962  <= Ie9e7630af25f39a0e820181918edd029;
                    Icc939d3c403d238cf5c9c196cac91886  <=  0;
                end else begin
                    Iece8968796771c1ef094808823da8962  <=  ~Ie9e7630af25f39a0e820181918edd029 + 1;
                    Icc939d3c403d238cf5c9c196cac91886  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I507f8602a99a1096e4c293ba3c235bbb == Ia3fb4901b185e64ccb788dcc1d7cfb1b ) begin
                    I05c7cb4a076239b8976a76d418ad6149  <= I0e1f07f30cfe36f189e9dcb4e713b5c8;
                    I0bd90c7dbb94917bb46a3e008484f582  <=  0;
                end else begin
                    I05c7cb4a076239b8976a76d418ad6149  <=  ~I0e1f07f30cfe36f189e9dcb4e713b5c8 + 1;
                    I0bd90c7dbb94917bb46a3e008484f582  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I507f8602a99a1096e4c293ba3c235bbb == I15a23e6922630f6d409706b1c4100d22 ) begin
                    I9076162e7b10bffbc9473e35b407e986  <= I31cee5e2a93635987776b0ea477e6211;
                    I6ec7620a49b53a8377767e363e88d471  <=  0;
                end else begin
                    I9076162e7b10bffbc9473e35b407e986  <=  ~I31cee5e2a93635987776b0ea477e6211 + 1;
                    I6ec7620a49b53a8377767e363e88d471  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == I08eb91ffc153d5007de61e2938407d18 ) begin
                    If702042844ed38f5e7103382ef4263eb  <= I84721f2bc5ae10db78d2e7e07cc28d94;
                    Ie512ccdcaff0cc5c29277e28f1ba5fa8  <=  0;
                end else begin
                    If702042844ed38f5e7103382ef4263eb  <=  ~I84721f2bc5ae10db78d2e7e07cc28d94 + 1;
                    Ie512ccdcaff0cc5c29277e28f1ba5fa8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == I642d63513e039da95a66c1cd4336f84f ) begin
                    Ide63b2762649761944db237c8efe69ae  <= I6c6d057e910da53aa47441566f95153e;
                    Ia115f92bd6dcb4167f0771941a18ad59  <=  0;
                end else begin
                    Ide63b2762649761944db237c8efe69ae  <=  ~I6c6d057e910da53aa47441566f95153e + 1;
                    Ia115f92bd6dcb4167f0771941a18ad59  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == I1e35f6f8ac9e61787a3b263e5e4ac62c ) begin
                    I1cec628c6d6e22895a0f0c0258851171  <= Iecbf70768fbaaab8da98eaa9a2b956ee;
                    I7c8174a3579ed90c0ec89941ac53e287  <=  0;
                end else begin
                    I1cec628c6d6e22895a0f0c0258851171  <=  ~Iecbf70768fbaaab8da98eaa9a2b956ee + 1;
                    I7c8174a3579ed90c0ec89941ac53e287  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == I5af04bd644d9c14f56884acd1f6674a7 ) begin
                    I46b0b74552e89df91c0027f0f093e1f5  <= I71b8492d70b423e95938995c07395def;
                    I7d6b68dbc5ac773ce97df3a6726c6836  <=  0;
                end else begin
                    I46b0b74552e89df91c0027f0f093e1f5  <=  ~I71b8492d70b423e95938995c07395def + 1;
                    I7d6b68dbc5ac773ce97df3a6726c6836  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == Ia9bc04087c3926bdf993858e683dc3f6 ) begin
                    I68dbff67a1910346ddc0281b445f4439  <= Iae469bcbba9598bb46aa7ccf9fa06a37;
                    I5045f1311d1e891577f3f8a09078fe79  <=  0;
                end else begin
                    I68dbff67a1910346ddc0281b445f4439  <=  ~Iae469bcbba9598bb46aa7ccf9fa06a37 + 1;
                    I5045f1311d1e891577f3f8a09078fe79  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == Ia8c23f2c6c80bc389fd66aee524975cf ) begin
                    Ia42f547c0b02c2de66f2ff383ca1741b  <= Ie2e854376f4b6509ec41507401173269;
                    I105c3326421f25d3b9931e2178c794d4  <=  0;
                end else begin
                    Ia42f547c0b02c2de66f2ff383ca1741b  <=  ~Ie2e854376f4b6509ec41507401173269 + 1;
                    I105c3326421f25d3b9931e2178c794d4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == I74ff51ab0824be97bf311b50b4ce5401 ) begin
                    If456045711d535cea07d9dd5ef9b04c6  <= I7b1401c3c2c389d9bf05658c88ff6b40;
                    I838c5c183e758ef4f28ad86d16befd87  <=  0;
                end else begin
                    If456045711d535cea07d9dd5ef9b04c6  <=  ~I7b1401c3c2c389d9bf05658c88ff6b40 + 1;
                    I838c5c183e758ef4f28ad86d16befd87  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == I22cf21c1e88c0b8ff5d5b43835b1f61f ) begin
                    I9585ff28ce0f3bca71d582b1cb8937d7  <= I88ee95aeb6c744eca0e127e8497b5dc9;
                    I33c782b29a89c2ec375038b88919b564  <=  0;
                end else begin
                    I9585ff28ce0f3bca71d582b1cb8937d7  <=  ~I88ee95aeb6c744eca0e127e8497b5dc9 + 1;
                    I33c782b29a89c2ec375038b88919b564  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == I2fc87e59765765e16bae0761ab5741ec ) begin
                    Iac3dfb28a343cbb391fdf58684e091ef  <= I5573e18ade3430ef3eff5e6d960e44eb;
                    Ia21ec0ad85852d1eea449283d1d45a7c  <=  0;
                end else begin
                    Iac3dfb28a343cbb391fdf58684e091ef  <=  ~I5573e18ade3430ef3eff5e6d960e44eb + 1;
                    Ia21ec0ad85852d1eea449283d1d45a7c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibdf2178bd18783c4797c21e642388d16 == I6c6297e7aca3c7d8a9f8c3542f8b070c ) begin
                    I82650d4bf0a9b51e245665259f40fe60  <= Id6260fa8a9be077673e82344c736b1c4;
                    Iae32e0aebc2719c3e476a5300f1bfdea  <=  0;
                end else begin
                    I82650d4bf0a9b51e245665259f40fe60  <=  ~Id6260fa8a9be077673e82344c736b1c4 + 1;
                    Iae32e0aebc2719c3e476a5300f1bfdea  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == Ifbc2ba75815cb3aece1d327a5c15dba4 ) begin
                    Ib21e67aa9696222891a0b33c414b1bbd  <= Ic052eadb342350c52d89e73d5fea80bb;
                    I6914a92b8da6d6db6f2e8806c7efc5aa  <=  0;
                end else begin
                    Ib21e67aa9696222891a0b33c414b1bbd  <=  ~Ic052eadb342350c52d89e73d5fea80bb + 1;
                    I6914a92b8da6d6db6f2e8806c7efc5aa  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == Ib1bba2d65c2224f05a444c6170aba187 ) begin
                    I1e168bf1a0dd18ff31d3560be00095f1  <= I98b8d024432fc54ebf2f15d99968f2e0;
                    I60cad827424e4799360141222a80ac57  <=  0;
                end else begin
                    I1e168bf1a0dd18ff31d3560be00095f1  <=  ~I98b8d024432fc54ebf2f15d99968f2e0 + 1;
                    I60cad827424e4799360141222a80ac57  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == Id75ce45a6df04b3d173b288b52d82138 ) begin
                    I97e6d2bc8c1ad455f7c61de81e8d4826  <= I98f54ab8454940141a484332f2a05369;
                    Ie3389948b5dd781ac9087e62cf93dd2d  <=  0;
                end else begin
                    I97e6d2bc8c1ad455f7c61de81e8d4826  <=  ~I98f54ab8454940141a484332f2a05369 + 1;
                    Ie3389948b5dd781ac9087e62cf93dd2d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == Icd148cb7a25bc30aafd0271e00356527 ) begin
                    Ie1170db51d408ccc7360ce53c94a9644  <= I9d94ad2da06ac1fef4da7dcc56abffca;
                    I566475d003c9fc40aebaba87655a0668  <=  0;
                end else begin
                    Ie1170db51d408ccc7360ce53c94a9644  <=  ~I9d94ad2da06ac1fef4da7dcc56abffca + 1;
                    I566475d003c9fc40aebaba87655a0668  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == I80e8b0fdd6bfadac9c8a788bd9be4b97 ) begin
                    If58c2c1e1dffe04295f3313595ffe319  <= I51262e3abe460148e3c2d2b74989c2b8;
                    Idb2467b1104f5b924d419208f2573df4  <=  0;
                end else begin
                    If58c2c1e1dffe04295f3313595ffe319  <=  ~I51262e3abe460148e3c2d2b74989c2b8 + 1;
                    Idb2467b1104f5b924d419208f2573df4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == I471dd2bc897a40a9463f4984952d4fa6 ) begin
                    I9a9fb4da9fdf5bd42cef32c7d8fa65d9  <= I560583680bb2f5a0b5ede42ceaafcf8b;
                    Ie0a8d219223bc68ea3040cbbd349caac  <=  0;
                end else begin
                    I9a9fb4da9fdf5bd42cef32c7d8fa65d9  <=  ~I560583680bb2f5a0b5ede42ceaafcf8b + 1;
                    Ie0a8d219223bc68ea3040cbbd349caac  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == Ic61bade7088606659ef8568dc134f686 ) begin
                    I785e4a1f2556289db0bd024e429bbd3e  <= I389f83346ffaffe8186fb0074d71f43c;
                    Ide01b9dcf3a3019d689d79f4d7ce0f32  <=  0;
                end else begin
                    I785e4a1f2556289db0bd024e429bbd3e  <=  ~I389f83346ffaffe8186fb0074d71f43c + 1;
                    Ide01b9dcf3a3019d689d79f4d7ce0f32  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == I298e98803772a458fbeed1de632c0555 ) begin
                    Ib6ca0cbcbaadb956d19a482fc099b175  <= Ie89c2a1b3943d12197bb972bd12595b0;
                    If33bbe9993ff895a7bd07bb8ee4ca970  <=  0;
                end else begin
                    Ib6ca0cbcbaadb956d19a482fc099b175  <=  ~Ie89c2a1b3943d12197bb972bd12595b0 + 1;
                    If33bbe9993ff895a7bd07bb8ee4ca970  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == I605674982abba50698d4d3c2220b0db8 ) begin
                    Id52b94ae6662bb2137d8b9d53280bcdd  <= Ic7be56919976a2d1088114c21c3c1ffb;
                    If9a84cb15af69dab2d9e4ed921f4deab  <=  0;
                end else begin
                    Id52b94ae6662bb2137d8b9d53280bcdd  <=  ~Ic7be56919976a2d1088114c21c3c1ffb + 1;
                    If9a84cb15af69dab2d9e4ed921f4deab  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2c690809d9b9e3482fe5a133b5c00afa == I201d44bd3cdf2b34fd2564188190b27b ) begin
                    Ic3975e4171d618ba53e1569e4fc93440  <= Icb5dab0df062ab46bd3d1a73e85ef4c2;
                    Ieba9f76cfb4c1a8069e2bfae0320ab0d  <=  0;
                end else begin
                    Ic3975e4171d618ba53e1569e4fc93440  <=  ~Icb5dab0df062ab46bd3d1a73e85ef4c2 + 1;
                    Ieba9f76cfb4c1a8069e2bfae0320ab0d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == Ia764576ce7e8ec4fc7120bcb8c038422 ) begin
                    Ib4e0f05afd881adf14a5eab850c75a3b  <= I27a568cfc2df13cf689d366a25e5d05f;
                    Ic85dfb2e44272dea346bdb4352a88c44  <=  0;
                end else begin
                    Ib4e0f05afd881adf14a5eab850c75a3b  <=  ~I27a568cfc2df13cf689d366a25e5d05f + 1;
                    Ic85dfb2e44272dea346bdb4352a88c44  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == I66d5eccef31484a090c91507a3d38a85 ) begin
                    Ifb875d675aa28de930d889ae4d37b48e  <= Ia6688964078f1ea87b742352877aac45;
                    I9f0f8b22b39af997db900c486fc37a18  <=  0;
                end else begin
                    Ifb875d675aa28de930d889ae4d37b48e  <=  ~Ia6688964078f1ea87b742352877aac45 + 1;
                    I9f0f8b22b39af997db900c486fc37a18  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == I93cee05370c836746d1ddeb0f74456bb ) begin
                    If98948e5f60b2c3ba1d7338e24dc0df6  <= I180deab4fe0d03104cf2ee035f6a9b8c;
                    Iebc1dd048a5c7e83175ba1030a4bb587  <=  0;
                end else begin
                    If98948e5f60b2c3ba1d7338e24dc0df6  <=  ~I180deab4fe0d03104cf2ee035f6a9b8c + 1;
                    Iebc1dd048a5c7e83175ba1030a4bb587  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == Iaa19be06695f47ff7d10667289dbde36 ) begin
                    I732bb69d248d700bcfdb287932839da8  <= Iff6cd034bb64d13c21910c11bd92266e;
                    Ie8340c2226ffbab8f79e95ef17594210  <=  0;
                end else begin
                    I732bb69d248d700bcfdb287932839da8  <=  ~Iff6cd034bb64d13c21910c11bd92266e + 1;
                    Ie8340c2226ffbab8f79e95ef17594210  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == I21adefc729265cc5ae67ce279a0a78a2 ) begin
                    I403a8ece76036b3ce6277435609548a5  <= I7c34057a77f2bdda93c422506959818d;
                    Ic7dcd6d9c98422e20947712d0f4adc62  <=  0;
                end else begin
                    I403a8ece76036b3ce6277435609548a5  <=  ~I7c34057a77f2bdda93c422506959818d + 1;
                    Ic7dcd6d9c98422e20947712d0f4adc62  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == Ibc0592b70bd60e475066554f0c7c4171 ) begin
                    I5a6cf1bdbcb2a342e548fb44c171aaf4  <= I7ff7d3fd63fa67cd72d1591c1a373180;
                    I7df25ee69290c62782cd05715b0a6ecb  <=  0;
                end else begin
                    I5a6cf1bdbcb2a342e548fb44c171aaf4  <=  ~I7ff7d3fd63fa67cd72d1591c1a373180 + 1;
                    I7df25ee69290c62782cd05715b0a6ecb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == I14f80574ea80b02ce13079854991febd ) begin
                    I83a16a5be8d92896234bb9f2a36a22c9  <= If910e75bf10cf02a5b414cbb4fad1304;
                    If904894b9cd6236c35bd9de268fab07d  <=  0;
                end else begin
                    I83a16a5be8d92896234bb9f2a36a22c9  <=  ~If910e75bf10cf02a5b414cbb4fad1304 + 1;
                    If904894b9cd6236c35bd9de268fab07d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == I09aae1dd6d02bd2a65dc7fa06fd848ca ) begin
                    I6cad1cb66561eb6f0e3bfe5070b290c2  <= I266697a6eca2b73a76fd375a0ad72a05;
                    I5b890a24c074e7f2ebfee20ce4e15951  <=  0;
                end else begin
                    I6cad1cb66561eb6f0e3bfe5070b290c2  <=  ~I266697a6eca2b73a76fd375a0ad72a05 + 1;
                    I5b890a24c074e7f2ebfee20ce4e15951  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == Idd698fb3a64825b43803642fc91bf674 ) begin
                    Ia50c447d5838d7979b2e19796be6221b  <= Iba188abd7715fcbdad3b1f3d985c6fc3;
                    I22f4468c482ed815d200d72ac2da570a  <=  0;
                end else begin
                    Ia50c447d5838d7979b2e19796be6221b  <=  ~Iba188abd7715fcbdad3b1f3d985c6fc3 + 1;
                    I22f4468c482ed815d200d72ac2da570a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I369ffa98995ba0834f8029ecce705c56 == I73c9bd7e52f6049b733b3a594ad6fae7 ) begin
                    Ief62ab0263b74086ae23a208da23e9c7  <= Ic60c640562e3e45c89a1de78af509b6a;
                    I091ae78d995382a96c68c47a60844a9b  <=  0;
                end else begin
                    Ief62ab0263b74086ae23a208da23e9c7  <=  ~Ic60c640562e3e45c89a1de78af509b6a + 1;
                    I091ae78d995382a96c68c47a60844a9b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == I0fa2b3408156b2b0f656db4947670fe3 ) begin
                    I564999dcc2f67c8f82fb5cd16af0ee12  <= I0456494b33e4ec852c123cb3003b9886;
                    Icbddf0d9df1bad66ea2f7352834bc759  <=  0;
                end else begin
                    I564999dcc2f67c8f82fb5cd16af0ee12  <=  ~I0456494b33e4ec852c123cb3003b9886 + 1;
                    Icbddf0d9df1bad66ea2f7352834bc759  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == Ifd85deef561f76562208a8798b540b99 ) begin
                    Ifb0e4775ffb73bb2533844db969ab900  <= I2ed7c217fe3e21fcb27e04f68b95dd6b;
                    I9a0db2b202a01aad173d2c8109cc596d  <=  0;
                end else begin
                    Ifb0e4775ffb73bb2533844db969ab900  <=  ~I2ed7c217fe3e21fcb27e04f68b95dd6b + 1;
                    I9a0db2b202a01aad173d2c8109cc596d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == I9d6eec32202aeaf66e7815492ac483b2 ) begin
                    Ib109fcaa55c3094cadb0c1f5f40ca752  <= Ifda5780b42bf451a7ce834f17b3fdd20;
                    I724071f9e582e988d8f2d4c98ab9c070  <=  0;
                end else begin
                    Ib109fcaa55c3094cadb0c1f5f40ca752  <=  ~Ifda5780b42bf451a7ce834f17b3fdd20 + 1;
                    I724071f9e582e988d8f2d4c98ab9c070  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == Id771356ebafcbb0e2bb8b03e49148b99 ) begin
                    I56aeb1bd0b0e9857d9cfd2c6b347fe91  <= Iadca92fd39d1fd6032feb8415ca5246f;
                    I31e8ca0bb1f64410501bb3c55bbb60fd  <=  0;
                end else begin
                    I56aeb1bd0b0e9857d9cfd2c6b347fe91  <=  ~Iadca92fd39d1fd6032feb8415ca5246f + 1;
                    I31e8ca0bb1f64410501bb3c55bbb60fd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == I7f4f192560919410f2526392d10776a1 ) begin
                    I02651642fc35059fe9b4141c2fa1f34a  <= I613453382f19dd7eb9bdf51e945a33b0;
                    Ib7b1834c1a9867cb8f42c9ab177dc11c  <=  0;
                end else begin
                    I02651642fc35059fe9b4141c2fa1f34a  <=  ~I613453382f19dd7eb9bdf51e945a33b0 + 1;
                    Ib7b1834c1a9867cb8f42c9ab177dc11c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == I4e2247be1d2dd1af7467039a05447631 ) begin
                    I1f1e04979c8a5badc8a103809f76dadb  <= Ideafa683e6a3a38848fb8bee22eba11b;
                    Iaf22f59aaf7fa5f0e87a8d7504427627  <=  0;
                end else begin
                    I1f1e04979c8a5badc8a103809f76dadb  <=  ~Ideafa683e6a3a38848fb8bee22eba11b + 1;
                    Iaf22f59aaf7fa5f0e87a8d7504427627  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == I5146e2d888c120b7afc430cc8d1dd34c ) begin
                    I19fe22e1104703ddc9bbc94a5368bbc2  <= Ie4226e7e17c7971f07aaf0cfaeae495a;
                    Iea702a29812bf0e4b61cf21351648fe4  <=  0;
                end else begin
                    I19fe22e1104703ddc9bbc94a5368bbc2  <=  ~Ie4226e7e17c7971f07aaf0cfaeae495a + 1;
                    Iea702a29812bf0e4b61cf21351648fe4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == Ib34be78c56c66ff7d85745612cd59f60 ) begin
                    I4386a95203c4fe83c6db7e25a288fc4c  <= Ifbbfa268bd4c31c7eed45cd43fe6a405;
                    I05fa85d0596e05c1df86434a2083c4e1  <=  0;
                end else begin
                    I4386a95203c4fe83c6db7e25a288fc4c  <=  ~Ifbbfa268bd4c31c7eed45cd43fe6a405 + 1;
                    I05fa85d0596e05c1df86434a2083c4e1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == Ic6f48b24e0247c43666af5f25f03c1dc ) begin
                    I2ddabc0b4bc45698fdd877c93bcbe280  <= Ib2d99d95f7a31e4745211c5ff96f851c;
                    Ic61a806c6bc223d2c23cf24dbf3e85db  <=  0;
                end else begin
                    I2ddabc0b4bc45698fdd877c93bcbe280  <=  ~Ib2d99d95f7a31e4745211c5ff96f851c + 1;
                    Ic61a806c6bc223d2c23cf24dbf3e85db  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ccef4c47ae7cfab43584de0f2e193d3 == If9f312c27d80be62969c60eb9b67586c ) begin
                    I5adddbf99d0d39c5d70ec6a0978f3ef5  <= I692c0a91b415b400a3640e2d9a40edad;
                    I8284c12f98671842255420333096213f  <=  0;
                end else begin
                    I5adddbf99d0d39c5d70ec6a0978f3ef5  <=  ~I692c0a91b415b400a3640e2d9a40edad + 1;
                    I8284c12f98671842255420333096213f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ief31fe169c1b360d5933558208dbb602 == Ic7e3298aeb02d5829de1904288687002 ) begin
                    Ia24d776498719aa6cfbdb5df69d648e3  <= If8c4dc70212e8873167e1cad8e8e5692;
                    Ide2e42206ceb5cc9ddd1646dea75776f  <=  0;
                end else begin
                    Ia24d776498719aa6cfbdb5df69d648e3  <=  ~If8c4dc70212e8873167e1cad8e8e5692 + 1;
                    Ide2e42206ceb5cc9ddd1646dea75776f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ief31fe169c1b360d5933558208dbb602 == Ib45f271c90e7bb32cba9dbaad5334c67 ) begin
                    I038ff8eadf1c551dc42d09fbadaea5b9  <= Ib2f75e91bf9e1d32a3f170fc85244139;
                    I47512947d0532033dfa2b015aa107642  <=  0;
                end else begin
                    I038ff8eadf1c551dc42d09fbadaea5b9  <=  ~Ib2f75e91bf9e1d32a3f170fc85244139 + 1;
                    I47512947d0532033dfa2b015aa107642  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ief31fe169c1b360d5933558208dbb602 == I727821089976c74cd540ec58ecce2da2 ) begin
                    I102dc8709a274d21c09abae1d2ac1272  <= I3606dc61f24567cb1ace443cea62a43b;
                    Ia5ec36569a57a6256966da94a52875d1  <=  0;
                end else begin
                    I102dc8709a274d21c09abae1d2ac1272  <=  ~I3606dc61f24567cb1ace443cea62a43b + 1;
                    Ia5ec36569a57a6256966da94a52875d1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ief31fe169c1b360d5933558208dbb602 == I4ed27d0c804891ee239ae8259d200712 ) begin
                    I136256458e71d84e850b61a950f279e7  <= Ie402c9f793b7306323efb8fe23533250;
                    I07ea72a5755bd2b0da6e89389df44f69  <=  0;
                end else begin
                    I136256458e71d84e850b61a950f279e7  <=  ~Ie402c9f793b7306323efb8fe23533250 + 1;
                    I07ea72a5755bd2b0da6e89389df44f69  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ief31fe169c1b360d5933558208dbb602 == I421ad50f600133f1e7f6a52625181d36 ) begin
                    Icda6fe755f2d840f8e404d84b231e827  <= I54652565023310e2eccfc4cb87c56b43;
                    I89b6e7810b2a5d45238819a6a171dac6  <=  0;
                end else begin
                    Icda6fe755f2d840f8e404d84b231e827  <=  ~I54652565023310e2eccfc4cb87c56b43 + 1;
                    I89b6e7810b2a5d45238819a6a171dac6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ief31fe169c1b360d5933558208dbb602 == I172379505892287217e08c060285018b ) begin
                    I1f6cd53f31f27d86d78d5079e84c9716  <= I616b7a5987edbc001e0ae1b638f25a39;
                    I2e6141be9be5edab8e67a1e7f640903f  <=  0;
                end else begin
                    I1f6cd53f31f27d86d78d5079e84c9716  <=  ~I616b7a5987edbc001e0ae1b638f25a39 + 1;
                    I2e6141be9be5edab8e67a1e7f640903f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ief31fe169c1b360d5933558208dbb602 == I8ac36cb7b4e56689efd4a3de1fafa0cc ) begin
                    Ia1f69042d447cb17772b29f634344b53  <= I06604bac478ee906b3fe8ff307cdf046;
                    Ib438d8ef5fdd32b2811e0e755acdfefb  <=  0;
                end else begin
                    Ia1f69042d447cb17772b29f634344b53  <=  ~I06604bac478ee906b3fe8ff307cdf046 + 1;
                    Ib438d8ef5fdd32b2811e0e755acdfefb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ief31fe169c1b360d5933558208dbb602 == I002e83f2fb7e5b07710a802aa505b2bc ) begin
                    I84648f139f0fd470a62f0638aeee9e97  <= I135dd8a85aca863db660f2ad4f80ca2e;
                    I21cc09d0a95b4598c5614b7af3c6fe03  <=  0;
                end else begin
                    I84648f139f0fd470a62f0638aeee9e97  <=  ~I135dd8a85aca863db660f2ad4f80ca2e + 1;
                    I21cc09d0a95b4598c5614b7af3c6fe03  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 == I26fe780ca6becdc9f86a7be04c6257d2 ) begin
                    I6ebc0ad14d76d3a80a4929ba8b5e7848  <= I8715d73b58270dfa33b903e9cfb50be8;
                    Ia7a6617c92f999d7c19d3c338cc60e8f  <=  0;
                end else begin
                    I6ebc0ad14d76d3a80a4929ba8b5e7848  <=  ~I8715d73b58270dfa33b903e9cfb50be8 + 1;
                    Ia7a6617c92f999d7c19d3c338cc60e8f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 == I3a8d18e570ec3aefcdc29d7bc783dfde ) begin
                    I26cba2d4920ff7fc40b1723c29ed8391  <= I7f60cb59895af6d314f5d0f401c80350;
                    I5ea3e9e13e199daf8df53389a405cd0a  <=  0;
                end else begin
                    I26cba2d4920ff7fc40b1723c29ed8391  <=  ~I7f60cb59895af6d314f5d0f401c80350 + 1;
                    I5ea3e9e13e199daf8df53389a405cd0a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 == I4ddf83c90adcc1bec65f265e898568fd ) begin
                    I27980b3a1936a92a1751588f91a5f542  <= I3e25e6e9de5ee9242a472ce957056762;
                    I5a202e3ec847e13fa21134123db7a027  <=  0;
                end else begin
                    I27980b3a1936a92a1751588f91a5f542  <=  ~I3e25e6e9de5ee9242a472ce957056762 + 1;
                    I5a202e3ec847e13fa21134123db7a027  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 == I0c06a37e120e59f19578c68801a4b6ec ) begin
                    I5464cf638e0ca778d4e113b216084180  <= I4c5f36517aaf872e7f05de2f7f76a6ce;
                    Ie697e69bd62cf7bef4a4934843967cec  <=  0;
                end else begin
                    I5464cf638e0ca778d4e113b216084180  <=  ~I4c5f36517aaf872e7f05de2f7f76a6ce + 1;
                    Ie697e69bd62cf7bef4a4934843967cec  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 == Ic290ad8aeb51c16106f9311b06134a2d ) begin
                    I1804dfc05236c728f563342eb011f4f8  <= I0e993e6f98616632f17835a2994f45e3;
                    I6979425ff99d598782f2a45b1d463f8d  <=  0;
                end else begin
                    I1804dfc05236c728f563342eb011f4f8  <=  ~I0e993e6f98616632f17835a2994f45e3 + 1;
                    I6979425ff99d598782f2a45b1d463f8d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 == Ic4c7c898ca601e4d44076ec5bb475979 ) begin
                    Id219264de5f6b67cff866b2bafc660b5  <= I281f996740b16568b9d29ca41a3fa50d;
                    Ie735fb63c3d40f44ede25d0a213847a8  <=  0;
                end else begin
                    Id219264de5f6b67cff866b2bafc660b5  <=  ~I281f996740b16568b9d29ca41a3fa50d + 1;
                    Ie735fb63c3d40f44ede25d0a213847a8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 == I380cd867541300f76fc359d72f49bdbc ) begin
                    I03e4f803d4b82aa774662e02b188b0a6  <= I55bbb73d68871d9dbce4d590c029aeab;
                    I2f132b8b367a5eb3d7029b1c27991dbe  <=  0;
                end else begin
                    I03e4f803d4b82aa774662e02b188b0a6  <=  ~I55bbb73d68871d9dbce4d590c029aeab + 1;
                    I2f132b8b367a5eb3d7029b1c27991dbe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8c0317dafcfb91b3da5eb5afae1f2e2 == I350f20848080cffa45a31e2f1e553a3a ) begin
                    I32e079707d9ce4b31aea8fd2c998c27c  <= Ida491561008f4984480d1b0f09d2fa77;
                    I55291a60dc5b1255d71ab749eaba0404  <=  0;
                end else begin
                    I32e079707d9ce4b31aea8fd2c998c27c  <=  ~Ida491561008f4984480d1b0f09d2fa77 + 1;
                    I55291a60dc5b1255d71ab749eaba0404  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd == I912b9be8432d4eb792d79566a8280703 ) begin
                    I488f60405ded7af04c941bdbf55290f8  <= I624e237f248d292c0417ff85056857b0;
                    I804b17fba020affb1ed32666d73607ae  <=  0;
                end else begin
                    I488f60405ded7af04c941bdbf55290f8  <=  ~I624e237f248d292c0417ff85056857b0 + 1;
                    I804b17fba020affb1ed32666d73607ae  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd == Ifaed59e29ee3ee9166192bbbf04bc682 ) begin
                    I26d314b69785bdb0ca8cd52c258c3b35  <= Ic7c1fd79ba76dbb254c6183017f40b3e;
                    I478f85d129f1f538304e6cc74b9d2234  <=  0;
                end else begin
                    I26d314b69785bdb0ca8cd52c258c3b35  <=  ~Ic7c1fd79ba76dbb254c6183017f40b3e + 1;
                    I478f85d129f1f538304e6cc74b9d2234  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd == I7eaa9f70586b12e371db5964758ee7c2 ) begin
                    Ia490437ab050e63e611dfb4d9366017c  <= I546d683af76dc209a5205c6274abe908;
                    I71ef5d9d9f272131a3c7bf864c0b4863  <=  0;
                end else begin
                    Ia490437ab050e63e611dfb4d9366017c  <=  ~I546d683af76dc209a5205c6274abe908 + 1;
                    I71ef5d9d9f272131a3c7bf864c0b4863  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd == I9a8946bbda4bfe72fab3c2f59533b3ae ) begin
                    Ia6cc50c8b7f83dd80d7058eea40338e9  <= I7b4bb785489c5bb22c84d9778192fe44;
                    I65ed551a24cd36ae20d1ffeac42fb99b  <=  0;
                end else begin
                    Ia6cc50c8b7f83dd80d7058eea40338e9  <=  ~I7b4bb785489c5bb22c84d9778192fe44 + 1;
                    I65ed551a24cd36ae20d1ffeac42fb99b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd == I29fd8dea7c3c39722614210cb7f65851 ) begin
                    I3652208cee3ca6dcdef63b7df53e4329  <= Ifc6af7d7aeb7162d554b8604a44f3361;
                    I4c99cb1e56179799079d9a484edf2a02  <=  0;
                end else begin
                    I3652208cee3ca6dcdef63b7df53e4329  <=  ~Ifc6af7d7aeb7162d554b8604a44f3361 + 1;
                    I4c99cb1e56179799079d9a484edf2a02  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd == I54bed2059ffd24ac2fa91b038c0256ae ) begin
                    Ia9a4760f6a2bf8f8f660e2b0c31dd823  <= I5b650c4c3291670b480a7f1095093dfb;
                    Ibd985ec8f6f4eed7f14ae2692367cc00  <=  0;
                end else begin
                    Ia9a4760f6a2bf8f8f660e2b0c31dd823  <=  ~I5b650c4c3291670b480a7f1095093dfb + 1;
                    Ibd985ec8f6f4eed7f14ae2692367cc00  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd == Ic3608e6a6c45ee04ccd8198c88c69003 ) begin
                    I5ec267a535ad08c629940d70c61894a5  <= I2f5f88cb5e5e4723bd8a83c5fa80cc4c;
                    Ic7eb65782a34589e2b015442172d7568  <=  0;
                end else begin
                    I5ec267a535ad08c629940d70c61894a5  <=  ~I2f5f88cb5e5e4723bd8a83c5fa80cc4c + 1;
                    Ic7eb65782a34589e2b015442172d7568  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I54e3f08f6f4cf784da57ac39f246b8fd == I37da881d3575c055944719409ddb66f1 ) begin
                    I17fadd913ac1008fcbefff48ad366d8f  <= Ic174b361182c98486e65b7f87b073274;
                    I3bb60f8d4ccc5e40e97af6f6718c90c9  <=  0;
                end else begin
                    I17fadd913ac1008fcbefff48ad366d8f  <=  ~Ic174b361182c98486e65b7f87b073274 + 1;
                    I3bb60f8d4ccc5e40e97af6f6718c90c9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I16c7f1b874b0d05c6d120bbede254416 == I2b6999fd13f9e57ea33c0b4602594c66 ) begin
                    I275728fecbd15ba77f57860bb329da16  <= I7ba2f7201745258dbf224de087a25233;
                    Ib109c4220b1113561ec1319a0ac74498  <=  0;
                end else begin
                    I275728fecbd15ba77f57860bb329da16  <=  ~I7ba2f7201745258dbf224de087a25233 + 1;
                    Ib109c4220b1113561ec1319a0ac74498  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I16c7f1b874b0d05c6d120bbede254416 == Idee62819bc831a9ba7c73dea46f3da9a ) begin
                    I8d0bc446761559f2188e78200eb0a895  <= I131a4bd335fc23ee10f7ccb1881ab9cd;
                    I91ec97b5793a453f81b1780157e12d47  <=  0;
                end else begin
                    I8d0bc446761559f2188e78200eb0a895  <=  ~I131a4bd335fc23ee10f7ccb1881ab9cd + 1;
                    I91ec97b5793a453f81b1780157e12d47  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I16c7f1b874b0d05c6d120bbede254416 == I48c95e9ee4d7dd54b6bf21a9a5b20635 ) begin
                    If9fc4683c2f0545e1f077541fd25da66  <= I90cb3e06b42f25956b788a792eef371f;
                    Icae10f8dc7273f91884f011b6a88cf91  <=  0;
                end else begin
                    If9fc4683c2f0545e1f077541fd25da66  <=  ~I90cb3e06b42f25956b788a792eef371f + 1;
                    Icae10f8dc7273f91884f011b6a88cf91  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I16c7f1b874b0d05c6d120bbede254416 == I26b2a20b53a3ef8531d6798c4b272422 ) begin
                    I1c8e7559160d5a1fe1fa0002cc414d1c  <= I56302770a8d56932e7bb5dcff56c71e2;
                    I8b7efa4f096bf761a8df08d1a3f1b77f  <=  0;
                end else begin
                    I1c8e7559160d5a1fe1fa0002cc414d1c  <=  ~I56302770a8d56932e7bb5dcff56c71e2 + 1;
                    I8b7efa4f096bf761a8df08d1a3f1b77f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I16c7f1b874b0d05c6d120bbede254416 == Ib814d21cc76c4f3135a4aa813dcb748d ) begin
                    I059014ede8b9092d817c0aaa1c7ed388  <= Id3b8c058b3838c388eb5ddcb31dfc799;
                    Ib0dfb26e39fd974f64d54a0f9c0cd552  <=  0;
                end else begin
                    I059014ede8b9092d817c0aaa1c7ed388  <=  ~Id3b8c058b3838c388eb5ddcb31dfc799 + 1;
                    Ib0dfb26e39fd974f64d54a0f9c0cd552  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I16c7f1b874b0d05c6d120bbede254416 == I44dcb4df87d1cf32ee2c9bea836223ea ) begin
                    I6294fc2c9181871210e0cfbb9834c3c7  <= I7ca8ce63dfb821d10304958bada71737;
                    Ida3a51bb8109fd4c3e494b736889efaf  <=  0;
                end else begin
                    I6294fc2c9181871210e0cfbb9834c3c7  <=  ~I7ca8ce63dfb821d10304958bada71737 + 1;
                    Ida3a51bb8109fd4c3e494b736889efaf  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I16c7f1b874b0d05c6d120bbede254416 == I96ea91e1bf398f6b2973e815a6a10aaa ) begin
                    Id24dd0ede5504678fbd809ffbacd0dcb  <= I06ad44414b45d262f9542015d2dead8d;
                    I6a47d611882f8af53484f22ce5b74fe6  <=  0;
                end else begin
                    Id24dd0ede5504678fbd809ffbacd0dcb  <=  ~I06ad44414b45d262f9542015d2dead8d + 1;
                    I6a47d611882f8af53484f22ce5b74fe6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I16c7f1b874b0d05c6d120bbede254416 == I75458b8dd7bf267526c36af5cbfcaad1 ) begin
                    I496994e784eb114337ac9e78ec0c4d3f  <= I833ef4acfed17e4699d65cbaa3e7dbd5;
                    I52af26697dd18d51e902642e19045d9a  <=  0;
                end else begin
                    I496994e784eb114337ac9e78ec0c4d3f  <=  ~I833ef4acfed17e4699d65cbaa3e7dbd5 + 1;
                    I52af26697dd18d51e902642e19045d9a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == I230ed2d0ad383ba3a6b5b69ce09ab4b6 ) begin
                    I44c28351f261765c28a066a581c27c13  <= Ia77e3db939408af719e0a8555dcb68ed;
                    I38b0b02379864bed0b097754dac42dec  <=  0;
                end else begin
                    I44c28351f261765c28a066a581c27c13  <=  ~Ia77e3db939408af719e0a8555dcb68ed + 1;
                    I38b0b02379864bed0b097754dac42dec  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == I6c09d773366bca735c15703f7c2c5a11 ) begin
                    I84419e016619a3a33224eeaba85e68b3  <= I57ab4999187992eda55a82bf0f09b31f;
                    Ic3f80e7837ab46f58cfd4b6c775d4e72  <=  0;
                end else begin
                    I84419e016619a3a33224eeaba85e68b3  <=  ~I57ab4999187992eda55a82bf0f09b31f + 1;
                    Ic3f80e7837ab46f58cfd4b6c775d4e72  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == I146e4737d01377560ffeb78fce84973d ) begin
                    I67d114d975d5d65f575bbb8c819fa22b  <= I21f7b5402ae8e8954d99931bd5108250;
                    I87b9dff79eb8389488e97e427d59d767  <=  0;
                end else begin
                    I67d114d975d5d65f575bbb8c819fa22b  <=  ~I21f7b5402ae8e8954d99931bd5108250 + 1;
                    I87b9dff79eb8389488e97e427d59d767  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == Iaa4c0cb6fd4dcc74d6ffd2bde42b7947 ) begin
                    I6a452adc2501774b55e5fe73c642ea26  <= I3627708869b47d460182bc5040092f9a;
                    I44926d094aefc5aa52713fb52704f84f  <=  0;
                end else begin
                    I6a452adc2501774b55e5fe73c642ea26  <=  ~I3627708869b47d460182bc5040092f9a + 1;
                    I44926d094aefc5aa52713fb52704f84f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == I49d021b0957d65a6c2608de826c2676e ) begin
                    I33792929f4428ddf0629231288e459ec  <= Ifd88f0f0abd1c037434dc16e34550d2a;
                    I57127b05215e4faa4e32d5ca38611eb2  <=  0;
                end else begin
                    I33792929f4428ddf0629231288e459ec  <=  ~Ifd88f0f0abd1c037434dc16e34550d2a + 1;
                    I57127b05215e4faa4e32d5ca38611eb2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == I72393e4bfc85c2b9ee24a4395b3568eb ) begin
                    Id0013f18ab77416e08d994c360b13473  <= I27eec53da48406e7e1202345a0810e08;
                    I79aadc384d50af92ae1af6760ffe3b3b  <=  0;
                end else begin
                    Id0013f18ab77416e08d994c360b13473  <=  ~I27eec53da48406e7e1202345a0810e08 + 1;
                    I79aadc384d50af92ae1af6760ffe3b3b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == Ic9f855b66d25668256912f2e434b4854 ) begin
                    I5683f67c7d462c01c55b8be9b6d1fca6  <= I682d42afaaf103550ce4fbdba6192c88;
                    I28effe4aa10b24a221d5e1c84f2c21ff  <=  0;
                end else begin
                    I5683f67c7d462c01c55b8be9b6d1fca6  <=  ~I682d42afaaf103550ce4fbdba6192c88 + 1;
                    I28effe4aa10b24a221d5e1c84f2c21ff  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == I27fe4e83261eb6a1789a8f7d77a0caf1 ) begin
                    I4a5e3cf3066a4c2f7f5f8dbe824ff88f  <= If225534847db8723768941c3819ed7c0;
                    Ia0d7cfa22522e5b4f7b545aacff7fa59  <=  0;
                end else begin
                    I4a5e3cf3066a4c2f7f5f8dbe824ff88f  <=  ~If225534847db8723768941c3819ed7c0 + 1;
                    Ia0d7cfa22522e5b4f7b545aacff7fa59  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == I45c158cf7145668cb8524f7fa06f9302 ) begin
                    I93879adfa4333a80be696d846e34d799  <= I43a91b2232a47d1f6731bafc15ced5db;
                    Ifdac0b0a75dfcc09291fd95e842e68f1  <=  0;
                end else begin
                    I93879adfa4333a80be696d846e34d799  <=  ~I43a91b2232a47d1f6731bafc15ced5db + 1;
                    Ifdac0b0a75dfcc09291fd95e842e68f1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c3cb2de514ecab0dd311e86a4dc3cdb == I16d2a9270452f0d8b6eda06ea939fc6a ) begin
                    I199e944b303446e2cdafb6f34d0d12c7  <= Ic54026604afd19b0c7c71ea1ac0f1c4e;
                    I1bbd0d48cc6bd8a4d4d520d38798f74c  <=  0;
                end else begin
                    I199e944b303446e2cdafb6f34d0d12c7  <=  ~Ic54026604afd19b0c7c71ea1ac0f1c4e + 1;
                    I1bbd0d48cc6bd8a4d4d520d38798f74c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == I1ab974ad9718ea8350d76bbc1510d2d1 ) begin
                    I91d282de42df72b1c439fede384d6336  <= I218bd69f079aa21f0dda241ae6e387ad;
                    I06ede5ab6bc97827c4f866dca1aa17bc  <=  0;
                end else begin
                    I91d282de42df72b1c439fede384d6336  <=  ~I218bd69f079aa21f0dda241ae6e387ad + 1;
                    I06ede5ab6bc97827c4f866dca1aa17bc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == I31467f39d6b5c20d4e155d19afa34e95 ) begin
                    I8a06d2c278af9d552fa36a61128b8a9b  <= Iaaacca4d06ad0f202d839fd7674f1829;
                    I4b7f22e0b9e1589fbc1d558b37cceb37  <=  0;
                end else begin
                    I8a06d2c278af9d552fa36a61128b8a9b  <=  ~Iaaacca4d06ad0f202d839fd7674f1829 + 1;
                    I4b7f22e0b9e1589fbc1d558b37cceb37  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == Ia8762fb956b52535ad6921e9191288d0 ) begin
                    I5a36e45af7599ec00703dfc81f9d1176  <= Iecddac410bb2121da0df2d73c2d23cb8;
                    I6e63e4047456268e73ad16a5cde93681  <=  0;
                end else begin
                    I5a36e45af7599ec00703dfc81f9d1176  <=  ~Iecddac410bb2121da0df2d73c2d23cb8 + 1;
                    I6e63e4047456268e73ad16a5cde93681  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == Ia018c4c165c5af9a329a63aa365ac038 ) begin
                    Iae09429ca8733186fdb3c50f36895746  <= I1aabc0c0b7b602297ad592ae48b23452;
                    Iec7997b0018f4fb3572579a5bf1e4728  <=  0;
                end else begin
                    Iae09429ca8733186fdb3c50f36895746  <=  ~I1aabc0c0b7b602297ad592ae48b23452 + 1;
                    Iec7997b0018f4fb3572579a5bf1e4728  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == Id85085de57a0152aad8cf5e27a195052 ) begin
                    Ie5f74b33d06ddb8b32b57c8c82392001  <= Ida3aaf7237b1383cfe95eeccf3971a8e;
                    I11cb6032d99f05b3f908418a70fd3d6e  <=  0;
                end else begin
                    Ie5f74b33d06ddb8b32b57c8c82392001  <=  ~Ida3aaf7237b1383cfe95eeccf3971a8e + 1;
                    I11cb6032d99f05b3f908418a70fd3d6e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == I461b443279e5bf47de450846e3da7d8e ) begin
                    I7d3cdb71cdab3a85122130207d872476  <= Idd2a8ed39edf6697b0988ee4eb4f2d95;
                    Idba56a073e34e530c36025914f7646d9  <=  0;
                end else begin
                    I7d3cdb71cdab3a85122130207d872476  <=  ~Idd2a8ed39edf6697b0988ee4eb4f2d95 + 1;
                    Idba56a073e34e530c36025914f7646d9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == I71d07a22b66aed8c24fe4dd203869fa1 ) begin
                    I68ae9f2a14b161c940f6685073eca97e  <= I735c660d5232e03dd8fb129e2ca4b445;
                    I3a7582a1c86f2b49979372132ce98c87  <=  0;
                end else begin
                    I68ae9f2a14b161c940f6685073eca97e  <=  ~I735c660d5232e03dd8fb129e2ca4b445 + 1;
                    I3a7582a1c86f2b49979372132ce98c87  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == I173b85306dc75e596cfe67f7c518f36b ) begin
                    I778f907b5eacdfac02b0bc4547af4ea3  <= Ia04d6065987df3f007658614406cbc28;
                    Ifaed912ee00082f8458ae37bd47179a5  <=  0;
                end else begin
                    I778f907b5eacdfac02b0bc4547af4ea3  <=  ~Ia04d6065987df3f007658614406cbc28 + 1;
                    Ifaed912ee00082f8458ae37bd47179a5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == Id57948138d3091aa350db0d906b06b34 ) begin
                    Ibcea5bf1e21fa764ac9f2d2702c8f79a  <= I7aeddde5b60828ac7f8b6c2addaf220b;
                    Ibecc30f33083404bf48eb0005e14bb83  <=  0;
                end else begin
                    Ibcea5bf1e21fa764ac9f2d2702c8f79a  <=  ~I7aeddde5b60828ac7f8b6c2addaf220b + 1;
                    Ibecc30f33083404bf48eb0005e14bb83  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icc5ba4554d7a44bc3b43377efbe3b5f8 == If6b37dd338e28ffd7fb888bc56f716d1 ) begin
                    I93a3e1a8e414d4775f19c0c9f16d07a8  <= I150c28296847348d69cce123f20656c3;
                    I87009d289b53c6e366b73e275e414caf  <=  0;
                end else begin
                    I93a3e1a8e414d4775f19c0c9f16d07a8  <=  ~I150c28296847348d69cce123f20656c3 + 1;
                    I87009d289b53c6e366b73e275e414caf  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == Idd412a66c4a434eaaf337b6b4ab6b0a5 ) begin
                    I8772034840834e51187950d320f9eb40  <= Ib94d38d19b3791fa2d1b42fdfde8435e;
                    I5d5b08cc3fd13b96621143655a806c7d  <=  0;
                end else begin
                    I8772034840834e51187950d320f9eb40  <=  ~Ib94d38d19b3791fa2d1b42fdfde8435e + 1;
                    I5d5b08cc3fd13b96621143655a806c7d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == I5829341b8f12f906ffc53c9d716e6556 ) begin
                    I3d0aa00b61d4684ad46f49329197c901  <= I94865622898b2e481e86a244f7aa2759;
                    I94ce074b29f44c5e4a63ff6e00d2b9c4  <=  0;
                end else begin
                    I3d0aa00b61d4684ad46f49329197c901  <=  ~I94865622898b2e481e86a244f7aa2759 + 1;
                    I94ce074b29f44c5e4a63ff6e00d2b9c4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == I449b6fdea575e92fa4603f141ff359e8 ) begin
                    I146866a6d46604c47d87afa3c88308c6  <= I1a4a432e735367f515ca747cef7d7d04;
                    I2fd3e923d1adff22ef7718dae5632b29  <=  0;
                end else begin
                    I146866a6d46604c47d87afa3c88308c6  <=  ~I1a4a432e735367f515ca747cef7d7d04 + 1;
                    I2fd3e923d1adff22ef7718dae5632b29  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == Ic6581fe8d97a45b71a1ca8d9ec97f97b ) begin
                    I84cf7aa78617faed2f1762bb1961cc0e  <= Ib3a2b744d8f38671a63da6f8f8f1a6a1;
                    Ibe2d184a52eb5d33cac0ca4a5dab55f6  <=  0;
                end else begin
                    I84cf7aa78617faed2f1762bb1961cc0e  <=  ~Ib3a2b744d8f38671a63da6f8f8f1a6a1 + 1;
                    Ibe2d184a52eb5d33cac0ca4a5dab55f6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == I4af6879c6d4d2b96562b1c2ada8f92b0 ) begin
                    Ib1f43a0b9c86d236b2ed71c35c296b9c  <= I87716ad5a64592abb812ffe041ccc163;
                    I0907dde542619e162f45f3dac8c0c16f  <=  0;
                end else begin
                    Ib1f43a0b9c86d236b2ed71c35c296b9c  <=  ~I87716ad5a64592abb812ffe041ccc163 + 1;
                    I0907dde542619e162f45f3dac8c0c16f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == I7a176a15ab2c5396639be387bc43896c ) begin
                    I88aaa7538f9007ce204319ec639d1c7e  <= I71b259faefbea7ce8f47e0ffb556a0be;
                    I9bdfa0d38ed6d215e7ef7ecb12185b60  <=  0;
                end else begin
                    I88aaa7538f9007ce204319ec639d1c7e  <=  ~I71b259faefbea7ce8f47e0ffb556a0be + 1;
                    I9bdfa0d38ed6d215e7ef7ecb12185b60  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == I38c29f53b042f039a908cca7d09cc2bf ) begin
                    Ie3a171564602e9936d7960e83bb0fb3a  <= I2161b2ff3514dbdbb79d25da87eeec2b;
                    Ie0e096809efa587a070562473e9a2fff  <=  0;
                end else begin
                    Ie3a171564602e9936d7960e83bb0fb3a  <=  ~I2161b2ff3514dbdbb79d25da87eeec2b + 1;
                    Ie0e096809efa587a070562473e9a2fff  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == I1e5c60072bcfdc56b1928040edf9ecb2 ) begin
                    I732b452fd9521b3a13ff1f965c443325  <= I860a3c9fca8d240c68ce3825192353b0;
                    I8c2c0b7861868365bc3935ef8d0fe309  <=  0;
                end else begin
                    I732b452fd9521b3a13ff1f965c443325  <=  ~I860a3c9fca8d240c68ce3825192353b0 + 1;
                    I8c2c0b7861868365bc3935ef8d0fe309  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == I03998667df412d12539d57112b6b6f76 ) begin
                    I16cd75fd747b600e90763d8ce9c08210  <= Ie4eb18c7e906c9a25c12e9980a9f61cb;
                    Idde6e2f615f8ec0aa66b7397e5581651  <=  0;
                end else begin
                    I16cd75fd747b600e90763d8ce9c08210  <=  ~Ie4eb18c7e906c9a25c12e9980a9f61cb + 1;
                    Idde6e2f615f8ec0aa66b7397e5581651  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5e51f49adb6dce65a9f19ff736526c4b == I2ae5c6ae2de0db31a656018e19d086b9 ) begin
                    Ic6a7d6bfb12f40ae8823db716cfe017a  <= I20a24846a74af76fa4470d6350546a9a;
                    I3098e45c14ec08213883f7879c30150c  <=  0;
                end else begin
                    Ic6a7d6bfb12f40ae8823db716cfe017a  <=  ~I20a24846a74af76fa4470d6350546a9a + 1;
                    I3098e45c14ec08213883f7879c30150c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == I1e27f59e10400144106861daca51e721 ) begin
                    Iea38a3c260d0caae4ae042264a0f4787  <= I90d40f6e9721a7d075512b8b81907453;
                    Ide3c2fa1d5da990a0566c65a12d1d7da  <=  0;
                end else begin
                    Iea38a3c260d0caae4ae042264a0f4787  <=  ~I90d40f6e9721a7d075512b8b81907453 + 1;
                    Ide3c2fa1d5da990a0566c65a12d1d7da  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == Iba8577f8233fe013584171e588868e69 ) begin
                    Id6240152bd22a9655b18bdfd91812e03  <= Ifc4525a25f38affb399004b057d1318c;
                    I6ece8c59f986da73f00e104ff5966189  <=  0;
                end else begin
                    Id6240152bd22a9655b18bdfd91812e03  <=  ~Ifc4525a25f38affb399004b057d1318c + 1;
                    I6ece8c59f986da73f00e104ff5966189  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == I1d0a95c7cced8ede694d02936af63047 ) begin
                    I07eeb34c9dfb9baadb9f263b6f095ecc  <= Icc93649a2050b9ded1e625be936b411f;
                    I5c002c1ec0c63a2c04ca2711fde50254  <=  0;
                end else begin
                    I07eeb34c9dfb9baadb9f263b6f095ecc  <=  ~Icc93649a2050b9ded1e625be936b411f + 1;
                    I5c002c1ec0c63a2c04ca2711fde50254  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == I8b072ed41d990e6afa6fb5d22990f4df ) begin
                    Iedb57db3cbaca9f9a469d91ed81466a8  <= Ibcc30c960ae0f29c4efb1266c9e490ac;
                    Icb5a521ae9f45d8c9101fdde8925e64f  <=  0;
                end else begin
                    Iedb57db3cbaca9f9a469d91ed81466a8  <=  ~Ibcc30c960ae0f29c4efb1266c9e490ac + 1;
                    Icb5a521ae9f45d8c9101fdde8925e64f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == Iab0f19858a1a01fe09fa3c99d92a79fb ) begin
                    I2972b771a4e99ddfa2178349a805b16f  <= I3b2ffa79fd2227a24c6468a89f2bd989;
                    I7b72bfdf546647380e6b1f9a810fd1d1  <=  0;
                end else begin
                    I2972b771a4e99ddfa2178349a805b16f  <=  ~I3b2ffa79fd2227a24c6468a89f2bd989 + 1;
                    I7b72bfdf546647380e6b1f9a810fd1d1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == Id88441b410f55c15465eff4cfa216691 ) begin
                    I6a61cdadaf987763080e6ce4d1605ee6  <= Ib489a11dfdd8a2b3ad561c965b3d7d2a;
                    I84581a99221f2aab1e7cbbcc80296ad4  <=  0;
                end else begin
                    I6a61cdadaf987763080e6ce4d1605ee6  <=  ~Ib489a11dfdd8a2b3ad561c965b3d7d2a + 1;
                    I84581a99221f2aab1e7cbbcc80296ad4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == I894540936535dd20ff1ea5c47546e5fe ) begin
                    I12e430f1ccaa6099ba9ff803c85d9532  <= Ifa51cf9f9d3d1b91c72387f5daf05c79;
                    I27d48bcfb04bf11d76b496d459ee1b48  <=  0;
                end else begin
                    I12e430f1ccaa6099ba9ff803c85d9532  <=  ~Ifa51cf9f9d3d1b91c72387f5daf05c79 + 1;
                    I27d48bcfb04bf11d76b496d459ee1b48  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == Ibb40a1e09cc59e00ce8ba1460e0712d4 ) begin
                    I2cc3c84149c81572357c01219248aa3b  <= Ifda20d77c574c8f13816620c56fff950;
                    Ib89fb8b901f12120ab0bdff5207c74f0  <=  0;
                end else begin
                    I2cc3c84149c81572357c01219248aa3b  <=  ~Ifda20d77c574c8f13816620c56fff950 + 1;
                    Ib89fb8b901f12120ab0bdff5207c74f0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == I5349c1efb5233e8cc6c472ecae80ccc3 ) begin
                    I6d4b18dbba5c2b058f93a8d46bed38ec  <= I03ce0915d3a170429959221b6c8cd16c;
                    Ic2324007897bedbb70a77faa1fd301ef  <=  0;
                end else begin
                    I6d4b18dbba5c2b058f93a8d46bed38ec  <=  ~I03ce0915d3a170429959221b6c8cd16c + 1;
                    Ic2324007897bedbb70a77faa1fd301ef  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id57092394c7cda397f42374df4aa3fec == Id90c5bcfdae1c4abdfa194477917dfbb ) begin
                    I32ca5d01c39fe736d6ed57d70fcbd555  <= I9c2da511df8277b7e61cf8611d04dd32;
                    Ic75af8091015d4615d0c059ceb16371b  <=  0;
                end else begin
                    I32ca5d01c39fe736d6ed57d70fcbd555  <=  ~I9c2da511df8277b7e61cf8611d04dd32 + 1;
                    Ic75af8091015d4615d0c059ceb16371b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idd6a4f8ae94c431f2fa3312b4fd287ba == I1dafa9e7b2a353dee90a0b0f9685a826 ) begin
                    I8807f2f633d64cb064fbc149ebd30412  <= Ib8c628f3d97ffdf8a8b5db0fe90bbfa8;
                    I5b98fb653fa4d3d4ce2ebccd24085f95  <=  0;
                end else begin
                    I8807f2f633d64cb064fbc149ebd30412  <=  ~Ib8c628f3d97ffdf8a8b5db0fe90bbfa8 + 1;
                    I5b98fb653fa4d3d4ce2ebccd24085f95  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idd6a4f8ae94c431f2fa3312b4fd287ba == Ia75e6368415ff53bdbfe81ac2bdfb290 ) begin
                    I822d3b3516499e58ee7777b99259a206  <= I42e0e42ae26723497a1da5e86e855499;
                    Ic9320f9ad332f511422f5b805de9488a  <=  0;
                end else begin
                    I822d3b3516499e58ee7777b99259a206  <=  ~I42e0e42ae26723497a1da5e86e855499 + 1;
                    Ic9320f9ad332f511422f5b805de9488a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idd6a4f8ae94c431f2fa3312b4fd287ba == I91217ca822fb03fdad03b8d005edadc9 ) begin
                    Ie706bf8dd49322fc1d5d83e40fb20f04  <= Id7e44a94fcaa2ca22ac9eb6756ecb830;
                    I71574a4f01fc2e2fdd051a90b9115524  <=  0;
                end else begin
                    Ie706bf8dd49322fc1d5d83e40fb20f04  <=  ~Id7e44a94fcaa2ca22ac9eb6756ecb830 + 1;
                    I71574a4f01fc2e2fdd051a90b9115524  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idd6a4f8ae94c431f2fa3312b4fd287ba == Iccc6e66d1f26c4a5874ba02980dad6a7 ) begin
                    I9975f2ca851119d7ec85cfdefda150f0  <= Ie91db5e628b828dfaa8c1bd7d614d986;
                    Ia59c01c2e6f19ee93a091dbd1a1da83c  <=  0;
                end else begin
                    I9975f2ca851119d7ec85cfdefda150f0  <=  ~Ie91db5e628b828dfaa8c1bd7d614d986 + 1;
                    Ia59c01c2e6f19ee93a091dbd1a1da83c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9f1f8590dcf596097bc81001d51684b9 == I15e9479f1c9aae3c1f12f0f301ee275b ) begin
                    I2e0639bf4e48a7b1486beebcc9ad7c0c  <= I683ebfd7677d9e175d7a86479a5b42c6;
                    I5e8e70c7ad583c0c4f09cacb60602c00  <=  0;
                end else begin
                    I2e0639bf4e48a7b1486beebcc9ad7c0c  <=  ~I683ebfd7677d9e175d7a86479a5b42c6 + 1;
                    I5e8e70c7ad583c0c4f09cacb60602c00  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9f1f8590dcf596097bc81001d51684b9 == I14692ccb24148a020dda28c6f61e3611 ) begin
                    I6131789039de7dc431c3b9b59ecb7654  <= I11090ba16ce17a70438618b474837c33;
                    Ia180d785ba74d63500c25e3a04d21c03  <=  0;
                end else begin
                    I6131789039de7dc431c3b9b59ecb7654  <=  ~I11090ba16ce17a70438618b474837c33 + 1;
                    Ia180d785ba74d63500c25e3a04d21c03  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9f1f8590dcf596097bc81001d51684b9 == Id237c89ded30e926343fb68d786a76d0 ) begin
                    Ia20482fd064712397fe2f9f77f4d854b  <= I845dd61995152e9d39cea7f0370b5a4d;
                    I4dbcb057b2076d4efd4e05e818d976c9  <=  0;
                end else begin
                    Ia20482fd064712397fe2f9f77f4d854b  <=  ~I845dd61995152e9d39cea7f0370b5a4d + 1;
                    I4dbcb057b2076d4efd4e05e818d976c9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9f1f8590dcf596097bc81001d51684b9 == Ib56bd244f7a9876fab3d51a21ef163c7 ) begin
                    If052875ec5a78a68428a1ff09df623df  <= Ia3e4dff8c98b38b6aebec9094ed26421;
                    I24e240c3d018053712e0fb7f861acad7  <=  0;
                end else begin
                    If052875ec5a78a68428a1ff09df623df  <=  ~Ia3e4dff8c98b38b6aebec9094ed26421 + 1;
                    I24e240c3d018053712e0fb7f861acad7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icecd765baa87877675b0f3972d78c02f == Ic1db9806badd4e959a0f0a769e15b6c0 ) begin
                    I2e27abc9297a3fa647f50859af7cb094  <= Id69a54dc4854348a482f052c64a736ca;
                    I78d4209646fe0f2b8027988024b947ae  <=  0;
                end else begin
                    I2e27abc9297a3fa647f50859af7cb094  <=  ~Id69a54dc4854348a482f052c64a736ca + 1;
                    I78d4209646fe0f2b8027988024b947ae  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icecd765baa87877675b0f3972d78c02f == I3649823bb60a4740b6a7f94dd26e45a1 ) begin
                    I5d5e3b64ed1ca16d65d8eadb8100fa06  <= I0f56c52253603ac01a22f3b942429262;
                    I62fa50cc71ade42b52be1de668da6b7b  <=  0;
                end else begin
                    I5d5e3b64ed1ca16d65d8eadb8100fa06  <=  ~I0f56c52253603ac01a22f3b942429262 + 1;
                    I62fa50cc71ade42b52be1de668da6b7b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icecd765baa87877675b0f3972d78c02f == I8d7596d25b93595ffa1ef7d273c98c14 ) begin
                    Ie91a08b49b9bf23270dd3fa331e64968  <= I718f82404f82fe0e822ee20d33ad20a2;
                    I5145e1005293c49c849599347a4a2b46  <=  0;
                end else begin
                    Ie91a08b49b9bf23270dd3fa331e64968  <=  ~I718f82404f82fe0e822ee20d33ad20a2 + 1;
                    I5145e1005293c49c849599347a4a2b46  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icecd765baa87877675b0f3972d78c02f == If607fe1cc3901fc74590a81a26ccb4a8 ) begin
                    Ib599712a1e8fadbdf7e3712bca6c0b74  <= I6c86073aaa32b64a43d06eb1a2d9fba8;
                    Id77a6df77f3d714b6b1f60bad2462f2b  <=  0;
                end else begin
                    Ib599712a1e8fadbdf7e3712bca6c0b74  <=  ~I6c86073aaa32b64a43d06eb1a2d9fba8 + 1;
                    Id77a6df77f3d714b6b1f60bad2462f2b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I401a38ea1d71dcc71d17a4694ceb0988 == Ibe2cd0729747659786b76f044f3caa6e ) begin
                    I1791c009b0838ef10233015f80a5c4af  <= Ie0c8e27167e6ba97a83dd238086f45e6;
                    I6cbfcd474a5a76538db10b8c3235986b  <=  0;
                end else begin
                    I1791c009b0838ef10233015f80a5c4af  <=  ~Ie0c8e27167e6ba97a83dd238086f45e6 + 1;
                    I6cbfcd474a5a76538db10b8c3235986b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I401a38ea1d71dcc71d17a4694ceb0988 == I38e96074261512c31ebd15c6de4b440b ) begin
                    I3dead2d8d18ea8503a578469625f3aa3  <= I6bb5e8ee16a2bc0c3b77c882cfb659e7;
                    I17c80f6af6d201a1214d251778a9e534  <=  0;
                end else begin
                    I3dead2d8d18ea8503a578469625f3aa3  <=  ~I6bb5e8ee16a2bc0c3b77c882cfb659e7 + 1;
                    I17c80f6af6d201a1214d251778a9e534  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I401a38ea1d71dcc71d17a4694ceb0988 == Ie72e9c0aa298ff1809a47908ff86b6c4 ) begin
                    I2fc47140b9df2544d7ae9c82cd38ebd6  <= Ieef625ad664ddadc849be46d1c083748;
                    I468342d7ba88b0a9313f38d0ec2a81e5  <=  0;
                end else begin
                    I2fc47140b9df2544d7ae9c82cd38ebd6  <=  ~Ieef625ad664ddadc849be46d1c083748 + 1;
                    I468342d7ba88b0a9313f38d0ec2a81e5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I401a38ea1d71dcc71d17a4694ceb0988 == Id6e349e3f114f328958052a680a95411 ) begin
                    Ice09150d69c67cd2d08d6e63b8a9bbc7  <= Ice91b069200a91b2ad48fbf87bb2e766;
                    I189be0be892f48991d69acf5a0d42533  <=  0;
                end else begin
                    Ice09150d69c67cd2d08d6e63b8a9bbc7  <=  ~Ice91b069200a91b2ad48fbf87bb2e766 + 1;
                    I189be0be892f48991d69acf5a0d42533  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e == I6dff6c5c76c92ba9626512b35a573ac8 ) begin
                    Id67765c4a6b11f6ee0a4524ebb2d1ca7  <= I9d4c7c85b4da5f7003ff05ed3a240a2e;
                    Ib5bdc1c490d7d2fd11359fc6c79372cb  <=  0;
                end else begin
                    Id67765c4a6b11f6ee0a4524ebb2d1ca7  <=  ~I9d4c7c85b4da5f7003ff05ed3a240a2e + 1;
                    Ib5bdc1c490d7d2fd11359fc6c79372cb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e == I5145ca1a0b7eb68adb93316264ed0084 ) begin
                    Ia17bbf4b7f063de0bf0701276b7b0c20  <= Ia8f1616f8a65025446a5ab4cc1624f9b;
                    I85e112a43fa9046e94da6bdb7b3a13d7  <=  0;
                end else begin
                    Ia17bbf4b7f063de0bf0701276b7b0c20  <=  ~Ia8f1616f8a65025446a5ab4cc1624f9b + 1;
                    I85e112a43fa9046e94da6bdb7b3a13d7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e == Icff67cd5e9472e77380eb812deb625b6 ) begin
                    I9f9075a7745d475331f0b25bad830421  <= I29848deb21ad480cdf155d849dc7bd48;
                    I03ad487e845cce369a813b0c7f32e59d  <=  0;
                end else begin
                    I9f9075a7745d475331f0b25bad830421  <=  ~I29848deb21ad480cdf155d849dc7bd48 + 1;
                    I03ad487e845cce369a813b0c7f32e59d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e == I88adcddd217c9b2363fe254b0be469e2 ) begin
                    I4d832ef88af4d4244516b0bdfd2b461c  <= I1ae69988f89b200bd0e48f640211321c;
                    I85aeb073e949fc999464ce61479790db  <=  0;
                end else begin
                    I4d832ef88af4d4244516b0bdfd2b461c  <=  ~I1ae69988f89b200bd0e48f640211321c + 1;
                    I85aeb073e949fc999464ce61479790db  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e == If149258ed84a848bc38011bef172b6ea ) begin
                    Ib2038174dd555b1d058778fa904aee65  <= I7ddcc3c9f4d21aacc07d8eb285dee83e;
                    I7534524f9d9c64bdf0bb88ba351b3ca5  <=  0;
                end else begin
                    Ib2038174dd555b1d058778fa904aee65  <=  ~I7ddcc3c9f4d21aacc07d8eb285dee83e + 1;
                    I7534524f9d9c64bdf0bb88ba351b3ca5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3db9b61e28a51e974e2d5e323ad53c1e == Ie70f8bcc335351e60eecd70b90d4432c ) begin
                    I959dff5d57b4c2adb85c3602d5874c90  <= I28f7cf50ea7ac81667ff1353e0e121bd;
                    Ic4a902801adb86fdb2481f5b868daa8b  <=  0;
                end else begin
                    I959dff5d57b4c2adb85c3602d5874c90  <=  ~I28f7cf50ea7ac81667ff1353e0e121bd + 1;
                    Ic4a902801adb86fdb2481f5b868daa8b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96d0a4387f9b959bc779ac13351182cc == I5277100478097db96b41fe0988046442 ) begin
                    I30dd112c5a6793cf37bfaaf8dfdebcaf  <= I09b7dd699ae0c4d34a7d1588efc90452;
                    I1141271b2c1fa529b7f4e4ce9ac10c95  <=  0;
                end else begin
                    I30dd112c5a6793cf37bfaaf8dfdebcaf  <=  ~I09b7dd699ae0c4d34a7d1588efc90452 + 1;
                    I1141271b2c1fa529b7f4e4ce9ac10c95  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96d0a4387f9b959bc779ac13351182cc == I0aced2534542d8d2c488c7082ca214ca ) begin
                    I4d4a0930420b4d7da8b6e91b2b25bc51  <= Ic937101cc53e67403e56ac85011aa9ba;
                    Ie62709fd754ca31b0e5d830901bd6433  <=  0;
                end else begin
                    I4d4a0930420b4d7da8b6e91b2b25bc51  <=  ~Ic937101cc53e67403e56ac85011aa9ba + 1;
                    Ie62709fd754ca31b0e5d830901bd6433  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96d0a4387f9b959bc779ac13351182cc == Ifad6157e5199a5b5dbd2465f4cae5b3a ) begin
                    I7ae1d318fd0df386e0c8bcf0f0a94e4b  <= Ib42b03d2f76b8939ff3183008b17a969;
                    I6c6a99a66fe46ca1532fa898123a6131  <=  0;
                end else begin
                    I7ae1d318fd0df386e0c8bcf0f0a94e4b  <=  ~Ib42b03d2f76b8939ff3183008b17a969 + 1;
                    I6c6a99a66fe46ca1532fa898123a6131  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96d0a4387f9b959bc779ac13351182cc == I2bf55a177a00da61ccd463a450de2bb0 ) begin
                    I06cc62e12d5a261d672b5428dbc9767b  <= I4b99f00b1c2cdcee6bf4f1d2e8199ee4;
                    I963a6698cd1f83ce4e7ecaff7f53ce25  <=  0;
                end else begin
                    I06cc62e12d5a261d672b5428dbc9767b  <=  ~I4b99f00b1c2cdcee6bf4f1d2e8199ee4 + 1;
                    I963a6698cd1f83ce4e7ecaff7f53ce25  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96d0a4387f9b959bc779ac13351182cc == I521e3e69d81a6034183d2ba861ec7726 ) begin
                    I9798b16b4658501d739d46182d7ab169  <= I01e153b020e1349eb66b47de581408df;
                    I451d9f14e13b272ea041178627ef7f56  <=  0;
                end else begin
                    I9798b16b4658501d739d46182d7ab169  <=  ~I01e153b020e1349eb66b47de581408df + 1;
                    I451d9f14e13b272ea041178627ef7f56  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96d0a4387f9b959bc779ac13351182cc == Ife32264cdbf7445987f5f39d6361d1e4 ) begin
                    I90bc85b7a6e56250bf13407ddd32bf11  <= I8ca1a48206ed8f1dc7ca57d77d0331a2;
                    I3e7f571589d773eaf3435c03bd13c9ca  <=  0;
                end else begin
                    I90bc85b7a6e56250bf13407ddd32bf11  <=  ~I8ca1a48206ed8f1dc7ca57d77d0331a2 + 1;
                    I3e7f571589d773eaf3435c03bd13c9ca  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 == Ied102cd26c4fc50aa354b16a35d3490b ) begin
                    I88990d32bd34da606660f1c078b36ce0  <= I40e8430f50206db37e500c22f461b0c7;
                    Ie823a06acbb6935875c5cb9088389b27  <=  0;
                end else begin
                    I88990d32bd34da606660f1c078b36ce0  <=  ~I40e8430f50206db37e500c22f461b0c7 + 1;
                    Ie823a06acbb6935875c5cb9088389b27  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 == I5900a9bf6a83b1965f0dd9749d90e317 ) begin
                    Ib32ce57f2840a45fce8e66f71b37719d  <= I521128b7d945e025ded04037494c850a;
                    Ia4c876fe77f09258fb130d03b8cdc67b  <=  0;
                end else begin
                    Ib32ce57f2840a45fce8e66f71b37719d  <=  ~I521128b7d945e025ded04037494c850a + 1;
                    Ia4c876fe77f09258fb130d03b8cdc67b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 == I1b4d2bc08a78865fb281a44e84088fa5 ) begin
                    Ib0179c2048d6c9d1865d171b48c521ff  <= Ic24dbb1a30bb9a32c1992afcba90d4fb;
                    Ie6bf8e5060074ce2dfcf7ddcbb158bff  <=  0;
                end else begin
                    Ib0179c2048d6c9d1865d171b48c521ff  <=  ~Ic24dbb1a30bb9a32c1992afcba90d4fb + 1;
                    Ie6bf8e5060074ce2dfcf7ddcbb158bff  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 == I70724327149d97d4d4f3f71a1500427e ) begin
                    Icc8ffcc0641f0f9405590338e6b5e517  <= I06cc903106b42e397fa7c4bc6c5edea4;
                    I706ad22942f1cfbfae4fde958450189b  <=  0;
                end else begin
                    Icc8ffcc0641f0f9405590338e6b5e517  <=  ~I06cc903106b42e397fa7c4bc6c5edea4 + 1;
                    I706ad22942f1cfbfae4fde958450189b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 == If91997f00102c66a7630ffb2d041d949 ) begin
                    I5d6cb688ef094e1f119d8536f0f56766  <= I765dff22de01d419a6626919d23850f2;
                    Ic64d1cde239aef0df4f227a64762f9f2  <=  0;
                end else begin
                    I5d6cb688ef094e1f119d8536f0f56766  <=  ~I765dff22de01d419a6626919d23850f2 + 1;
                    Ic64d1cde239aef0df4f227a64762f9f2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64082bc75fdbeb69a52a4361ed2d5883 == I25da82603d45fc12f685407e8dc2f6f1 ) begin
                    Ia5aa7c66d2818982a661e4d048876d1c  <= Ie9538b63a057a50371de2d17898d3ad7;
                    I719f60bd29522fded995c8230b4f3a34  <=  0;
                end else begin
                    Ia5aa7c66d2818982a661e4d048876d1c  <=  ~Ie9538b63a057a50371de2d17898d3ad7 + 1;
                    I719f60bd29522fded995c8230b4f3a34  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I62929057b7c214bd38fd532e20ba5623 == Id2fdc5b6c996c567743aaf021a5e6371 ) begin
                    I449e514b6afb3e8e337691fc64f7431c  <= If93a5596528db9017b8783fa0cf1dbc2;
                    I1bd8505e6f316488bb1cdd74932c0314  <=  0;
                end else begin
                    I449e514b6afb3e8e337691fc64f7431c  <=  ~If93a5596528db9017b8783fa0cf1dbc2 + 1;
                    I1bd8505e6f316488bb1cdd74932c0314  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I62929057b7c214bd38fd532e20ba5623 == I8d57ad30940b8351a829b8ca99921a10 ) begin
                    Ibbd5f0906646560a903abcf6848ee80e  <= I68016caaf170fbe2734c5b6aaf089894;
                    I63e645f447ddd1fc9409879872479bef  <=  0;
                end else begin
                    Ibbd5f0906646560a903abcf6848ee80e  <=  ~I68016caaf170fbe2734c5b6aaf089894 + 1;
                    I63e645f447ddd1fc9409879872479bef  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I62929057b7c214bd38fd532e20ba5623 == I2ccb382adcd7799634c86273c8a39199 ) begin
                    Iee607ab8132caf0f678324d20394f533  <= I169b0fac6d01a713986b636bf8dfc3fb;
                    Ia8298013e67424c2d5fbe03634170080  <=  0;
                end else begin
                    Iee607ab8132caf0f678324d20394f533  <=  ~I169b0fac6d01a713986b636bf8dfc3fb + 1;
                    Ia8298013e67424c2d5fbe03634170080  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I62929057b7c214bd38fd532e20ba5623 == Ie521ecd231d7bfedc8de182c5050f6de ) begin
                    Icc90fd3c992755ac7e4aec1370600e06  <= Iddb14d68b464d04fe9e0b4e62789601a;
                    Ib404a1296714f45ddca6351a918ee875  <=  0;
                end else begin
                    Icc90fd3c992755ac7e4aec1370600e06  <=  ~Iddb14d68b464d04fe9e0b4e62789601a + 1;
                    Ib404a1296714f45ddca6351a918ee875  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I62929057b7c214bd38fd532e20ba5623 == I855892c34f1706745dda4ffc3e5e5a98 ) begin
                    I81e0ea92e07ed7d29b4ab769443b55d3  <= Ie5b71f77beb734a6ab7f7be6c6f9c252;
                    Ic08905e9ffee26c630277db86cd5be95  <=  0;
                end else begin
                    I81e0ea92e07ed7d29b4ab769443b55d3  <=  ~Ie5b71f77beb734a6ab7f7be6c6f9c252 + 1;
                    Ic08905e9ffee26c630277db86cd5be95  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I62929057b7c214bd38fd532e20ba5623 == Ib945fab3df6e5a7494b7fe463384ff4b ) begin
                    Ie7554e9d2bb6287b440973a9effefb50  <= I59f9fa0b81ca88915c338ece1d1e08d5;
                    I674e937c017f29d18946139b00db02d8  <=  0;
                end else begin
                    Ie7554e9d2bb6287b440973a9effefb50  <=  ~I59f9fa0b81ca88915c338ece1d1e08d5 + 1;
                    I674e937c017f29d18946139b00db02d8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I641179f37fef63e7deec603b3291381c == Id4fa22c6f8634ae38892953bd6ab55b5 ) begin
                    I3fd483389e4ddb927e7be7636441f0f1  <= I4f27922ccb21b65dcfe2dc0fcc97cdf3;
                    Ib3f5f61eaba0c2dfdf6c75e46e4233f0  <=  0;
                end else begin
                    I3fd483389e4ddb927e7be7636441f0f1  <=  ~I4f27922ccb21b65dcfe2dc0fcc97cdf3 + 1;
                    Ib3f5f61eaba0c2dfdf6c75e46e4233f0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I641179f37fef63e7deec603b3291381c == I3d8295457058e1d34bb136753b69aaae ) begin
                    I3d7a6bd63d9f66b068c08cf9046474f7  <= Idd7ae55ba748fb36e49684037212936d;
                    Iff1039ba558287ef96daa7dfd15d6294  <=  0;
                end else begin
                    I3d7a6bd63d9f66b068c08cf9046474f7  <=  ~Idd7ae55ba748fb36e49684037212936d + 1;
                    Iff1039ba558287ef96daa7dfd15d6294  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I641179f37fef63e7deec603b3291381c == Ib8df0659486e8ecfb5c52bc2db3a8436 ) begin
                    Ifdb5bd8e8237676fd8d2816bfa53f0c0  <= Ib8da505d1572487e814e7b0682e6dfa9;
                    I017268444024bc19b209dbb4322de15c  <=  0;
                end else begin
                    Ifdb5bd8e8237676fd8d2816bfa53f0c0  <=  ~Ib8da505d1572487e814e7b0682e6dfa9 + 1;
                    I017268444024bc19b209dbb4322de15c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I641179f37fef63e7deec603b3291381c == Ice8927db6ef88a90daf77ea5be2a34bb ) begin
                    If2865b698bf9c511fcf6724856074335  <= Idedb59a6fa2f6ad049f81ac652c645d8;
                    I22e4741c472c64c846742391d81f682c  <=  0;
                end else begin
                    If2865b698bf9c511fcf6724856074335  <=  ~Idedb59a6fa2f6ad049f81ac652c645d8 + 1;
                    I22e4741c472c64c846742391d81f682c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I641179f37fef63e7deec603b3291381c == Ifde5beb333f350ce581a137dae22b99b ) begin
                    I077ad1ef2fe0a7e791fdb45026788641  <= I7d50b49718ab2007accda67ac77a65d0;
                    Ie3c87a536250268b1012b6166173108b  <=  0;
                end else begin
                    I077ad1ef2fe0a7e791fdb45026788641  <=  ~I7d50b49718ab2007accda67ac77a65d0 + 1;
                    Ie3c87a536250268b1012b6166173108b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I641179f37fef63e7deec603b3291381c == I9fe47549e560319ae8decf04a9db5240 ) begin
                    I4c67ed6284da547b599a4602a3cc51dd  <= I27e0600689451a7475a36143f0eb1079;
                    I54204328537dbc383a3a03352e9d6fb6  <=  0;
                end else begin
                    I4c67ed6284da547b599a4602a3cc51dd  <=  ~I27e0600689451a7475a36143f0eb1079 + 1;
                    I54204328537dbc383a3a03352e9d6fb6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 == Idcda31b4dea85b3acd88cad806aef569 ) begin
                    I3d0babc64a3400a1ee57fff14920d1e3  <= Iba6724b61ecb74552b9bb3cab96480c6;
                    Ic5d81213c2d23b0549006ed162d9e6dd  <=  0;
                end else begin
                    I3d0babc64a3400a1ee57fff14920d1e3  <=  ~Iba6724b61ecb74552b9bb3cab96480c6 + 1;
                    Ic5d81213c2d23b0549006ed162d9e6dd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 == I54da9f6048b299dd7e94962912b86407 ) begin
                    Ica1731833fd3d6a881b3a17a5916f7e7  <= I0abb44bd896fbc695e880fee67fb0c42;
                    I0ac628860f9fb9e6daae572ff007f34a  <=  0;
                end else begin
                    Ica1731833fd3d6a881b3a17a5916f7e7  <=  ~I0abb44bd896fbc695e880fee67fb0c42 + 1;
                    I0ac628860f9fb9e6daae572ff007f34a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 == Ib1da5f847077624a37594c2db1b444fc ) begin
                    Id5705e57bc5c050342e82a302b73902e  <= Ifd714548110aa979e735cc6e13d3ef57;
                    I2487101836608b77528a49d037c40fb6  <=  0;
                end else begin
                    Id5705e57bc5c050342e82a302b73902e  <=  ~Ifd714548110aa979e735cc6e13d3ef57 + 1;
                    I2487101836608b77528a49d037c40fb6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 == I80c640a2bc35e9012dfdda839dc5ed1a ) begin
                    I4606e0ec878c615753206459716b5d25  <= Ieeb6c7cdf1379ee3d2933d81bc812dbc;
                    I99d49fb5c921d2d837ac7b02716d9ada  <=  0;
                end else begin
                    I4606e0ec878c615753206459716b5d25  <=  ~Ieeb6c7cdf1379ee3d2933d81bc812dbc + 1;
                    I99d49fb5c921d2d837ac7b02716d9ada  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 == Ic81ffedc7f65fc4d390acd0a30d5e427 ) begin
                    I5ac4f231a175a60f63db8d4d71cfabaf  <= Id682af5250edce8e3811d418ecf2dd10;
                    If4d0af4a78a49e861adbdb1a3f6e7ae9  <=  0;
                end else begin
                    I5ac4f231a175a60f63db8d4d71cfabaf  <=  ~Id682af5250edce8e3811d418ecf2dd10 + 1;
                    If4d0af4a78a49e861adbdb1a3f6e7ae9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iff04b7ec87148f5bd408b4ec4b0590a5 == Ied3448df1f31122d619b1a4cb316f200 ) begin
                    I26a3cd9ec3a564df04ad20559039598f  <= I1d02127e28fb2e9aaf352815627960e7;
                    Iccefd72e7e22a425ced6974251245da8  <=  0;
                end else begin
                    I26a3cd9ec3a564df04ad20559039598f  <=  ~I1d02127e28fb2e9aaf352815627960e7 + 1;
                    Iccefd72e7e22a425ced6974251245da8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa == I017d4243cafbd5d4d615393de3a29aa8 ) begin
                    I26801bb91e66797982b66ce815da85a8  <= Ibee34260749dc92b8523e83cd64d6a40;
                    I3fcc5c32415df9710be01f0f35ac68e5  <=  0;
                end else begin
                    I26801bb91e66797982b66ce815da85a8  <=  ~Ibee34260749dc92b8523e83cd64d6a40 + 1;
                    I3fcc5c32415df9710be01f0f35ac68e5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa == Icb2adb3572c2ac780b4fb413c6ebb375 ) begin
                    I3b617a013c15e8b623ad517e08df3a00  <= Ie9a2a59c7b3571194198dca0c679c5f6;
                    I0bf8339802110abb8bc94e481647f25f  <=  0;
                end else begin
                    I3b617a013c15e8b623ad517e08df3a00  <=  ~Ie9a2a59c7b3571194198dca0c679c5f6 + 1;
                    I0bf8339802110abb8bc94e481647f25f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa == I711042dda213300a90c51b09057b64b4 ) begin
                    I65f5f9a3f7f68f4b2fd7695ce6bf4629  <= Ie4b5a941feb385e88498a98e5f8ddc01;
                    I6ae57b8d68417d1ea8ef70d43a943e0b  <=  0;
                end else begin
                    I65f5f9a3f7f68f4b2fd7695ce6bf4629  <=  ~Ie4b5a941feb385e88498a98e5f8ddc01 + 1;
                    I6ae57b8d68417d1ea8ef70d43a943e0b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa == I59b7772e832e814877d4f9e7726f5143 ) begin
                    I7d405b59e360b17d7f2eb1805b796fa9  <= I30b2b34a0cecfdbdeecba5f286befccd;
                    I07dd0ed55fbdeaace398ab7644a5189f  <=  0;
                end else begin
                    I7d405b59e360b17d7f2eb1805b796fa9  <=  ~I30b2b34a0cecfdbdeecba5f286befccd + 1;
                    I07dd0ed55fbdeaace398ab7644a5189f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa == Ida6ee8eeec2fa7a6bc1eeb8b5c3fbffd ) begin
                    I033ad5c570f42830b265d7bf6a102757  <= I8ce739ddc344cacb2de7f2c88a882170;
                    I69cfa3967387c5e8e48994b6466673a0  <=  0;
                end else begin
                    I033ad5c570f42830b265d7bf6a102757  <=  ~I8ce739ddc344cacb2de7f2c88a882170 + 1;
                    I69cfa3967387c5e8e48994b6466673a0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I198bfb18d6f91c8f62777e6f592a88fa == Ic7fb6a8351310bd93953232556a692ab ) begin
                    Ia00376ef5aca6a428280f2dbf25ab1cb  <= I8b00260bb93e928e66e9d4aaeb0d9b55;
                    I2ce599e7a40a71d9fe09f80269accc31  <=  0;
                end else begin
                    Ia00376ef5aca6a428280f2dbf25ab1cb  <=  ~I8b00260bb93e928e66e9d4aaeb0d9b55 + 1;
                    I2ce599e7a40a71d9fe09f80269accc31  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 == Ib2ff62fd117b50bc0c190b8111b85f4b ) begin
                    I252b17144e39018fda208bd18b555c09  <= I9c1ca916654bad308af37d040b486cf8;
                    Id424746e76cc70f9292ed41659973621  <=  0;
                end else begin
                    I252b17144e39018fda208bd18b555c09  <=  ~I9c1ca916654bad308af37d040b486cf8 + 1;
                    Id424746e76cc70f9292ed41659973621  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 == I4d46847f77bb17019eaba7ead1549a87 ) begin
                    Idb756c313694457c14b02431f3f076c7  <= I05749703a8a131453c563ed2264680a7;
                    I45528f9be6a8f9a0f646d83223307e79  <=  0;
                end else begin
                    Idb756c313694457c14b02431f3f076c7  <=  ~I05749703a8a131453c563ed2264680a7 + 1;
                    I45528f9be6a8f9a0f646d83223307e79  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 == I1d6145f5c5d5049a1ba3f3ef8a09924e ) begin
                    I0c1545b312d755b14ee27b399a1d3079  <= I4b76fe5f9863a41733b76decf9867d16;
                    Iabcd2910bddf2e544c707c553b2ef370  <=  0;
                end else begin
                    I0c1545b312d755b14ee27b399a1d3079  <=  ~I4b76fe5f9863a41733b76decf9867d16 + 1;
                    Iabcd2910bddf2e544c707c553b2ef370  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 == Ie5e08b5111cd2baacecc68000f84a9ef ) begin
                    I903842d13327b74a952be0aa6c7ab0e8  <= I2805bb16fd574a64de548b39a532cd8a;
                    If01521dbf7dd9aa5196a9130ba47b149  <=  0;
                end else begin
                    I903842d13327b74a952be0aa6c7ab0e8  <=  ~I2805bb16fd574a64de548b39a532cd8a + 1;
                    If01521dbf7dd9aa5196a9130ba47b149  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 == I3d61c9137cc0cdc892bc50c659fa8c47 ) begin
                    Ic461c1b7bd09b59297193d388c525ece  <= Ide6a696c06f17f455d56bb28cad98bd0;
                    I9284cc53534eaf3d6e5b4e9d9d93bea5  <=  0;
                end else begin
                    Ic461c1b7bd09b59297193d388c525ece  <=  ~Ide6a696c06f17f455d56bb28cad98bd0 + 1;
                    I9284cc53534eaf3d6e5b4e9d9d93bea5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia1562c88b4f56d8935c3a5d6ead0f816 == I15411a1495f104308964c62a1ac7fe6a ) begin
                    Ia14490057ef27f5df5f1b23ca6440a65  <= I39bce1f71ede4663c187ddfd6501eda1;
                    Id5fdf11f0bf10ec37b11ced0a3268ad7  <=  0;
                end else begin
                    Ia14490057ef27f5df5f1b23ca6440a65  <=  ~I39bce1f71ede4663c187ddfd6501eda1 + 1;
                    Id5fdf11f0bf10ec37b11ced0a3268ad7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 == I99f350aa0b468f89e8ac4b3da627a81a ) begin
                    I2d3c1e36bd952fdbe4fac5f3af07e666  <= Id0e769bee61ae0a90c167fab061f5965;
                    I36cc6827c8e4c7831078c8f9972ee78a  <=  0;
                end else begin
                    I2d3c1e36bd952fdbe4fac5f3af07e666  <=  ~Id0e769bee61ae0a90c167fab061f5965 + 1;
                    I36cc6827c8e4c7831078c8f9972ee78a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 == Ie23efd54df7880569e2d45a8572c02ba ) begin
                    I7fcea0a5f9987b2414ab443bd07c05ad  <= I83e03af8657a4a237641a9da7922e502;
                    Ied6cdc5d7aa6335b2c32d8ab6ee6d889  <=  0;
                end else begin
                    I7fcea0a5f9987b2414ab443bd07c05ad  <=  ~I83e03af8657a4a237641a9da7922e502 + 1;
                    Ied6cdc5d7aa6335b2c32d8ab6ee6d889  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 == I29de3d73d38639aacb693c8080f4a168 ) begin
                    If0f5bf08d96033f6281121230c1e47c9  <= I7565e071282ca6e77bb469afc522f1a2;
                    I70709dd8c55168e62143f56d0bda1239  <=  0;
                end else begin
                    If0f5bf08d96033f6281121230c1e47c9  <=  ~I7565e071282ca6e77bb469afc522f1a2 + 1;
                    I70709dd8c55168e62143f56d0bda1239  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 == I09fe5010524903c8b34892f6c308d670 ) begin
                    I19412627d5c573ceaa981cd7f1027e83  <= I5d0dc5d40385ab67bc7f540f212b6a97;
                    I73ce9bd4312ce9a6cdc0c6b6aec72a55  <=  0;
                end else begin
                    I19412627d5c573ceaa981cd7f1027e83  <=  ~I5d0dc5d40385ab67bc7f540f212b6a97 + 1;
                    I73ce9bd4312ce9a6cdc0c6b6aec72a55  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 == Id1af840781c6093921ea2feef85b6bb7 ) begin
                    I7c72a1709b233f745fb0323d04bfeb1a  <= I548cac395730b8386670cc4c7a64319a;
                    I9d0fc48c488109406aa9cfef80ac3b48  <=  0;
                end else begin
                    I7c72a1709b233f745fb0323d04bfeb1a  <=  ~I548cac395730b8386670cc4c7a64319a + 1;
                    I9d0fc48c488109406aa9cfef80ac3b48  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iaccba3030d9d9f8a56f86d6e34ed6325 == Iab8c6e113a90faf59bb550681b0dc7f7 ) begin
                    I2639cefc25ac6f4982e4eeccf8fa810e  <= Ic6d9bbbfb7890540edd10aa5758b0c4b;
                    Ie09336ee55ee45ac0297849f7b814f4d  <=  0;
                end else begin
                    I2639cefc25ac6f4982e4eeccf8fa810e  <=  ~Ic6d9bbbfb7890540edd10aa5758b0c4b + 1;
                    Ie09336ee55ee45ac0297849f7b814f4d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 == I2110f3928229bc70d8ec9ec7f1c92520 ) begin
                    I76340f05f74b295583bd9353884979be  <= I7beb1f915a881a302f93c869d81417d1;
                    If919b9778437e1c4366017968d1ea582  <=  0;
                end else begin
                    I76340f05f74b295583bd9353884979be  <=  ~I7beb1f915a881a302f93c869d81417d1 + 1;
                    If919b9778437e1c4366017968d1ea582  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 == I0befd079483b2da8d410fa137f71d801 ) begin
                    I00974459262f29ec2b5472472e49faf6  <= I5fc389bbc1ce31f7b326da719dc576d4;
                    I71cdff133cb7a645e623c4bf06588fc3  <=  0;
                end else begin
                    I00974459262f29ec2b5472472e49faf6  <=  ~I5fc389bbc1ce31f7b326da719dc576d4 + 1;
                    I71cdff133cb7a645e623c4bf06588fc3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 == Icd1a2b8c1a50f9a1bab48ebfbb87ca73 ) begin
                    I075efbd3c4d87df8d733f0b3db008b1f  <= I922e6f05f7c6e0f6f0b1a5c9548df238;
                    Ie7fd0410103d16e27611f9ac30c657da  <=  0;
                end else begin
                    I075efbd3c4d87df8d733f0b3db008b1f  <=  ~I922e6f05f7c6e0f6f0b1a5c9548df238 + 1;
                    Ie7fd0410103d16e27611f9ac30c657da  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 == I4422278d28ff2a983cc3a4ad8f2d655f ) begin
                    If8bd6a5d380075f1ee7f7a4542531dbe  <= I8c6bb234a1ca3deba637adf746672194;
                    Iab93975104312336985d4736015098b4  <=  0;
                end else begin
                    If8bd6a5d380075f1ee7f7a4542531dbe  <=  ~I8c6bb234a1ca3deba637adf746672194 + 1;
                    Iab93975104312336985d4736015098b4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 == I3fc4400a93546df2e2aad374a4d8c7e4 ) begin
                    Ib81b730d107434503c988ab9f00e1605  <= Ide24ebd7423d4c4f43577b019f2e30e4;
                    I564a4d4a94f9951d85287b2ac35479fe  <=  0;
                end else begin
                    Ib81b730d107434503c988ab9f00e1605  <=  ~Ide24ebd7423d4c4f43577b019f2e30e4 + 1;
                    I564a4d4a94f9951d85287b2ac35479fe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I953dfeeacee8c44c08d0a425fa549e49 == I6c6a02b572e98d30ea5a0406be5cfd11 ) begin
                    Ib05cffa1bb31054450391bf9e17f8ef9  <= Ifc412122eab7560c9021a17d7f8700c4;
                    I09c5b4146a3c48ae706d3041ddfe074d  <=  0;
                end else begin
                    Ib05cffa1bb31054450391bf9e17f8ef9  <=  ~Ifc412122eab7560c9021a17d7f8700c4 + 1;
                    I09c5b4146a3c48ae706d3041ddfe074d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 == I91c29953d4b53657da39b53d8c909fd8 ) begin
                    I627097c06e3be5a4385171f3ec7ae5c9  <= Ia5a56ed2c6b98e72002c6c5f946e7264;
                    If205c7d745e5372ea61afa389f1af2c2  <=  0;
                end else begin
                    I627097c06e3be5a4385171f3ec7ae5c9  <=  ~Ia5a56ed2c6b98e72002c6c5f946e7264 + 1;
                    If205c7d745e5372ea61afa389f1af2c2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 == I10441dc2915fcece28b38aa6b4156f5c ) begin
                    I76e2c6001e1ae97670539bd471fc74e8  <= Ia888ed8885f66084b777f66e25cef1e7;
                    Ief37a022c34d4e670413f5b7db306876  <=  0;
                end else begin
                    I76e2c6001e1ae97670539bd471fc74e8  <=  ~Ia888ed8885f66084b777f66e25cef1e7 + 1;
                    Ief37a022c34d4e670413f5b7db306876  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 == Id26aa7283f70b13f1eb0b97ab1222da7 ) begin
                    I8b4433056d26f4aa60f18418b0114930  <= I248229aecef00b87a70ce88920e407f5;
                    I5ac36d471eec2b3ac068a2d20283f674  <=  0;
                end else begin
                    I8b4433056d26f4aa60f18418b0114930  <=  ~I248229aecef00b87a70ce88920e407f5 + 1;
                    I5ac36d471eec2b3ac068a2d20283f674  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 == I98b4bf6c27d9420941d252a98806344c ) begin
                    I99601176686afd8fb85a85ec43849e6f  <= I3d162a0ec918f220a7d5f4efdf89cb58;
                    I68acc6967dd156d6373abd6cc620f247  <=  0;
                end else begin
                    I99601176686afd8fb85a85ec43849e6f  <=  ~I3d162a0ec918f220a7d5f4efdf89cb58 + 1;
                    I68acc6967dd156d6373abd6cc620f247  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 == I7814b43f7573d005d6b9350b311f93df ) begin
                    Iad8276d5be3d9c6fc085465f05ac2aed  <= I1ca0372f60e48f2f803778c9017023c0;
                    Ic830033c7861645951982dc630e3385b  <=  0;
                end else begin
                    Iad8276d5be3d9c6fc085465f05ac2aed  <=  ~I1ca0372f60e48f2f803778c9017023c0 + 1;
                    Ic830033c7861645951982dc630e3385b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I214a50bf9f879fe747904f4679fdd1f6 == Ia378bb83b0f76d4bf7de347a8bfd20cb ) begin
                    I5e5dfce3ceb4fbbfce344bd471901736  <= Ieb9693d54f0808b0ba463fd3c316a80e;
                    I7f9305c8bfe731300ad0a9d1ece97db4  <=  0;
                end else begin
                    I5e5dfce3ceb4fbbfce344bd471901736  <=  ~Ieb9693d54f0808b0ba463fd3c316a80e + 1;
                    I7f9305c8bfe731300ad0a9d1ece97db4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d == Ie814322ac906e4bc9baa42fef66e9b8e ) begin
                    I22ace766690e445ff36176eac2473368  <= I63da03315d7e51fcacb0bc0298e506ed;
                    I0bb61f163279dc993a94e647611f6e06  <=  0;
                end else begin
                    I22ace766690e445ff36176eac2473368  <=  ~I63da03315d7e51fcacb0bc0298e506ed + 1;
                    I0bb61f163279dc993a94e647611f6e06  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d == Ic3f5c7e9a546509687973efde6a8a8f7 ) begin
                    I896c57162e4384f021d822789b4c01a3  <= I918f5a12e96bb96941f019940f27a5be;
                    Ib5effb1b2c147179bc8c8febce7657c7  <=  0;
                end else begin
                    I896c57162e4384f021d822789b4c01a3  <=  ~I918f5a12e96bb96941f019940f27a5be + 1;
                    Ib5effb1b2c147179bc8c8febce7657c7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d == I5a7668981b781cea8cd3de0aa6687bc1 ) begin
                    I3d0367a799090b3c9048235436a39063  <= Ib4fb115f442ff544fa3d21b4e9d3f075;
                    I81dd944eccdd3dd6fd84727d21efd0ac  <=  0;
                end else begin
                    I3d0367a799090b3c9048235436a39063  <=  ~Ib4fb115f442ff544fa3d21b4e9d3f075 + 1;
                    I81dd944eccdd3dd6fd84727d21efd0ac  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d == I4951067363d095f73676e08c2be255fa ) begin
                    Ic0f25799f0dc7cc33de95e47ebcc083a  <= I387403482432a3196109484d1120d584;
                    I986e7c899df08e35fa2347e282e8c90e  <=  0;
                end else begin
                    Ic0f25799f0dc7cc33de95e47ebcc083a  <=  ~I387403482432a3196109484d1120d584 + 1;
                    I986e7c899df08e35fa2347e282e8c90e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d == Ia02db0467aa519e8920344525ed30dfb ) begin
                    I7186b368e297d0db1f746c6241eae65d  <= I619af17eaa4a56726d6ab322a74dd0a4;
                    Idb764022b3ae49281c7b82f6e309cca9  <=  0;
                end else begin
                    I7186b368e297d0db1f746c6241eae65d  <=  ~I619af17eaa4a56726d6ab322a74dd0a4 + 1;
                    Idb764022b3ae49281c7b82f6e309cca9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic88f2c344a8ad254fc7d7034cb594f6d == I303114e80311c7f6552446bbcb0fe6a9 ) begin
                    I21d63f6fe5c72798aa4636527c02613d  <= I7a67ed3bb370520d0d25ce407ab8cd8b;
                    I311eb64d22cff4b1424f3ccdd33dec45  <=  0;
                end else begin
                    I21d63f6fe5c72798aa4636527c02613d  <=  ~I7a67ed3bb370520d0d25ce407ab8cd8b + 1;
                    I311eb64d22cff4b1424f3ccdd33dec45  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If299d1a4e044acbc70bc3b7bce9f86e9 == I7a5c09537045dcd633095a86a6c530ed ) begin
                    I15e0219f2da6f52177e76580198d0e6c  <= I7629b35ca548190a81021a2c13d8919b;
                    I128183dffb32a1461db0c2b851559f68  <=  0;
                end else begin
                    I15e0219f2da6f52177e76580198d0e6c  <=  ~I7629b35ca548190a81021a2c13d8919b + 1;
                    I128183dffb32a1461db0c2b851559f68  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If299d1a4e044acbc70bc3b7bce9f86e9 == I6aac30f1ecc270161a81bccffab85efa ) begin
                    I4cac308bee8801c4f9716673e39da4ab  <= I004851d3828f135ebe4d2e6ab83936bf;
                    I817fbe1f44196264e2531197ca8da9ea  <=  0;
                end else begin
                    I4cac308bee8801c4f9716673e39da4ab  <=  ~I004851d3828f135ebe4d2e6ab83936bf + 1;
                    I817fbe1f44196264e2531197ca8da9ea  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If299d1a4e044acbc70bc3b7bce9f86e9 == I79b86b24bfa472a80487e7ea64f9dd82 ) begin
                    I6f4f7b4e45a495fe139955e0605ff208  <= I0e2c382b2e62ed43b76697230e34b719;
                    I3e74c445193a1c9ec9dcb31f4aef2117  <=  0;
                end else begin
                    I6f4f7b4e45a495fe139955e0605ff208  <=  ~I0e2c382b2e62ed43b76697230e34b719 + 1;
                    I3e74c445193a1c9ec9dcb31f4aef2117  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If299d1a4e044acbc70bc3b7bce9f86e9 == I208d1c07cebe2f45b25b562dd9109f7e ) begin
                    I79ae5f2981b7dd91141b0a22f012f4b1  <= I36dac27d10701db70fb2b5996a3f038f;
                    I70f3cac8f36ef943672bbe7a9d6be5ed  <=  0;
                end else begin
                    I79ae5f2981b7dd91141b0a22f012f4b1  <=  ~I36dac27d10701db70fb2b5996a3f038f + 1;
                    I70f3cac8f36ef943672bbe7a9d6be5ed  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idb373d2cf788f6a93a0e5df7f9179292 == I86a3b6dc06c6c99cb1fa88023d920423 ) begin
                    Id4b4d757e50bc2721e8725ae10d88c9e  <= I51d62ebd160eb0d073a7efb64d20079a;
                    I26b4d738c45246201073f4b4a786078a  <=  0;
                end else begin
                    Id4b4d757e50bc2721e8725ae10d88c9e  <=  ~I51d62ebd160eb0d073a7efb64d20079a + 1;
                    I26b4d738c45246201073f4b4a786078a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idb373d2cf788f6a93a0e5df7f9179292 == I9c0e0297c0e5042f1ed791d9d97a6f37 ) begin
                    I4513152c34d5d00ddcc4f099481f659d  <= Ib3545a88d68631af1c94ca2cb1f379af;
                    I6c4f341b9eeda21a97806084196421d3  <=  0;
                end else begin
                    I4513152c34d5d00ddcc4f099481f659d  <=  ~Ib3545a88d68631af1c94ca2cb1f379af + 1;
                    I6c4f341b9eeda21a97806084196421d3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idb373d2cf788f6a93a0e5df7f9179292 == I3af891fd5da91085a79886d82e6bdf48 ) begin
                    I7bd4e77993fdd5a0833f1cdc7a382b56  <= I81ad7b044118734f4dc32a1a4e8eba31;
                    Ibdf325321ebd9a7baa25435537c159bb  <=  0;
                end else begin
                    I7bd4e77993fdd5a0833f1cdc7a382b56  <=  ~I81ad7b044118734f4dc32a1a4e8eba31 + 1;
                    Ibdf325321ebd9a7baa25435537c159bb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idb373d2cf788f6a93a0e5df7f9179292 == Ia1c63f27861c8e594f01ffb31a29ba0a ) begin
                    I13b0d404e7a96cd53147b574b242ef41  <= I5ad8c235d46349b6d310d0f175f84288;
                    I626a4c66bf0cca36dfa2bcd8c24bff35  <=  0;
                end else begin
                    I13b0d404e7a96cd53147b574b242ef41  <=  ~I5ad8c235d46349b6d310d0f175f84288 + 1;
                    I626a4c66bf0cca36dfa2bcd8c24bff35  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic73b8c8f76a985330d4ac1fa0cc28e7f == I62b87c6aa6ba054ab5e80842ea738020 ) begin
                    I4acc3bfa99b152c6ef6d11608f639b70  <= Ibc00920378e2427df2a63a47dc3eaded;
                    Icd6ab7be501038196ab2674cdf764453  <=  0;
                end else begin
                    I4acc3bfa99b152c6ef6d11608f639b70  <=  ~Ibc00920378e2427df2a63a47dc3eaded + 1;
                    Icd6ab7be501038196ab2674cdf764453  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic73b8c8f76a985330d4ac1fa0cc28e7f == I429241122829d9e51a3db90b33a44ac3 ) begin
                    Ia1ec7ba972ec6f0049c4cf00b9d42125  <= Ic5195bbaa69d95059cca6e152dc9f705;
                    I31c6d68ecdb4d0a6790a12343f59731b  <=  0;
                end else begin
                    Ia1ec7ba972ec6f0049c4cf00b9d42125  <=  ~Ic5195bbaa69d95059cca6e152dc9f705 + 1;
                    I31c6d68ecdb4d0a6790a12343f59731b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic73b8c8f76a985330d4ac1fa0cc28e7f == I162416616ce392c679d22b115c192356 ) begin
                    I4fb5494e6f04e29d76bb8d3bc8bf6cd9  <= Ia01f20e0bcf35c2ee4963e9c392c1004;
                    I8eb06ffb6aca72c66cea97d9caa26f1c  <=  0;
                end else begin
                    I4fb5494e6f04e29d76bb8d3bc8bf6cd9  <=  ~Ia01f20e0bcf35c2ee4963e9c392c1004 + 1;
                    I8eb06ffb6aca72c66cea97d9caa26f1c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic73b8c8f76a985330d4ac1fa0cc28e7f == I62edec03adbb7bbda313abc2220a6a5f ) begin
                    Iaffb0ef4e18bb7b582275b43684fcf3d  <= I9f6f48fea88d1cd73ef2b24c7e819964;
                    I35ecf6ebd98d91d12361beef01dadfbe  <=  0;
                end else begin
                    Iaffb0ef4e18bb7b582275b43684fcf3d  <=  ~I9f6f48fea88d1cd73ef2b24c7e819964 + 1;
                    I35ecf6ebd98d91d12361beef01dadfbe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I134dfb2c57d8cdffd2789e2f442c3247 == Ic3e192f5abb5526a54ea249e736702b7 ) begin
                    Ia5e3649f8e32a81606ee34353c54350a  <= I847feea780cc8a06caea2d2ea79ad281;
                    If73961b42bf31d49c78c3fbe86f8d2cb  <=  0;
                end else begin
                    Ia5e3649f8e32a81606ee34353c54350a  <=  ~I847feea780cc8a06caea2d2ea79ad281 + 1;
                    If73961b42bf31d49c78c3fbe86f8d2cb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I134dfb2c57d8cdffd2789e2f442c3247 == I1ae99cfc5ded208c2dbadbabf36fd629 ) begin
                    Ic675cf7eac5ece436feb5a8acd642f6b  <= I7ef6f4aeda7fd6775839c068c681f9bc;
                    I560157aede2c2c3b6dce019e2fb4314c  <=  0;
                end else begin
                    Ic675cf7eac5ece436feb5a8acd642f6b  <=  ~I7ef6f4aeda7fd6775839c068c681f9bc + 1;
                    I560157aede2c2c3b6dce019e2fb4314c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I134dfb2c57d8cdffd2789e2f442c3247 == I1ef8bfbeda31b3dbbff053cd36de4859 ) begin
                    I71357943bbe307c9ae9099d4bcbff882  <= I0645e741da20a4957747188273a655b1;
                    I075a8e7435a4fbe97304b4d379bcfee4  <=  0;
                end else begin
                    I71357943bbe307c9ae9099d4bcbff882  <=  ~I0645e741da20a4957747188273a655b1 + 1;
                    I075a8e7435a4fbe97304b4d379bcfee4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I134dfb2c57d8cdffd2789e2f442c3247 == I6d76fd8af44893ab0f82a282aca12377 ) begin
                    Ib2684f54caebb1a1c079a2a4f2cf0dab  <= I71125dffdd2d37e44dbb46143c1e8d9a;
                    I09a1ad6a0fba78d4984fee238fd95bd7  <=  0;
                end else begin
                    Ib2684f54caebb1a1c079a2a4f2cf0dab  <=  ~I71125dffdd2d37e44dbb46143c1e8d9a + 1;
                    I09a1ad6a0fba78d4984fee238fd95bd7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c735e43be8030078ec10bdb6882e79c == I86247340bd399afebac1ffe403a3331e ) begin
                    If19836577f9a254b365f0dcfe0ae55ce  <= I50c166f958b22ce866cd40334918274c;
                    I5c03de756d46517f2158e4ffb019edd3  <=  0;
                end else begin
                    If19836577f9a254b365f0dcfe0ae55ce  <=  ~I50c166f958b22ce866cd40334918274c + 1;
                    I5c03de756d46517f2158e4ffb019edd3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c735e43be8030078ec10bdb6882e79c == Id932053ac235b3035e2f3d5986b7d398 ) begin
                    I2f47a00b58779b836c08b472d305b031  <= Icd225144fd331b870847044b4d02bed0;
                    Ia897f60b5c256180be523c5ff8ba6b77  <=  0;
                end else begin
                    I2f47a00b58779b836c08b472d305b031  <=  ~Icd225144fd331b870847044b4d02bed0 + 1;
                    Ia897f60b5c256180be523c5ff8ba6b77  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c735e43be8030078ec10bdb6882e79c == I4b43b5eb71dffb4bcb9ee541a537b427 ) begin
                    I8b2593fd0e35c37f68097187a41596e2  <= I5e876482090ce6007c2a2f2101c24654;
                    I81a7d30b51b1d7f9d9bc9a97d2f3caac  <=  0;
                end else begin
                    I8b2593fd0e35c37f68097187a41596e2  <=  ~I5e876482090ce6007c2a2f2101c24654 + 1;
                    I81a7d30b51b1d7f9d9bc9a97d2f3caac  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c735e43be8030078ec10bdb6882e79c == Ib481c772e0ef5d172f6b079dc8df1ae1 ) begin
                    Ibbcdc1c30d3333cbec65d264890cf3e5  <= I026ded06f56d9ca93f47fd85aec4f7ad;
                    If46a830ca08eeb2b8b3d8b2f996491e8  <=  0;
                end else begin
                    Ibbcdc1c30d3333cbec65d264890cf3e5  <=  ~I026ded06f56d9ca93f47fd85aec4f7ad + 1;
                    If46a830ca08eeb2b8b3d8b2f996491e8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0c735e43be8030078ec10bdb6882e79c == I2e046a6e848cf2da29e103872a10c26d ) begin
                    Iec6e9640b0494777c013c97613855ce7  <= Iec596e94ec168a564bccbbaa7df833c9;
                    I13e6271176ef80d03f8878441893c467  <=  0;
                end else begin
                    Iec6e9640b0494777c013c97613855ce7  <=  ~Iec596e94ec168a564bccbbaa7df833c9 + 1;
                    I13e6271176ef80d03f8878441893c467  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9951415c1d599570af1787767caa2dc == I2a64ca51e05db642281525ccc7cf9a06 ) begin
                    Ic10f396b52dda0dcfbf2a847cfed617c  <= Ib514e01c261e43a725582a10596eed32;
                    Idb5b4ae9bb42a053d9db8b8c71a0b9cc  <=  0;
                end else begin
                    Ic10f396b52dda0dcfbf2a847cfed617c  <=  ~Ib514e01c261e43a725582a10596eed32 + 1;
                    Idb5b4ae9bb42a053d9db8b8c71a0b9cc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9951415c1d599570af1787767caa2dc == I4275f1683058cfab72e02f2631d2ee96 ) begin
                    I94ebfb633f3272b8f40303ce768f0ade  <= Ic19a62cdecb2329370f7e11c48d3738d;
                    I96c6deed53888cfe0b1fcbe6832a1d61  <=  0;
                end else begin
                    I94ebfb633f3272b8f40303ce768f0ade  <=  ~Ic19a62cdecb2329370f7e11c48d3738d + 1;
                    I96c6deed53888cfe0b1fcbe6832a1d61  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9951415c1d599570af1787767caa2dc == I592fab4d3d2c1bb3956b89eabc06dc56 ) begin
                    Ie975a6fd78adbad8b8a56bd6a3802e4f  <= Ib2f5691baa59adfbaad62f6ffc71fb05;
                    Ibb40e3b624d2f19eeccfe071e540021a  <=  0;
                end else begin
                    Ie975a6fd78adbad8b8a56bd6a3802e4f  <=  ~Ib2f5691baa59adfbaad62f6ffc71fb05 + 1;
                    Ibb40e3b624d2f19eeccfe071e540021a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9951415c1d599570af1787767caa2dc == I6520a98d1357fc57d687f9ea9a60508b ) begin
                    Ib852991e38422ba6de5e18a879ddc3f9  <= I9bdfaca6112385deb86e24ad7e45bbaa;
                    I93bd27a068e6fd416060bd5d919b3451  <=  0;
                end else begin
                    Ib852991e38422ba6de5e18a879ddc3f9  <=  ~I9bdfaca6112385deb86e24ad7e45bbaa + 1;
                    I93bd27a068e6fd416060bd5d919b3451  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9951415c1d599570af1787767caa2dc == I8a022ff37fcd6f34531af4dc7f31a223 ) begin
                    Ife665c9aa6794cccffd04923f4359047  <= I0e647bb8351cfe7828423e7099525585;
                    Iaf516c91fe1544bd0a6f671635eda05d  <=  0;
                end else begin
                    Ife665c9aa6794cccffd04923f4359047  <=  ~I0e647bb8351cfe7828423e7099525585 + 1;
                    Iaf516c91fe1544bd0a6f671635eda05d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2630f187d63ba9b0af52c77093e6b760 == Ia95cd411b17d1c5aaf9e5b583e9398a6 ) begin
                    I076cbc669ff4fb135ffc85910c888241  <= I185b758fb3e50bcfb1464fe2ab593cfe;
                    I6029a024d76e9357223c6fea077501c3  <=  0;
                end else begin
                    I076cbc669ff4fb135ffc85910c888241  <=  ~I185b758fb3e50bcfb1464fe2ab593cfe + 1;
                    I6029a024d76e9357223c6fea077501c3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2630f187d63ba9b0af52c77093e6b760 == I526597e8561c75326b96e85743420a1e ) begin
                    I50245c953aab8c513b17b894afb36a6c  <= Ie25e944f9e3100c39b69bb38dffca177;
                    I8dd3c6c27d8fea2b67906c78715c5854  <=  0;
                end else begin
                    I50245c953aab8c513b17b894afb36a6c  <=  ~Ie25e944f9e3100c39b69bb38dffca177 + 1;
                    I8dd3c6c27d8fea2b67906c78715c5854  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2630f187d63ba9b0af52c77093e6b760 == If2c489abf57879ea491d9a95ce7e1cc1 ) begin
                    I33ac557ef59d79e8b1b359e499a00119  <= I8e77032a54376578b3d16799e30c97f7;
                    I244ab0a87c282939527938b5d43c90e8  <=  0;
                end else begin
                    I33ac557ef59d79e8b1b359e499a00119  <=  ~I8e77032a54376578b3d16799e30c97f7 + 1;
                    I244ab0a87c282939527938b5d43c90e8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2630f187d63ba9b0af52c77093e6b760 == I1dfa9cd65fb0f7c62439bc0d9539e45d ) begin
                    I173fd30c1a5367b61e3fda352365f557  <= I4cd2a7f8f8ec378200b00d03e447ac92;
                    I8b9861dd9f6dbeaedffc07a3e088cf49  <=  0;
                end else begin
                    I173fd30c1a5367b61e3fda352365f557  <=  ~I4cd2a7f8f8ec378200b00d03e447ac92 + 1;
                    I8b9861dd9f6dbeaedffc07a3e088cf49  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2630f187d63ba9b0af52c77093e6b760 == I5799e21b9e2fdc554f8ec65b98120544 ) begin
                    Id6f5041043fa4fd352e74016c4e7de48  <= I1b3c55aca0da232cf3f81d6d0914729f;
                    I71c3dc98a45a807f146ec052c8a9fb82  <=  0;
                end else begin
                    Id6f5041043fa4fd352e74016c4e7de48  <=  ~I1b3c55aca0da232cf3f81d6d0914729f + 1;
                    I71c3dc98a45a807f146ec052c8a9fb82  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 == Id109dde61c0ee952c9053905ee54ccd8 ) begin
                    I6d863254c7f0b52f803b2af4b184f99d  <= I34c76f1a126120c4474e750e9b51e034;
                    Iaa6c753b09c2244d22a8680d73670deb  <=  0;
                end else begin
                    I6d863254c7f0b52f803b2af4b184f99d  <=  ~I34c76f1a126120c4474e750e9b51e034 + 1;
                    Iaa6c753b09c2244d22a8680d73670deb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 == Iafef3ac31f22ba4f5ef06b13165e97eb ) begin
                    I1eeb9c94908cc9ddeb8e3904a145ec6e  <= I0edb624c344787066a2267757052196b;
                    Id8e40a0bd35259f34ffc971eaa7f2fc5  <=  0;
                end else begin
                    I1eeb9c94908cc9ddeb8e3904a145ec6e  <=  ~I0edb624c344787066a2267757052196b + 1;
                    Id8e40a0bd35259f34ffc971eaa7f2fc5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 == Ifc59d693d6dc2fa6848f37a134fbb316 ) begin
                    I6211e241282624fc50fb4ca1842ff9db  <= Ia8443f199838742595ac114f35c00143;
                    I59df806ee758f4db794635ec24232ae9  <=  0;
                end else begin
                    I6211e241282624fc50fb4ca1842ff9db  <=  ~Ia8443f199838742595ac114f35c00143 + 1;
                    I59df806ee758f4db794635ec24232ae9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 == Ie83012a17bd2730837939cf0454395c3 ) begin
                    Iba09e22ece1eb1639d2bb940d3273fe0  <= Ib25b8a538c9d64880e114bf4a80ca42e;
                    I7bd8b1c89a39e4dccbde5c5e040c162f  <=  0;
                end else begin
                    Iba09e22ece1eb1639d2bb940d3273fe0  <=  ~Ib25b8a538c9d64880e114bf4a80ca42e + 1;
                    I7bd8b1c89a39e4dccbde5c5e040c162f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I83db667ace2f04ef4950e2c186e0e6a4 == I1f37257664651a57575f7ae53ab4e180 ) begin
                    I2fe99e4fb8c660d83508bff50ab4929b  <= I25f6a3d7bb869082e4dbbd0ee8574c95;
                    Id3d37273d55ba1de64f97f6d11e704d7  <=  0;
                end else begin
                    I2fe99e4fb8c660d83508bff50ab4929b  <=  ~I25f6a3d7bb869082e4dbbd0ee8574c95 + 1;
                    Id3d37273d55ba1de64f97f6d11e704d7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 == Ibdf8f7dadf142fe8a166328bb5461308 ) begin
                    Ia73db0428763da3c0feffc94a8a8f4f1  <= If96057023747a1538d9f06966af48bc2;
                    I4ff07696ccaf99e49d575694d3a2670e  <=  0;
                end else begin
                    Ia73db0428763da3c0feffc94a8a8f4f1  <=  ~If96057023747a1538d9f06966af48bc2 + 1;
                    I4ff07696ccaf99e49d575694d3a2670e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 == I0ce12cc00bd66d743ab82e89887190dc ) begin
                    I6542fbca90e189048b15deaa3af5d836  <= I199e995390462e06853b1f5cdbd46e0a;
                    Ib89e0144bfc6be3be9a06a08e4f297ca  <=  0;
                end else begin
                    I6542fbca90e189048b15deaa3af5d836  <=  ~I199e995390462e06853b1f5cdbd46e0a + 1;
                    Ib89e0144bfc6be3be9a06a08e4f297ca  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 == I70145dd478e7f0c74c0299cdc0ab8ad5 ) begin
                    Ieacf022fc976bf397946d6481468d6a4  <= Iec6325d585ddd0a9f86bb5cd0229960d;
                    Ife372091864d6ae9b770b69db66ff3ca  <=  0;
                end else begin
                    Ieacf022fc976bf397946d6481468d6a4  <=  ~Iec6325d585ddd0a9f86bb5cd0229960d + 1;
                    Ife372091864d6ae9b770b69db66ff3ca  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 == I03d54826d217e4209d0e0f82beda4100 ) begin
                    I1cef7e6e0555e076b68bbc57de8f289f  <= I4be1ccfec148a522fbf5b8375245cbb3;
                    Ie81b8b84cc2795e2e92168bfa496ece4  <=  0;
                end else begin
                    I1cef7e6e0555e076b68bbc57de8f289f  <=  ~I4be1ccfec148a522fbf5b8375245cbb3 + 1;
                    Ie81b8b84cc2795e2e92168bfa496ece4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie818c5ea3f3b879fded32e6cb06ca546 == I0aad448f6b0692670432efdd1b92d115 ) begin
                    Iadaaac832a1422494d4206edee770d63  <= I074386ff6a3d8d644f4b2501c69f26c7;
                    Ia6eb1062be96666c061e5fc1f830e1d3  <=  0;
                end else begin
                    Iadaaac832a1422494d4206edee770d63  <=  ~I074386ff6a3d8d644f4b2501c69f26c7 + 1;
                    Ia6eb1062be96666c061e5fc1f830e1d3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a67a175863091a52844aae6ad277da0 == Ia5a7e36b324b3a34be321ef63db22f50 ) begin
                    I905b0ec8983ba423798bbe8282728af8  <= I83b378e5534c553b57beb22c5178a3ce;
                    Ia0947c561ef360d78d0dae68baee6161  <=  0;
                end else begin
                    I905b0ec8983ba423798bbe8282728af8  <=  ~I83b378e5534c553b57beb22c5178a3ce + 1;
                    Ia0947c561ef360d78d0dae68baee6161  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a67a175863091a52844aae6ad277da0 == I01399ecad74618d26fea1ef278a3125f ) begin
                    Ic646b82fb6e3d0afb3a58c4e0d68f06c  <= I14f79d67f75af6a495d6eb2986210cda;
                    I3cd67e0abb8ff03aa1068dcb61aa3468  <=  0;
                end else begin
                    Ic646b82fb6e3d0afb3a58c4e0d68f06c  <=  ~I14f79d67f75af6a495d6eb2986210cda + 1;
                    I3cd67e0abb8ff03aa1068dcb61aa3468  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a67a175863091a52844aae6ad277da0 == Ia56986ae4171b36a362b170920663c44 ) begin
                    Ie57f41c62e23092974664f967a27566d  <= Iacd805413ec1eb001b3083554f187554;
                    Ic64779388389bf13a0e5240613caefc7  <=  0;
                end else begin
                    Ie57f41c62e23092974664f967a27566d  <=  ~Iacd805413ec1eb001b3083554f187554 + 1;
                    Ic64779388389bf13a0e5240613caefc7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a67a175863091a52844aae6ad277da0 == I7785a1b6345c7a2086b3d2a032970fa8 ) begin
                    I34524ca1dddbeadcc060954238175e7f  <= I3e61e09fcc81a0011a79f5c5ce77bc46;
                    I767cd611a030d15fc5eebc6e1b9ea2dc  <=  0;
                end else begin
                    I34524ca1dddbeadcc060954238175e7f  <=  ~I3e61e09fcc81a0011a79f5c5ce77bc46 + 1;
                    I767cd611a030d15fc5eebc6e1b9ea2dc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a67a175863091a52844aae6ad277da0 == I778c7251ca1b16e1ea1a4720ec7ba2de ) begin
                    Iaf2a93993f99814321951a6bffd8bdd4  <= I6e6cbb7dba8eb3c02b5b4e4469e23cea;
                    I03e14765645af77dd39ed51320bf7a95  <=  0;
                end else begin
                    Iaf2a93993f99814321951a6bffd8bdd4  <=  ~I6e6cbb7dba8eb3c02b5b4e4469e23cea + 1;
                    I03e14765645af77dd39ed51320bf7a95  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia3aba80aead67feab12e4800fef82322 == I1fcb2b0e5beab6a80ce06aeca85610b6 ) begin
                    I97e4f7a9a8a42be813c6e4128936df3f  <= I8b25822c33f7d506ef69216af3fdab44;
                    I29e966dc25c12cd095c25c5e6fd6d872  <=  0;
                end else begin
                    I97e4f7a9a8a42be813c6e4128936df3f  <=  ~I8b25822c33f7d506ef69216af3fdab44 + 1;
                    I29e966dc25c12cd095c25c5e6fd6d872  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia3aba80aead67feab12e4800fef82322 == I3f8184c2f7e604f0581e5c02f5b9563b ) begin
                    I682a67100f862bac0155a870cae0528c  <= I06fd642cbc8aa2f65197801d7459cfa2;
                    Ie8b68c8c51e2e03a3797a2ec3f8a56ae  <=  0;
                end else begin
                    I682a67100f862bac0155a870cae0528c  <=  ~I06fd642cbc8aa2f65197801d7459cfa2 + 1;
                    Ie8b68c8c51e2e03a3797a2ec3f8a56ae  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia3aba80aead67feab12e4800fef82322 == I25be48f72f47043fb6e8b7f774db1912 ) begin
                    Id5296b03b99bbf52d3ec04dddf3e84b1  <= I22202e6c3de9b06c04ce9514af28933e;
                    Ibbcfb7c284a2c99332d9261a4de199f1  <=  0;
                end else begin
                    Id5296b03b99bbf52d3ec04dddf3e84b1  <=  ~I22202e6c3de9b06c04ce9514af28933e + 1;
                    Ibbcfb7c284a2c99332d9261a4de199f1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia3aba80aead67feab12e4800fef82322 == If75d53ea58491447eb2344e993b4881e ) begin
                    Ibb089d47014f9002f2ea6b431156d9af  <= Ib991cdbb91133cb82e154c575e00a174;
                    I3e33a1f3e03bdb35d7c03f17f4ba4ebd  <=  0;
                end else begin
                    Ibb089d47014f9002f2ea6b431156d9af  <=  ~Ib991cdbb91133cb82e154c575e00a174 + 1;
                    I3e33a1f3e03bdb35d7c03f17f4ba4ebd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia3aba80aead67feab12e4800fef82322 == I4951621739ec145bcf3004b0f72e26db ) begin
                    I83496522139d35aa028dc9cb8a78d442  <= I5590364df6874420e169aa444ab520b9;
                    I0f81337862e31b6a4a6db462533d17f3  <=  0;
                end else begin
                    I83496522139d35aa028dc9cb8a78d442  <=  ~I5590364df6874420e169aa444ab520b9 + 1;
                    I0f81337862e31b6a4a6db462533d17f3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc == I959793f388e50197e4e31dae019d64f2 ) begin
                    Ifd4ca5a83fa0c09b043ad54d25971410  <= I43a9e393037fb4aa84741dca22648459;
                    I5029faffc78b92bc6e76d08fc4cd822f  <=  0;
                end else begin
                    Ifd4ca5a83fa0c09b043ad54d25971410  <=  ~I43a9e393037fb4aa84741dca22648459 + 1;
                    I5029faffc78b92bc6e76d08fc4cd822f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc == I8bccd3ff9583b2e33bf26d779f1c6233 ) begin
                    I6efbc715be55b616551a7d4650a446dd  <= Ibb4d8301d90c66fdfac92b3fbc53c019;
                    I11262f431003b344ab224ab5488995c2  <=  0;
                end else begin
                    I6efbc715be55b616551a7d4650a446dd  <=  ~Ibb4d8301d90c66fdfac92b3fbc53c019 + 1;
                    I11262f431003b344ab224ab5488995c2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc == I177f26189ade299e79c1406cc8171ae0 ) begin
                    I572bf74835f5acdf5a17de2063c293fc  <= Ibae217fa4b808e4accbeb8f4a9a976ab;
                    I3f0fc144d868b4446b6d261b3ac80a67  <=  0;
                end else begin
                    I572bf74835f5acdf5a17de2063c293fc  <=  ~Ibae217fa4b808e4accbeb8f4a9a976ab + 1;
                    I3f0fc144d868b4446b6d261b3ac80a67  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc == I93f3cd21e4819405b800ade59c9ccdd4 ) begin
                    I5f8194ef67d22bcd38f415fe8d9a6ce7  <= Ia8bd7a3594f7084a57e64da023bf784c;
                    I463736cac698d2366442abf5fba61580  <=  0;
                end else begin
                    I5f8194ef67d22bcd38f415fe8d9a6ce7  <=  ~Ia8bd7a3594f7084a57e64da023bf784c + 1;
                    I463736cac698d2366442abf5fba61580  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1181d42b560fca7bb5c924a81a5db1fc == Ie655403fd0fb16aaa04783a2ff742064 ) begin
                    I3d3f2dff1f64ce14071e5f315bb8a57f  <= I3ce4b9d41f5472bf60ed2802a2ab10eb;
                    I6cc14595c5c11f3ef8daa2a0b0634f73  <=  0;
                end else begin
                    I3d3f2dff1f64ce14071e5f315bb8a57f  <=  ~I3ce4b9d41f5472bf60ed2802a2ab10eb + 1;
                    I6cc14595c5c11f3ef8daa2a0b0634f73  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf == I1c3163e355c43d0a134c88fa671c41f3 ) begin
                    I8e3880fe0374bc068ed14eeff9f6d009  <= I93ec9bc6fbd056e7e52496546493e727;
                    Ia2345aaec32840b490d4b58c6ab3f115  <=  0;
                end else begin
                    I8e3880fe0374bc068ed14eeff9f6d009  <=  ~I93ec9bc6fbd056e7e52496546493e727 + 1;
                    Ia2345aaec32840b490d4b58c6ab3f115  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf == Ie378961bdb2de01ac733e765bba5eaa4 ) begin
                    I51d8f49653c7468b2923390dc5932a2a  <= I2374b90dde1cf481baa40af31e1a43e3;
                    Ifdca49a87cf807777f2e460bd3d3a4fb  <=  0;
                end else begin
                    I51d8f49653c7468b2923390dc5932a2a  <=  ~I2374b90dde1cf481baa40af31e1a43e3 + 1;
                    Ifdca49a87cf807777f2e460bd3d3a4fb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf == Ife404037f29f17b3edcc4d1334298781 ) begin
                    Ibeb380f8f935c8e061fe00734675662a  <= I0cee595f488a909ade8a3b4c90dbb0c7;
                    I4fab81c713b53f66f545f4f614713462  <=  0;
                end else begin
                    Ibeb380f8f935c8e061fe00734675662a  <=  ~I0cee595f488a909ade8a3b4c90dbb0c7 + 1;
                    I4fab81c713b53f66f545f4f614713462  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf == I4109fd0e3086c344f926c4a83b378296 ) begin
                    I641f4280286c9343b7ce001a8b43fa21  <= Iba4c3d91d492b000ab1de7add9f171a9;
                    I1dd4557e3f4df4fa18a9198f9f36a98c  <=  0;
                end else begin
                    I641f4280286c9343b7ce001a8b43fa21  <=  ~Iba4c3d91d492b000ab1de7add9f171a9 + 1;
                    I1dd4557e3f4df4fa18a9198f9f36a98c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie4e5f3d7c5d2df30653f5666d14567bf == I5d9e11667955d8128b76d9144463e59c ) begin
                    I796970d7c73d8fbd7d25793d0dbf9872  <= I2b4152aa4c51cc1c1ffabac78cea267c;
                    Id2ac1ca1ab4cb5eaba4ebb9dcb31d857  <=  0;
                end else begin
                    I796970d7c73d8fbd7d25793d0dbf9872  <=  ~I2b4152aa4c51cc1c1ffabac78cea267c + 1;
                    Id2ac1ca1ab4cb5eaba4ebb9dcb31d857  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifd9345cf219c58291c0b437aac093d78 == I70c06d2f51ef27666c8c39e0a13ff5cb ) begin
                    Ied0b1d10ae09c523d1cd1cd3e5b184c6  <= Ie4c3dd5c191aff00a6d62006223c2b76;
                    Id40872fc0d4f1e9ce25d366069af2f1a  <=  0;
                end else begin
                    Ied0b1d10ae09c523d1cd1cd3e5b184c6  <=  ~Ie4c3dd5c191aff00a6d62006223c2b76 + 1;
                    Id40872fc0d4f1e9ce25d366069af2f1a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifd9345cf219c58291c0b437aac093d78 == Iacd270f7fbb94c91757a4f8780616e1e ) begin
                    I7d0d39d94d929741158c39f69e8169e4  <= Ie4c0ba9510f9b924999bb5f432137271;
                    If3b1c8b7c2296e5664f105adc761fd48  <=  0;
                end else begin
                    I7d0d39d94d929741158c39f69e8169e4  <=  ~Ie4c0ba9510f9b924999bb5f432137271 + 1;
                    If3b1c8b7c2296e5664f105adc761fd48  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifd9345cf219c58291c0b437aac093d78 == Ia95e1a8c5bce4673824d56d6fab81f4b ) begin
                    I2349636f6ea8796c7b798aa555641a9e  <= I5bad544a17b384973d5672acbe0ac0d5;
                    Idd694db68c0f91155fd81a106d596d8c  <=  0;
                end else begin
                    I2349636f6ea8796c7b798aa555641a9e  <=  ~I5bad544a17b384973d5672acbe0ac0d5 + 1;
                    Idd694db68c0f91155fd81a106d596d8c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifd9345cf219c58291c0b437aac093d78 == I49137af52922e3872901905fd7c70601 ) begin
                    Ia3739201eb91605fc115bf320d4c24f0  <= I231bfb8e19e1d9c4bbd29a0bd75c1ed3;
                    I89473d1b100eb64c951e986819a4bc59  <=  0;
                end else begin
                    Ia3739201eb91605fc115bf320d4c24f0  <=  ~I231bfb8e19e1d9c4bbd29a0bd75c1ed3 + 1;
                    I89473d1b100eb64c951e986819a4bc59  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifd9345cf219c58291c0b437aac093d78 == I548d9239de9b536e1b581327961b53df ) begin
                    Ic74cc511acc98510da011e126edaf3a3  <= I1ecf87e33de04d02db9e64590bcaffde;
                    I4351f5987566977330a1e69b78d4e6aa  <=  0;
                end else begin
                    Ic74cc511acc98510da011e126edaf3a3  <=  ~I1ecf87e33de04d02db9e64590bcaffde + 1;
                    I4351f5987566977330a1e69b78d4e6aa  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 == Ifad4cf6d79d76caa33927ba4a6b94b45 ) begin
                    I89b1312c0696711956ddcf787e37f3c9  <= I60c97bf58193f004e3fcfdbd6a03ce6e;
                    Ic067d44971ef80f6c63c6e187a583e3e  <=  0;
                end else begin
                    I89b1312c0696711956ddcf787e37f3c9  <=  ~I60c97bf58193f004e3fcfdbd6a03ce6e + 1;
                    Ic067d44971ef80f6c63c6e187a583e3e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 == Ie78dd544469009d2b182d2b76694df6a ) begin
                    Ib2ef1187c1743da2cd83eb9231a7ddf1  <= Ib71065a3fe70d3ab5f05b0c393278631;
                    I9d46fd2fca52ea2ecb6242801a4378a3  <=  0;
                end else begin
                    Ib2ef1187c1743da2cd83eb9231a7ddf1  <=  ~Ib71065a3fe70d3ab5f05b0c393278631 + 1;
                    I9d46fd2fca52ea2ecb6242801a4378a3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 == I69122b791a8f717c501f2842240a51f6 ) begin
                    I21710bdb6874ab83e2b2a2cffb026ab8  <= I984074a5c77445ad266463e20d77899e;
                    I916104565afa11bfd9b3ef53551ade1d  <=  0;
                end else begin
                    I21710bdb6874ab83e2b2a2cffb026ab8  <=  ~I984074a5c77445ad266463e20d77899e + 1;
                    I916104565afa11bfd9b3ef53551ade1d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 == Ib89ed0cfe4ba481ae28b835d4248babf ) begin
                    I2ec8afd22c84596550412a5d2c7129af  <= I50bb40691aa09c42e0b64a076b50a971;
                    I48812dfaa796a851f23d230227be8969  <=  0;
                end else begin
                    I2ec8afd22c84596550412a5d2c7129af  <=  ~I50bb40691aa09c42e0b64a076b50a971 + 1;
                    I48812dfaa796a851f23d230227be8969  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4f2d7bb48918ce51efe6b3b12f9f8e65 == I6ec25bbba8c41ebdf4efa95fc1d8e1b0 ) begin
                    I57056cc2fd4bd1ea6e980cf90c22e871  <= I753bff437b6c563f5fddf19685405504;
                    Ia2d3db44f16c9bf381145ce71ba2efd2  <=  0;
                end else begin
                    I57056cc2fd4bd1ea6e980cf90c22e871  <=  ~I753bff437b6c563f5fddf19685405504 + 1;
                    Ia2d3db44f16c9bf381145ce71ba2efd2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifa612e6208151c616c3a0319182a96f1 == I92953d645060c118de19fafee18e34a1 ) begin
                    I233becd31032d63e65371119edb2cf79  <= I21f2ec69bcc507756e2a5f85d3ead3e8;
                    I849110a991c42aefaead8d9500a18912  <=  0;
                end else begin
                    I233becd31032d63e65371119edb2cf79  <=  ~I21f2ec69bcc507756e2a5f85d3ead3e8 + 1;
                    I849110a991c42aefaead8d9500a18912  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifa612e6208151c616c3a0319182a96f1 == Id89c23eca2ed6103c87dc296082605ab ) begin
                    I0142623400f5994f581a4797fd9d327c  <= Iddec4486996054e475499d370016a685;
                    Ic4988fc07458064e44f882807bd13c4b  <=  0;
                end else begin
                    I0142623400f5994f581a4797fd9d327c  <=  ~Iddec4486996054e475499d370016a685 + 1;
                    Ic4988fc07458064e44f882807bd13c4b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifa612e6208151c616c3a0319182a96f1 == I070e631601f2529f8f18ad0be6a70316 ) begin
                    Id3e298c9f2709d8dc01c18626ea846e8  <= I3d3edd06f8907f4369b825062348da87;
                    I0fdd344f1ce42003661bb06c2c0d2fb5  <=  0;
                end else begin
                    Id3e298c9f2709d8dc01c18626ea846e8  <=  ~I3d3edd06f8907f4369b825062348da87 + 1;
                    I0fdd344f1ce42003661bb06c2c0d2fb5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifa612e6208151c616c3a0319182a96f1 == Ie1e3e5fbe2e2ae4cb3218616bcaa0ae1 ) begin
                    I1044e090bdf84a1bd30438137d6ed056  <= I72467ef10ecced8395a6870a39525787;
                    Ib2ab217127041c49acfc86ef2eba3350  <=  0;
                end else begin
                    I1044e090bdf84a1bd30438137d6ed056  <=  ~I72467ef10ecced8395a6870a39525787 + 1;
                    Ib2ab217127041c49acfc86ef2eba3350  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifa612e6208151c616c3a0319182a96f1 == I6b2795593e93e47b2733c1e0003a7806 ) begin
                    Iff0f43c1fb40bdb3271a3a38d89f4d6d  <= I9b74b672f55e7bf7560ba4dd2d0c79fd;
                    I5d6dfd14a38b207a97ba02a357965d5e  <=  0;
                end else begin
                    Iff0f43c1fb40bdb3271a3a38d89f4d6d  <=  ~I9b74b672f55e7bf7560ba4dd2d0c79fd + 1;
                    I5d6dfd14a38b207a97ba02a357965d5e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9cb28a0cc6358610854c8f8d1dd3c707 == I467646a701c26d253f43251aceac9527 ) begin
                    Ibc71a0c3641097c144513810bc9a0a7c  <= I285b012d2fb5e2279a79cf8edca24ac8;
                    I963472efe41928bdcd4c87ae5d6d9781  <=  0;
                end else begin
                    Ibc71a0c3641097c144513810bc9a0a7c  <=  ~I285b012d2fb5e2279a79cf8edca24ac8 + 1;
                    I963472efe41928bdcd4c87ae5d6d9781  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9cb28a0cc6358610854c8f8d1dd3c707 == I280a8abed1540ebaf599c094a0a75797 ) begin
                    I6ef3b025eb065f833efe6daaab699efb  <= I8faf911a7d1ea8b0abe54f6688068ca0;
                    Id8cde19539c6cdf7186230e34b96dc15  <=  0;
                end else begin
                    I6ef3b025eb065f833efe6daaab699efb  <=  ~I8faf911a7d1ea8b0abe54f6688068ca0 + 1;
                    Id8cde19539c6cdf7186230e34b96dc15  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9cb28a0cc6358610854c8f8d1dd3c707 == If75560cad0cb26bd315f3711d1e9711d ) begin
                    If76152e9435e7300b19095a9b070e0f4  <= I3dca974bf2d5631a47ebf8b945efab20;
                    Ia31ee8ac9735d3bd38298fd5d9812aa1  <=  0;
                end else begin
                    If76152e9435e7300b19095a9b070e0f4  <=  ~I3dca974bf2d5631a47ebf8b945efab20 + 1;
                    Ia31ee8ac9735d3bd38298fd5d9812aa1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9cb28a0cc6358610854c8f8d1dd3c707 == Id0d79e0b7361bae1b007c8a7d606f6fb ) begin
                    I5fa63303ab85db9c8cd268528eb604ca  <= I12141c45d147b058a9e392f3b7d7d06e;
                    I79bced0e80e2554a4e748644c5985896  <=  0;
                end else begin
                    I5fa63303ab85db9c8cd268528eb604ca  <=  ~I12141c45d147b058a9e392f3b7d7d06e + 1;
                    I79bced0e80e2554a4e748644c5985896  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40bcc924f5cf1f7d587aa35267022261 == Iac7bb2fe5935b53852a63923c53f13a1 ) begin
                    I69d6adcd3d35a24b393e97ed6a99c061  <= Ia527c96e30b782f837bc6206961400e4;
                    Id0216555323efdec39d0448568f59f23  <=  0;
                end else begin
                    I69d6adcd3d35a24b393e97ed6a99c061  <=  ~Ia527c96e30b782f837bc6206961400e4 + 1;
                    Id0216555323efdec39d0448568f59f23  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40bcc924f5cf1f7d587aa35267022261 == I4554a553586d9966e7d4e8d99a5c799d ) begin
                    I8980eca0e5973840121576b6eaaab736  <= I6adbdb64422a08be9bf9e538db97463b;
                    I35c6735d2fa06f57341b6010f5bb825d  <=  0;
                end else begin
                    I8980eca0e5973840121576b6eaaab736  <=  ~I6adbdb64422a08be9bf9e538db97463b + 1;
                    I35c6735d2fa06f57341b6010f5bb825d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40bcc924f5cf1f7d587aa35267022261 == I84a85d995e807610f153e72ea3df3ae0 ) begin
                    Iadbb5c4f7b7c02e151d5118a7ede1f0b  <= I958cdf5367c7b0bd58b70b763d3af8aa;
                    Id2e8b17327e8c85999d3d6b3dd31a164  <=  0;
                end else begin
                    Iadbb5c4f7b7c02e151d5118a7ede1f0b  <=  ~I958cdf5367c7b0bd58b70b763d3af8aa + 1;
                    Id2e8b17327e8c85999d3d6b3dd31a164  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40bcc924f5cf1f7d587aa35267022261 == Ic68f898ba0d0073df41bbfae0944c9de ) begin
                    Ifff90bff22a3bcc33261004136d2e655  <= I91b7b8e8887b5dd9853297463c55b78d;
                    Iccd9ca809045617acea3364a6c86fde9  <=  0;
                end else begin
                    Ifff90bff22a3bcc33261004136d2e655  <=  ~I91b7b8e8887b5dd9853297463c55b78d + 1;
                    Iccd9ca809045617acea3364a6c86fde9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5238f7273b05b8b9f376314acdc6cc42 == Iab98e00ea4dca63c81eb8f78a133b1bd ) begin
                    I8d13628f322640414a4b556ee48d3bdd  <= I6162978f0c57958ad0403246fb0530dd;
                    I8ce27f01f84ea9babfca8074bb57417a  <=  0;
                end else begin
                    I8d13628f322640414a4b556ee48d3bdd  <=  ~I6162978f0c57958ad0403246fb0530dd + 1;
                    I8ce27f01f84ea9babfca8074bb57417a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5238f7273b05b8b9f376314acdc6cc42 == I67aca5b07f66a9f3e8a5550020802c63 ) begin
                    If7d187cc56b1014b1582c5f5b94759f1  <= I508142e70fd04513977130556aa574ef;
                    If6bad1b3865cb4cec97a730043863b3d  <=  0;
                end else begin
                    If7d187cc56b1014b1582c5f5b94759f1  <=  ~I508142e70fd04513977130556aa574ef + 1;
                    If6bad1b3865cb4cec97a730043863b3d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5238f7273b05b8b9f376314acdc6cc42 == Id4b0e0110bcd34cf8f0a9a92108b88c2 ) begin
                    Ia01d5a33078abf4b2d6c625af01c25f6  <= I2afab673e4b803ffd888f187de47fa49;
                    I0c88089ad1c5fc9928c091c1c677ca66  <=  0;
                end else begin
                    Ia01d5a33078abf4b2d6c625af01c25f6  <=  ~I2afab673e4b803ffd888f187de47fa49 + 1;
                    I0c88089ad1c5fc9928c091c1c677ca66  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5238f7273b05b8b9f376314acdc6cc42 == I29ee6514004941d4280cf4a93e7baf5d ) begin
                    I4c74240688b5635b5323ce3a8ac666fb  <= I7a56f81596920126a9ea2c9fb3a19285;
                    Ida2ed38c156200b9511c3b4515f42e5e  <=  0;
                end else begin
                    I4c74240688b5635b5323ce3a8ac666fb  <=  ~I7a56f81596920126a9ea2c9fb3a19285 + 1;
                    Ida2ed38c156200b9511c3b4515f42e5e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7137f56eeb4c4ae08bbc238db4cd3441 == I3bb0ea6e5c41271be14ed45d4b8ece5b ) begin
                    I943e9afa0dc80fb50b5869cf34726823  <= Ic6252de2c819f2243476ddf82e22d137;
                    Id322e4a2b0197e5b0f67a220134ca540  <=  0;
                end else begin
                    I943e9afa0dc80fb50b5869cf34726823  <=  ~Ic6252de2c819f2243476ddf82e22d137 + 1;
                    Id322e4a2b0197e5b0f67a220134ca540  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7137f56eeb4c4ae08bbc238db4cd3441 == I0a1dc75c36d5fb043c80dde4e8c5e577 ) begin
                    I44d8779f30245bc7f1475e6feb762cec  <= Ieea8672b2f23711c6ba893de5c5d8bc2;
                    I935862d2f7c82e05768f55434167ba47  <=  0;
                end else begin
                    I44d8779f30245bc7f1475e6feb762cec  <=  ~Ieea8672b2f23711c6ba893de5c5d8bc2 + 1;
                    I935862d2f7c82e05768f55434167ba47  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7137f56eeb4c4ae08bbc238db4cd3441 == I89e39167f230c52eaf64e8c5ce8fc38d ) begin
                    I479e7456c445ad604ebc134872a0fbfa  <= I3a4dbdf517b8f9c93b567f91870e6160;
                    I1c6dd243cd7d2b8d00eb59e2ae30331c  <=  0;
                end else begin
                    I479e7456c445ad604ebc134872a0fbfa  <=  ~I3a4dbdf517b8f9c93b567f91870e6160 + 1;
                    I1c6dd243cd7d2b8d00eb59e2ae30331c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7137f56eeb4c4ae08bbc238db4cd3441 == Id6e88b1c05e5f4e7188f4b646f428b55 ) begin
                    I484f372e3a2e74e0791b06aa666b781e  <= I4731ee7a0e08c69e2bd2a8bcea0838c2;
                    I8ab7b4e7f78fa63ec77224c7e5a31198  <=  0;
                end else begin
                    I484f372e3a2e74e0791b06aa666b781e  <=  ~I4731ee7a0e08c69e2bd2a8bcea0838c2 + 1;
                    I8ab7b4e7f78fa63ec77224c7e5a31198  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I02335be013799e2560a98b6a82a0c528 == Id9b024743e4060a62c6dde2646b5c998 ) begin
                    I64b07241996c48963595f28e35a75be5  <= I1b6cbbcf01a65cd1c2f1e241f849c904;
                    If20d6cdf73bb1a925317f35de01b6f62  <=  0;
                end else begin
                    I64b07241996c48963595f28e35a75be5  <=  ~I1b6cbbcf01a65cd1c2f1e241f849c904 + 1;
                    If20d6cdf73bb1a925317f35de01b6f62  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I02335be013799e2560a98b6a82a0c528 == I2bc4cf6682dca441749b95f63592dd8e ) begin
                    Idf678798bf4e1cd316a49a2b413cb29f  <= I663aee79f824c854f57c19e87207529b;
                    I8c2bc7a3c5c7e798a9dbd0199d37bfd5  <=  0;
                end else begin
                    Idf678798bf4e1cd316a49a2b413cb29f  <=  ~I663aee79f824c854f57c19e87207529b + 1;
                    I8c2bc7a3c5c7e798a9dbd0199d37bfd5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I02335be013799e2560a98b6a82a0c528 == I05d8735777c75ecc9f1e5d2f972f5c21 ) begin
                    I35fd5e5e93f992ef5ff6b11f9d69609c  <= I34ff7299c9d83affa4512b7da302c199;
                    If814b033c7e3229ba1475b305fe98307  <=  0;
                end else begin
                    I35fd5e5e93f992ef5ff6b11f9d69609c  <=  ~I34ff7299c9d83affa4512b7da302c199 + 1;
                    If814b033c7e3229ba1475b305fe98307  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I02335be013799e2560a98b6a82a0c528 == Iaa201a0537ab3cbcb5bc065871e0153b ) begin
                    Ie72397edc1c597c0a8213b67a030a482  <= I70ca6c9d0a5c99e0036479f7b5dd760a;
                    I6e69f6d33a933441458f5a46decc4e8d  <=  0;
                end else begin
                    Ie72397edc1c597c0a8213b67a030a482  <=  ~I70ca6c9d0a5c99e0036479f7b5dd760a + 1;
                    I6e69f6d33a933441458f5a46decc4e8d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I02335be013799e2560a98b6a82a0c528 == Ib76deffcb8cd38d5643df9447f3b060b ) begin
                    Iae50178e99a07cee0eea6f7cfdcedf1f  <= I835bb7345787eaadc41816858e0a71a1;
                    Ie2bb4ef41cf43cbea46b7a6d492bf03b  <=  0;
                end else begin
                    Iae50178e99a07cee0eea6f7cfdcedf1f  <=  ~I835bb7345787eaadc41816858e0a71a1 + 1;
                    Ie2bb4ef41cf43cbea46b7a6d492bf03b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id327bb65156c8307901dfcb4184bb65f == I6483a59c7f2bc77b445b202f0448eb2a ) begin
                    Idd7082c7a65d7f8e0ea88142312a631e  <= I3c7f6fdd0e9cc7426df76027912d1ccb;
                    I757b0e2104a4d9913cf6b3a13ad7d6d6  <=  0;
                end else begin
                    Idd7082c7a65d7f8e0ea88142312a631e  <=  ~I3c7f6fdd0e9cc7426df76027912d1ccb + 1;
                    I757b0e2104a4d9913cf6b3a13ad7d6d6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id327bb65156c8307901dfcb4184bb65f == Ic1ffdfe961dc8458b1d4cb36642a386a ) begin
                    I4b580dc4cfac9e9315d03b60e2a915d9  <= I9ff512085174a7720705d0fb37c4ec34;
                    I46c7f4a6ef4b3ac3eb74b4ba2552fcdd  <=  0;
                end else begin
                    I4b580dc4cfac9e9315d03b60e2a915d9  <=  ~I9ff512085174a7720705d0fb37c4ec34 + 1;
                    I46c7f4a6ef4b3ac3eb74b4ba2552fcdd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id327bb65156c8307901dfcb4184bb65f == I0fb493a1f8f2810ddf67a6cbcb2c782c ) begin
                    I77cdc9841414221c3f6c3cf35397059f  <= I6a69cdf2bae1ea68c9be56dcc4e76a59;
                    I247479fee56f209f758feeb4770e50de  <=  0;
                end else begin
                    I77cdc9841414221c3f6c3cf35397059f  <=  ~I6a69cdf2bae1ea68c9be56dcc4e76a59 + 1;
                    I247479fee56f209f758feeb4770e50de  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id327bb65156c8307901dfcb4184bb65f == I2c555af9585a50d2cd6a27c223c8722c ) begin
                    Ie59619c3e78e616e1febd2db2fa940ae  <= I855ddead34ac131137ba644afbfea2b7;
                    I2ada4b104b94c163f3d9201808d21121  <=  0;
                end else begin
                    Ie59619c3e78e616e1febd2db2fa940ae  <=  ~I855ddead34ac131137ba644afbfea2b7 + 1;
                    I2ada4b104b94c163f3d9201808d21121  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id327bb65156c8307901dfcb4184bb65f == I5f93af2953a9f1aea5cf55a037f7af6e ) begin
                    I5bc8079a5896f59bc6137b59c4b7e750  <= Ib1a463388daf270eb0ce698d7b5ded4b;
                    Ic7f0721d5160d4ce266b21c53aad0b4e  <=  0;
                end else begin
                    I5bc8079a5896f59bc6137b59c4b7e750  <=  ~Ib1a463388daf270eb0ce698d7b5ded4b + 1;
                    Ic7f0721d5160d4ce266b21c53aad0b4e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56331cb7b310613016958553732cdf40 == I25b3e2b9f55ea811784ba8ad8c5f516d ) begin
                    I239bf978d991f702ad23bc6b4b8be1dc  <= I74e4bb7530c02073f9b15a6389659d4b;
                    I9af70dd16bd606c4b9588ce32ce9844d  <=  0;
                end else begin
                    I239bf978d991f702ad23bc6b4b8be1dc  <=  ~I74e4bb7530c02073f9b15a6389659d4b + 1;
                    I9af70dd16bd606c4b9588ce32ce9844d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56331cb7b310613016958553732cdf40 == I93fb55e460d75b8d36c19833849bc1d2 ) begin
                    I450351fbb31246b49cfb2d622b9e90b4  <= I6721b13abeddc76139bdc7380434cc2a;
                    I30c5fca5bab3bc9cf5c024c3302bbdbd  <=  0;
                end else begin
                    I450351fbb31246b49cfb2d622b9e90b4  <=  ~I6721b13abeddc76139bdc7380434cc2a + 1;
                    I30c5fca5bab3bc9cf5c024c3302bbdbd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56331cb7b310613016958553732cdf40 == Ic51082943371a401c48202b4e655e84c ) begin
                    Ia7c17a0979f3bbb9e9e821bf69a239b7  <= I84fba239c5705bcd92096e204cc9438c;
                    I09db79951c2115c2db0a3036bcb2b63f  <=  0;
                end else begin
                    Ia7c17a0979f3bbb9e9e821bf69a239b7  <=  ~I84fba239c5705bcd92096e204cc9438c + 1;
                    I09db79951c2115c2db0a3036bcb2b63f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56331cb7b310613016958553732cdf40 == Ib53122ae54dc4ac5b090ba8aa3ab9959 ) begin
                    Ic22975c34b92a39bc8940076e80d3c0b  <= I4d46e4d50176768fda897949545e2125;
                    Id76636b29db2c1a69d585b68731fc3b0  <=  0;
                end else begin
                    Ic22975c34b92a39bc8940076e80d3c0b  <=  ~I4d46e4d50176768fda897949545e2125 + 1;
                    Id76636b29db2c1a69d585b68731fc3b0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56331cb7b310613016958553732cdf40 == I459abcd025ce92565cbbfaada735a325 ) begin
                    Ia7be8cf38ecee4568a939cb2ef727619  <= I57086cfab3b163c3911c3cf7bfb3141a;
                    I2ce42f5733f4d0cf15d1a7944fe0344f  <=  0;
                end else begin
                    Ia7be8cf38ecee4568a939cb2ef727619  <=  ~I57086cfab3b163c3911c3cf7bfb3141a + 1;
                    I2ce42f5733f4d0cf15d1a7944fe0344f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 == If8abbbaf2986196395e63aa49b1022bb ) begin
                    I3e475cb1733d494f5f7c4b26a07d5852  <= Ice174debd5dc911fdf5d5756cff8d731;
                    I87e7191f5ec3f0847afbca81660a7608  <=  0;
                end else begin
                    I3e475cb1733d494f5f7c4b26a07d5852  <=  ~Ice174debd5dc911fdf5d5756cff8d731 + 1;
                    I87e7191f5ec3f0847afbca81660a7608  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 == I830ffb778558295001c003f114b66198 ) begin
                    Ib2c0df16678f6aac19f7af4ad4e53ef8  <= Ie369670edc5b602d305904f3a4a4381f;
                    I0f8f4304c88efcc90c021be7764be01b  <=  0;
                end else begin
                    Ib2c0df16678f6aac19f7af4ad4e53ef8  <=  ~Ie369670edc5b602d305904f3a4a4381f + 1;
                    I0f8f4304c88efcc90c021be7764be01b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 == I56e732494aa029b716ac04289d951e27 ) begin
                    I8bd2ef39eeb7089409db02e3806956ac  <= I41f66f79339962ef42fab3b88e571170;
                    Ie8b6b834bdde210d6f7a3e60fc78275d  <=  0;
                end else begin
                    I8bd2ef39eeb7089409db02e3806956ac  <=  ~I41f66f79339962ef42fab3b88e571170 + 1;
                    Ie8b6b834bdde210d6f7a3e60fc78275d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 == Id077045b00947ff1b4de86777d84a48f ) begin
                    Ie3669e34cd19462f524932b3d232b546  <= I5cbd2fad4d90bd77ba3d2448a37ac60f;
                    I591b99ab1b55e2eb4c10996efab5e0d0  <=  0;
                end else begin
                    Ie3669e34cd19462f524932b3d232b546  <=  ~I5cbd2fad4d90bd77ba3d2448a37ac60f + 1;
                    I591b99ab1b55e2eb4c10996efab5e0d0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3b00960f8af88a5aba7a2104dfca9a7 == I7ce7ba4f90dea6eb91d61cb456134df3 ) begin
                    I1ecea23a4e56948365dcb04c5bf6d6d6  <= Id86a2869148e2885633d9e277f7041c3;
                    I27402f7d7892626f9b5ea1fc39987c23  <=  0;
                end else begin
                    I1ecea23a4e56948365dcb04c5bf6d6d6  <=  ~Id86a2869148e2885633d9e277f7041c3 + 1;
                    I27402f7d7892626f9b5ea1fc39987c23  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 == Iaee8dd8470306340982baafd8c9e28b5 ) begin
                    Iac222e9e39e300d7161ed05153cd9ca0  <= Ifb7b585189db23efabfb522c9b45bede;
                    Ie6e9475310530f511d38602f2c58a28f  <=  0;
                end else begin
                    Iac222e9e39e300d7161ed05153cd9ca0  <=  ~Ifb7b585189db23efabfb522c9b45bede + 1;
                    Ie6e9475310530f511d38602f2c58a28f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 == I35088305c303ace3b0bd194f5efa557f ) begin
                    I292683f8453be58f65370a286c1a4505  <= I7763f0d28d8065d8c94ef8df96b2ab06;
                    I30eeb2d396c381acb08253d886025fe1  <=  0;
                end else begin
                    I292683f8453be58f65370a286c1a4505  <=  ~I7763f0d28d8065d8c94ef8df96b2ab06 + 1;
                    I30eeb2d396c381acb08253d886025fe1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 == If28f074339d099d0c8f0e582c11f57e8 ) begin
                    I1dff7459553fccefc94a6020cc248a49  <= I115ba88588187c7115977e95bd26ee5a;
                    I9a9a3b834bb25862cbe40375e20c2163  <=  0;
                end else begin
                    I1dff7459553fccefc94a6020cc248a49  <=  ~I115ba88588187c7115977e95bd26ee5a + 1;
                    I9a9a3b834bb25862cbe40375e20c2163  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 == I55b6efd25a905ab958ff62e0334d0116 ) begin
                    I9acec7aa4b420b7c820028b669a8bfb4  <= I6e7f2bdd0c8231a3689893ef4877fdba;
                    I1152ba49a018ec527bb8091c0cebd737  <=  0;
                end else begin
                    I9acec7aa4b420b7c820028b669a8bfb4  <=  ~I6e7f2bdd0c8231a3689893ef4877fdba + 1;
                    I1152ba49a018ec527bb8091c0cebd737  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7d1ef47f35b7a4c3ea2e4383732de398 == I859a2864cbe2fffc01b411e7b0a2c3d0 ) begin
                    I714b7d8b39c4135183b605dd97ff15d6  <= I546c513d5357ac1a6fe669888dfaf717;
                    I1cf3b72b3aa02961788688172c1ad2b2  <=  0;
                end else begin
                    I714b7d8b39c4135183b605dd97ff15d6  <=  ~I546c513d5357ac1a6fe669888dfaf717 + 1;
                    I1cf3b72b3aa02961788688172c1ad2b2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a == I3ede6ae83cec11aecdb308142c26f6d6 ) begin
                    Ie5856c36d9a310f890ecc5220590fc3e  <= Ib3e12c614471912d0b276cb9f0382b1b;
                    I09293a7f47ffb53331aad25a876d2562  <=  0;
                end else begin
                    Ie5856c36d9a310f890ecc5220590fc3e  <=  ~Ib3e12c614471912d0b276cb9f0382b1b + 1;
                    I09293a7f47ffb53331aad25a876d2562  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a == Icb7fa4f4271f536afd96934a45bbf0ff ) begin
                    I062b1d8d3b6fe6d8e158ede1f0af9eed  <= I7187a2499e3319da90b6d6fc64411b46;
                    Ic00d9c70df8f473695a4aa76827ef690  <=  0;
                end else begin
                    I062b1d8d3b6fe6d8e158ede1f0af9eed  <=  ~I7187a2499e3319da90b6d6fc64411b46 + 1;
                    Ic00d9c70df8f473695a4aa76827ef690  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a == I4dfd9e0bf539f3077f2d5a8bd3b5e469 ) begin
                    I0fbd5b5eef6da9adaf918390f6bdbc27  <= I9b46582473bb4dd5541a35ac708486f4;
                    I36132477ed96c4731e46d24e9ca1e9e8  <=  0;
                end else begin
                    I0fbd5b5eef6da9adaf918390f6bdbc27  <=  ~I9b46582473bb4dd5541a35ac708486f4 + 1;
                    I36132477ed96c4731e46d24e9ca1e9e8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a == I795091257b4f78363310623b731b347e ) begin
                    I73fb14b30841cf67e96ba329fdfa3e35  <= I929796fe327ee9c8a05e6bb683ae5d7c;
                    I2cb80c174e5ddbbaca6eabbfa7c669c7  <=  0;
                end else begin
                    I73fb14b30841cf67e96ba329fdfa3e35  <=  ~I929796fe327ee9c8a05e6bb683ae5d7c + 1;
                    I2cb80c174e5ddbbaca6eabbfa7c669c7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ibb013f036fc42687a04bdcbe2d0bbd8a == I6ff1f76a6ad568b5fa0cb300a67ceea9 ) begin
                    I6d6cfca51988c5ac32471fe8f4399bbc  <= Ib6638da8b69373c2026d3f5305825cde;
                    I359e17e055d03931cac7b41c77be575b  <=  0;
                end else begin
                    I6d6cfca51988c5ac32471fe8f4399bbc  <=  ~Ib6638da8b69373c2026d3f5305825cde + 1;
                    I359e17e055d03931cac7b41c77be575b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc == I5864383518b7c9a70f69b0fd1a64d4aa ) begin
                    Id7940e4951c96c3de9f45119043fbffd  <= I28c26bf4cf9693d1807818b2ca7883ac;
                    If466ac9d4d278b49b4aa91650b30ec2e  <=  0;
                end else begin
                    Id7940e4951c96c3de9f45119043fbffd  <=  ~I28c26bf4cf9693d1807818b2ca7883ac + 1;
                    If466ac9d4d278b49b4aa91650b30ec2e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc == I30959187f5ac883ab77af90ccfce5704 ) begin
                    Iea71361c5f846419eaa18ae4b9463ee8  <= I291fc4eef4b80d1020c96488b869727e;
                    I17d171b83e60410ce78a7e4fa9d17001  <=  0;
                end else begin
                    Iea71361c5f846419eaa18ae4b9463ee8  <=  ~I291fc4eef4b80d1020c96488b869727e + 1;
                    I17d171b83e60410ce78a7e4fa9d17001  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc == I0d2bcd2e24e64ad5703a580ddc415f3a ) begin
                    Ib67ac5fdd6e068ee799965b51aa893ba  <= I53006ed50f6211439681aa7659647e35;
                    Id79a4b98545d81fef573054b93ae80d4  <=  0;
                end else begin
                    Ib67ac5fdd6e068ee799965b51aa893ba  <=  ~I53006ed50f6211439681aa7659647e35 + 1;
                    Id79a4b98545d81fef573054b93ae80d4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc == I4d1ef379c32f93cdd18e2415ba83a5ea ) begin
                    I0bd84509dde112f3657bd5a12a8df72c  <= I47fe32973727237ae0cd4c306c7efbfb;
                    I4e8f5e83e32143008d70a8edf17e2ff5  <=  0;
                end else begin
                    I0bd84509dde112f3657bd5a12a8df72c  <=  ~I47fe32973727237ae0cd4c306c7efbfb + 1;
                    I4e8f5e83e32143008d70a8edf17e2ff5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I77eae49d321f1d1e39dd7c75829aaedc == I921c8abbe15effa3769c5c3f81427274 ) begin
                    I2caf86026460a024f752fa71b44f743f  <= Ic3e0c7d71f13a56a9a63e158c7f2cfa8;
                    I57cf1069290a2a5f30b75eb592752b88  <=  0;
                end else begin
                    I2caf86026460a024f752fa71b44f743f  <=  ~Ic3e0c7d71f13a56a9a63e158c7f2cfa8 + 1;
                    I57cf1069290a2a5f30b75eb592752b88  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 == I40cce0292c07026fb144dc28ba228485 ) begin
                    Id81d9c9ffa81c2653dea2e872ab2f71c  <= If383f241447cbea4e18f4f79fcdbf144;
                    I7447d4584dccf4dac9f0d359748ae327  <=  0;
                end else begin
                    Id81d9c9ffa81c2653dea2e872ab2f71c  <=  ~If383f241447cbea4e18f4f79fcdbf144 + 1;
                    I7447d4584dccf4dac9f0d359748ae327  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 == Ia1401fc86b9d014a28f1c5bfa7aefc2d ) begin
                    I0b4d1a08307d452870c3e762bd038568  <= Ia05354d3b4f61299d5897832639df2c2;
                    Ic4571481454a10eb7f8c0b58f9d35178  <=  0;
                end else begin
                    I0b4d1a08307d452870c3e762bd038568  <=  ~Ia05354d3b4f61299d5897832639df2c2 + 1;
                    Ic4571481454a10eb7f8c0b58f9d35178  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 == Id3899a9a35b467c103ed0dfef20dd4a1 ) begin
                    Id75cc40233cc8648e21a750d882d5ed4  <= I9faec40665477e8b3237773d606af2f0;
                    I00810b2849a3d3097e028efac18c0a06  <=  0;
                end else begin
                    Id75cc40233cc8648e21a750d882d5ed4  <=  ~I9faec40665477e8b3237773d606af2f0 + 1;
                    I00810b2849a3d3097e028efac18c0a06  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 == Icff78887751d68045a0bc21e69047c79 ) begin
                    I3ea9815ba887e373a0a477654f136856  <= Id231ab3133d4bed02aad7e5f560ee5f0;
                    I19be1cf97631f5bd782d8358fb55954b  <=  0;
                end else begin
                    I3ea9815ba887e373a0a477654f136856  <=  ~Id231ab3133d4bed02aad7e5f560ee5f0 + 1;
                    I19be1cf97631f5bd782d8358fb55954b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I420a4d69a077dc1996ddb4b715d63e15 == I9a2e36db1aa972536df63a24462eba98 ) begin
                    I8b26e270c3ca5563da39e7092ef830dc  <= I13616c8c7be221cf4d2c13ae87c38bed;
                    Id7fe36cc9d5c1d7cc54ee1040e6578de  <=  0;
                end else begin
                    I8b26e270c3ca5563da39e7092ef830dc  <=  ~I13616c8c7be221cf4d2c13ae87c38bed + 1;
                    Id7fe36cc9d5c1d7cc54ee1040e6578de  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I652202a4dc8f102d29334b4811f5628d == Id74033401d8494d013fcfd1f69537592 ) begin
                    Ib03f94d7e5ff830d5063cd514e7f7998  <= I8793bc728a4d423fb96a88c83bb9746f;
                    If6984aadfa0583c3281a04ba48f3d765  <=  0;
                end else begin
                    Ib03f94d7e5ff830d5063cd514e7f7998  <=  ~I8793bc728a4d423fb96a88c83bb9746f + 1;
                    If6984aadfa0583c3281a04ba48f3d765  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I652202a4dc8f102d29334b4811f5628d == Ib64741c15a5f128b008851c36d55c0ca ) begin
                    I00b05bb0b225b27562d6629725ac2126  <= I2fb6af0f152232550a3cadd55656df20;
                    Ia7750161c32ac0507e1ff6a8fe896148  <=  0;
                end else begin
                    I00b05bb0b225b27562d6629725ac2126  <=  ~I2fb6af0f152232550a3cadd55656df20 + 1;
                    Ia7750161c32ac0507e1ff6a8fe896148  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I652202a4dc8f102d29334b4811f5628d == Ie75e57f87e9c8cc7d29519f0419f1b22 ) begin
                    I1f273682cac5644f1fcc30ffa20f8cd8  <= I5144918fcd4ce1a061644240730fc52a;
                    I97d6084735a682ba654fc70a9e07f27d  <=  0;
                end else begin
                    I1f273682cac5644f1fcc30ffa20f8cd8  <=  ~I5144918fcd4ce1a061644240730fc52a + 1;
                    I97d6084735a682ba654fc70a9e07f27d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I652202a4dc8f102d29334b4811f5628d == I95bc08d218c4a924f810b69c7e2b923f ) begin
                    I483725645504999df82a4d0660873c1d  <= I1821eb21cdf8208ff6c2f28d963f7bd6;
                    I3e9d85c0ca08314fe2da0fa6977942b7  <=  0;
                end else begin
                    I483725645504999df82a4d0660873c1d  <=  ~I1821eb21cdf8208ff6c2f28d963f7bd6 + 1;
                    I3e9d85c0ca08314fe2da0fa6977942b7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0e33e0cdf39fc4cc99f6696e9f2784de == I6dd9a12bbad2fd4aded0354fbb09c6cb ) begin
                    I689dc18b56442b8db01bd7ca4c44d615  <= I80471575b1d4b69ef073056f798394ea;
                    Id28d0dd03217797390811bdd3564191b  <=  0;
                end else begin
                    I689dc18b56442b8db01bd7ca4c44d615  <=  ~I80471575b1d4b69ef073056f798394ea + 1;
                    Id28d0dd03217797390811bdd3564191b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0e33e0cdf39fc4cc99f6696e9f2784de == Ie78ca77c4a9cfac31f52cc1f49e5c6d1 ) begin
                    I805d665f394ff24f230bebfa6d252122  <= I890bf9b72cc3c71351547178d72796e5;
                    I0eb20560e7e211b67cfa8ca9e056c1da  <=  0;
                end else begin
                    I805d665f394ff24f230bebfa6d252122  <=  ~I890bf9b72cc3c71351547178d72796e5 + 1;
                    I0eb20560e7e211b67cfa8ca9e056c1da  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0e33e0cdf39fc4cc99f6696e9f2784de == I771cf2bb35d06a6009955936e2530f07 ) begin
                    Icfba3f165f1cdf2e6070239100e9ac3d  <= Icc9d28b84fa91028ae96cc9b8bae7555;
                    Id089d9523253f91c670099157325af05  <=  0;
                end else begin
                    Icfba3f165f1cdf2e6070239100e9ac3d  <=  ~Icc9d28b84fa91028ae96cc9b8bae7555 + 1;
                    Id089d9523253f91c670099157325af05  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0e33e0cdf39fc4cc99f6696e9f2784de == I2d9d14b5c585e74db793171f304e5d61 ) begin
                    I93c51f71db0e3df7f6e2978fd93fbb54  <= I0b0d167c415f8c14594bd61907d46d80;
                    I4db3f0e5ff2cc72e499ab5f1b9fd1d14  <=  0;
                end else begin
                    I93c51f71db0e3df7f6e2978fd93fbb54  <=  ~I0b0d167c415f8c14594bd61907d46d80 + 1;
                    I4db3f0e5ff2cc72e499ab5f1b9fd1d14  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib9479328689dec62f900946e56ba0eb4 == I1e7165374d01b2b7abb1e1883daa4463 ) begin
                    Ib7410e44d23eea21613074695b64bd2b  <= I9577d49a74520355e53a1818f479db0e;
                    I082972cc68873126a258e9db29e524f9  <=  0;
                end else begin
                    Ib7410e44d23eea21613074695b64bd2b  <=  ~I9577d49a74520355e53a1818f479db0e + 1;
                    I082972cc68873126a258e9db29e524f9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib9479328689dec62f900946e56ba0eb4 == I783fdf0d5058b09d9d0d5c87d9926c50 ) begin
                    I93cc273684a376d76a2e3468b3dc8bd7  <= Ie6e888d582ba9e600e91b119e2804642;
                    I3ba1cbc9ff352842d6d687b2218b6c0f  <=  0;
                end else begin
                    I93cc273684a376d76a2e3468b3dc8bd7  <=  ~Ie6e888d582ba9e600e91b119e2804642 + 1;
                    I3ba1cbc9ff352842d6d687b2218b6c0f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib9479328689dec62f900946e56ba0eb4 == I1c66ca0e94ab96e8420e97641a5a707b ) begin
                    Id133dc3fa65840136b1157fe97a1e962  <= Iccfac3d489b4b110d6b6e005a5ba45d8;
                    Id8fbc7f9a403b07efd27c20d6d78e661  <=  0;
                end else begin
                    Id133dc3fa65840136b1157fe97a1e962  <=  ~Iccfac3d489b4b110d6b6e005a5ba45d8 + 1;
                    Id8fbc7f9a403b07efd27c20d6d78e661  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib9479328689dec62f900946e56ba0eb4 == If5f2d3751eb3af97e20c680475976bb6 ) begin
                    Ib792104b6cf946d632f7591f2cd5e104  <= I69a67481ca8fd01dc5400dbe887b4f83;
                    I0628944b437e239b25736381fa59901d  <=  0;
                end else begin
                    Ib792104b6cf946d632f7591f2cd5e104  <=  ~I69a67481ca8fd01dc5400dbe887b4f83 + 1;
                    I0628944b437e239b25736381fa59901d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2728682c0f749d1a9e8afeacdf44bfb7 == I96f91ace9649929071ca3e6e87eda861 ) begin
                    Ia44bcc8308360d3e6fa351bc108df3fa  <= I1f36f045becec7f0528f4a935d3da2ff;
                    Icf6bf0aab709fb68c18e26f9fe7503b7  <=  0;
                end else begin
                    Ia44bcc8308360d3e6fa351bc108df3fa  <=  ~I1f36f045becec7f0528f4a935d3da2ff + 1;
                    Icf6bf0aab709fb68c18e26f9fe7503b7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2728682c0f749d1a9e8afeacdf44bfb7 == I27968f9d2e9dc75bfa55b1e5ad6f8c8e ) begin
                    Ib29a26c41a3ba089efd30c3256106a7c  <= I530fe7720e3bcda35e940aa4973a7da4;
                    I15947ee18296366e3e13cc9727ad2ebb  <=  0;
                end else begin
                    Ib29a26c41a3ba089efd30c3256106a7c  <=  ~I530fe7720e3bcda35e940aa4973a7da4 + 1;
                    I15947ee18296366e3e13cc9727ad2ebb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2728682c0f749d1a9e8afeacdf44bfb7 == Id53e488ea1a69e9d1e50dc276c14bb43 ) begin
                    I8999f385aaf15b67e4c12e56c7dba7cc  <= I03069dda9fa863172d8747408800eeba;
                    I23b16e4f6f2fab529ae42009d38cee85  <=  0;
                end else begin
                    I8999f385aaf15b67e4c12e56c7dba7cc  <=  ~I03069dda9fa863172d8747408800eeba + 1;
                    I23b16e4f6f2fab529ae42009d38cee85  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2728682c0f749d1a9e8afeacdf44bfb7 == I8440ba68619a5a3aad3510ad6ecaaea6 ) begin
                    I202980f6263e3b312c38061224992740  <= Ie7f36ee89f2b092555fbf8031d2347d9;
                    I51e128a639866ca032029880ae59e874  <=  0;
                end else begin
                    I202980f6263e3b312c38061224992740  <=  ~Ie7f36ee89f2b092555fbf8031d2347d9 + 1;
                    I51e128a639866ca032029880ae59e874  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I07da3bb5f943db6271fe1867a358df35 == I9e00e6e111b313b2efd5c9d32eae6a8e ) begin
                    I1fd9ed3763ff0ce0a671360f83bc3613  <= I18af7980562b28c537be3bea8dc5252b;
                    Ib14c75f869e8f09519517f3fcbdfaa7b  <=  0;
                end else begin
                    I1fd9ed3763ff0ce0a671360f83bc3613  <=  ~I18af7980562b28c537be3bea8dc5252b + 1;
                    Ib14c75f869e8f09519517f3fcbdfaa7b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I07da3bb5f943db6271fe1867a358df35 == I1836b01cfa5570153a8e4387baee29d6 ) begin
                    I4b58194aa6a5b5c825f14bb926a0ae9f  <= I22ec20f9396d28ed39c5fc4bf060c44a;
                    I9ceea65912b0a100eaa0afb42e84e5bd  <=  0;
                end else begin
                    I4b58194aa6a5b5c825f14bb926a0ae9f  <=  ~I22ec20f9396d28ed39c5fc4bf060c44a + 1;
                    I9ceea65912b0a100eaa0afb42e84e5bd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I07da3bb5f943db6271fe1867a358df35 == Icad06a6e006badf38d87cd3c4fd0981a ) begin
                    I706daad77f6a6eddf5576c238fa4714d  <= I105eac4e38f4661c7c7ca32161e42baa;
                    Id93be78cd06b38e1d7ec35ee66f878c3  <=  0;
                end else begin
                    I706daad77f6a6eddf5576c238fa4714d  <=  ~I105eac4e38f4661c7c7ca32161e42baa + 1;
                    Id93be78cd06b38e1d7ec35ee66f878c3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I07da3bb5f943db6271fe1867a358df35 == I8c061e6f5fb7e2be23d69254f0d0f59c ) begin
                    Ibceceead1cdcf8805e9a9f93b3b783ca  <= I5030734bfa54065cbef20c1350cd647d;
                    Ia61e18c0042f8ec7abb670e7f0648b45  <=  0;
                end else begin
                    Ibceceead1cdcf8805e9a9f93b3b783ca  <=  ~I5030734bfa54065cbef20c1350cd647d + 1;
                    Ia61e18c0042f8ec7abb670e7f0648b45  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I07da3bb5f943db6271fe1867a358df35 == I5411a76d49de45984ac852d98159ef5d ) begin
                    Ia5956c899daaaa0b2b0c16f524feaf98  <= Ieccf25e3abd6bae7dcf08baf815f3439;
                    I117b1ef192f2b24c6764c2d96864cc5f  <=  0;
                end else begin
                    Ia5956c899daaaa0b2b0c16f524feaf98  <=  ~Ieccf25e3abd6bae7dcf08baf815f3439 + 1;
                    I117b1ef192f2b24c6764c2d96864cc5f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61fc44808c85a75909b9d9fd4035f147 == I826369ad5207f64f64ff58abdb9f321e ) begin
                    I7f353333180ccbf6a271c9745430b199  <= I600c21fca7901299f8e95e8fa0ea0eb0;
                    If5224b5f45318dac2a64dcc72c6afad1  <=  0;
                end else begin
                    I7f353333180ccbf6a271c9745430b199  <=  ~I600c21fca7901299f8e95e8fa0ea0eb0 + 1;
                    If5224b5f45318dac2a64dcc72c6afad1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61fc44808c85a75909b9d9fd4035f147 == I4c266cd72fd1cd92f21511071a51c361 ) begin
                    I958f0106e3ffe429d0450f4b6e9ada3d  <= Ic4363dfd133124dd45ec2211499d0788;
                    I41710bb2545ba34f65e6d9a24086185b  <=  0;
                end else begin
                    I958f0106e3ffe429d0450f4b6e9ada3d  <=  ~Ic4363dfd133124dd45ec2211499d0788 + 1;
                    I41710bb2545ba34f65e6d9a24086185b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61fc44808c85a75909b9d9fd4035f147 == I76aac239cb31a0bdcebd7a3e3829f274 ) begin
                    Idf02454b4aacb6ff03288bb19a4771b1  <= I7c0bc779c09847e3beb0a139e8826511;
                    I15a9f9397a5d23e6885ac887723a8a19  <=  0;
                end else begin
                    Idf02454b4aacb6ff03288bb19a4771b1  <=  ~I7c0bc779c09847e3beb0a139e8826511 + 1;
                    I15a9f9397a5d23e6885ac887723a8a19  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61fc44808c85a75909b9d9fd4035f147 == Ief0092617ed13bebb791c57c0da0b12e ) begin
                    I42f39cecfe5c3d77b3fffb624cdb2c0b  <= If64db4386bf8f7d07292f14e3b313520;
                    I46f40fec14e2e6d5060c97f0a0d86696  <=  0;
                end else begin
                    I42f39cecfe5c3d77b3fffb624cdb2c0b  <=  ~If64db4386bf8f7d07292f14e3b313520 + 1;
                    I46f40fec14e2e6d5060c97f0a0d86696  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61fc44808c85a75909b9d9fd4035f147 == If1a6e0ead8f7aec9046bf22a1f59cf68 ) begin
                    Id7b0871cafd2630ba4dfc3e058613908  <= Ibf51e537b992c4b4c0539dda9948f45c;
                    I06e512c9097f76687d65c87f99c74764  <=  0;
                end else begin
                    Id7b0871cafd2630ba4dfc3e058613908  <=  ~Ibf51e537b992c4b4c0539dda9948f45c + 1;
                    I06e512c9097f76687d65c87f99c74764  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f == I26ee3d378528d4a8469eee34a7b5652e ) begin
                    I18c1c4d71799c5da8172f6cc63d2d37f  <= I9f83063bdc3c352024f702cb9dc71ce8;
                    I17759c97920685cd28c898441838531b  <=  0;
                end else begin
                    I18c1c4d71799c5da8172f6cc63d2d37f  <=  ~I9f83063bdc3c352024f702cb9dc71ce8 + 1;
                    I17759c97920685cd28c898441838531b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f == Ic8f3b5e177f927b64f1213625abc76c2 ) begin
                    I7d53f3ce487b0a2446d5205868c29175  <= I72127f6d422ec68dcd47126b87b3d3b1;
                    Ie7da1180f2c4eb8153421db4c6317a50  <=  0;
                end else begin
                    I7d53f3ce487b0a2446d5205868c29175  <=  ~I72127f6d422ec68dcd47126b87b3d3b1 + 1;
                    Ie7da1180f2c4eb8153421db4c6317a50  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f == Ia813a2600edc508e2eb59a9856e8fc4f ) begin
                    I37fb9120bfe27a0e7449583dda735479  <= I0b4a1b48d110b820d8d87f6e94d32988;
                    Ie6fe42c4fa7e64067960cab4edee83d5  <=  0;
                end else begin
                    I37fb9120bfe27a0e7449583dda735479  <=  ~I0b4a1b48d110b820d8d87f6e94d32988 + 1;
                    Ie6fe42c4fa7e64067960cab4edee83d5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f == Id04ad2fc64d6c346ae479abcbf3df41a ) begin
                    Ie7e15e6743a750cbf1b272da694b47dd  <= I2e3aeede695007fabe0d6247a93ed403;
                    Ic064e5425fd7a36be5860a40bc765994  <=  0;
                end else begin
                    Ie7e15e6743a750cbf1b272da694b47dd  <=  ~I2e3aeede695007fabe0d6247a93ed403 + 1;
                    Ic064e5425fd7a36be5860a40bc765994  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic5075ee0ad355c20dd45ed594f2a8c3f == I2827f1757a4ffc394869610f710291c4 ) begin
                    I66a1e62b25bce18e36d78c382b40b1df  <= I8c5ea3dc59fdcdea1c5f503dde1e815f;
                    Ifc8326ba561071589aec67a7de4276fb  <=  0;
                end else begin
                    I66a1e62b25bce18e36d78c382b40b1df  <=  ~I8c5ea3dc59fdcdea1c5f503dde1e815f + 1;
                    Ifc8326ba561071589aec67a7de4276fb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc == Ic8c6fbb1e7408869e5d11d0aea83203b ) begin
                    I9b81ec12daf51cb61f7dc0b9ad01cc1d  <= I873c4dbe95220e40d7388870520261bd;
                    Ibc55f69c8c895e9fad768b4b1a4a7a20  <=  0;
                end else begin
                    I9b81ec12daf51cb61f7dc0b9ad01cc1d  <=  ~I873c4dbe95220e40d7388870520261bd + 1;
                    Ibc55f69c8c895e9fad768b4b1a4a7a20  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc == Ibe0134da146c0c96af213013c5215943 ) begin
                    I9d76cb6c99a69086774f7fd471dadf53  <= I561fa67a9bfbedffcb04e7a4d6b76a64;
                    I50b89d077d160ee7d56376ae0abd9c6a  <=  0;
                end else begin
                    I9d76cb6c99a69086774f7fd471dadf53  <=  ~I561fa67a9bfbedffcb04e7a4d6b76a64 + 1;
                    I50b89d077d160ee7d56376ae0abd9c6a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc == I46a2e76ccab8ae201f78845054028074 ) begin
                    I4c59798356c8e05f8b2cdb4e202fc4bb  <= Ia55752d6c4f20378ff570a661ab31d9a;
                    I59a2c5b8dc1924b8503c24efa60c0c4a  <=  0;
                end else begin
                    I4c59798356c8e05f8b2cdb4e202fc4bb  <=  ~Ia55752d6c4f20378ff570a661ab31d9a + 1;
                    I59a2c5b8dc1924b8503c24efa60c0c4a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc == I1ee771cad3766a589cd62746062401c4 ) begin
                    I395b43b11730131a5f4331b2ce82717d  <= Ia13307be43e9155ed0333df62ccc8bf2;
                    I57a7c62f6cdf0fa0bd65df83a4904e36  <=  0;
                end else begin
                    I395b43b11730131a5f4331b2ce82717d  <=  ~Ia13307be43e9155ed0333df62ccc8bf2 + 1;
                    I57a7c62f6cdf0fa0bd65df83a4904e36  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic0a651f45a502ead495cf14f97d65bfc == Ic37d0375083a9415f7c0e9650ef0ecb7 ) begin
                    Ib3f07793c2e2cf7b6ac988be01a55829  <= I07b3d1451487a55fbbedda48b0cb6c73;
                    I733e71d48b2ae728b9d7b6a86261a156  <=  0;
                end else begin
                    Ib3f07793c2e2cf7b6ac988be01a55829  <=  ~I07b3d1451487a55fbbedda48b0cb6c73 + 1;
                    I733e71d48b2ae728b9d7b6a86261a156  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c == I73167dd9e24b49f6af3f7493cc2f9c0f ) begin
                    I05ad19dc723fe482f93cb524c8c86cf6  <= I9f8cf1a6cd0182fba35a49bd232f062a;
                    I20386e26c247b478dd7f2c89e73a1016  <=  0;
                end else begin
                    I05ad19dc723fe482f93cb524c8c86cf6  <=  ~I9f8cf1a6cd0182fba35a49bd232f062a + 1;
                    I20386e26c247b478dd7f2c89e73a1016  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c == I156970479a68c248bffd30be0097ff8f ) begin
                    I1db8d47c1852578aa6325919279419b1  <= Ie2e488a8589559deeec8598cf6726f1f;
                    Iaa6dcd47c9356b0b3b93d83f87c7fa05  <=  0;
                end else begin
                    I1db8d47c1852578aa6325919279419b1  <=  ~Ie2e488a8589559deeec8598cf6726f1f + 1;
                    Iaa6dcd47c9356b0b3b93d83f87c7fa05  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c == I851f4bdd95d1297f7ff05f01830c93fe ) begin
                    I98ec1bdbb599febfcdc06dbf807ab781  <= I9118ee5ff8c9ba9b125e5baa07bf52e0;
                    I8913043709d09e66411b5e70b0e3c969  <=  0;
                end else begin
                    I98ec1bdbb599febfcdc06dbf807ab781  <=  ~I9118ee5ff8c9ba9b125e5baa07bf52e0 + 1;
                    I8913043709d09e66411b5e70b0e3c969  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c == If6f8ef7f0cc4860dfb264b645ab0898f ) begin
                    I86f73b27c90bbd800b521fb8953d5506  <= I13b894057e2deae2c00787385de252a8;
                    Ifdcd9ff3c567f73e0366261dd09dee05  <=  0;
                end else begin
                    I86f73b27c90bbd800b521fb8953d5506  <=  ~I13b894057e2deae2c00787385de252a8 + 1;
                    Ifdcd9ff3c567f73e0366261dd09dee05  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic1c05ea22f708f620f626cc8c5ca309c == I5b983a4c1b35218893ed1bb0aaae26c8 ) begin
                    Id117870de7302febd51da982ab8b524e  <= I7797a3ea5b97b514a797243cf9fe890a;
                    I95af25eeba42e7fb3dc0dff9b702f61e  <=  0;
                end else begin
                    Id117870de7302febd51da982ab8b524e  <=  ~I7797a3ea5b97b514a797243cf9fe890a + 1;
                    I95af25eeba42e7fb3dc0dff9b702f61e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61a18378aadae4556da501ce997321b4 == Ifd281eb29091bcaf3a2929983366e637 ) begin
                    I6cff1d82f4c1bf7789e39b964dd9e6fe  <= I3af78697aacc410108d0be7fd13c686b;
                    Idf7fd041b837ee19551784f305c4efa1  <=  0;
                end else begin
                    I6cff1d82f4c1bf7789e39b964dd9e6fe  <=  ~I3af78697aacc410108d0be7fd13c686b + 1;
                    Idf7fd041b837ee19551784f305c4efa1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61a18378aadae4556da501ce997321b4 == I5ef5030a4e29e5e3c981d2616cae1ccd ) begin
                    I5d9786c9b4566669e7981654c3c10da7  <= I871cb63247618a543b444aa3f888fffe;
                    Ida9601d0e04fcfa1e448b681c4aa6bdc  <=  0;
                end else begin
                    I5d9786c9b4566669e7981654c3c10da7  <=  ~I871cb63247618a543b444aa3f888fffe + 1;
                    Ida9601d0e04fcfa1e448b681c4aa6bdc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61a18378aadae4556da501ce997321b4 == I3051150debf8f223b936ea5f169623f8 ) begin
                    I83dd9071e7e35d7165d556a67d2d1658  <= I124404013f8fc6b302661900b9ad8ed8;
                    Ibf6735fa3cd381ba501ab67979729a08  <=  0;
                end else begin
                    I83dd9071e7e35d7165d556a67d2d1658  <=  ~I124404013f8fc6b302661900b9ad8ed8 + 1;
                    Ibf6735fa3cd381ba501ab67979729a08  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61a18378aadae4556da501ce997321b4 == I9b76f1b49c0faf3f89256a1fe04c4597 ) begin
                    Id62c5db9d4a4e5eb91ca4b6876d36a9d  <= I8e413271c9d13748a1aa2d1a018ff28f;
                    Ic78e2d18e11538916e6726418f181e48  <=  0;
                end else begin
                    Id62c5db9d4a4e5eb91ca4b6876d36a9d  <=  ~I8e413271c9d13748a1aa2d1a018ff28f + 1;
                    Ic78e2d18e11538916e6726418f181e48  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61a18378aadae4556da501ce997321b4 == I62626dac5bf648ffad6e6e3cd836ab9c ) begin
                    Ibeb5414f37bbb8176c1a9ac51957dba0  <= I4d799e93b4dfcabd69977ddb25634a69;
                    I4b62c23b8d6b70c44af359b951424df1  <=  0;
                end else begin
                    Ibeb5414f37bbb8176c1a9ac51957dba0  <=  ~I4d799e93b4dfcabd69977ddb25634a69 + 1;
                    I4b62c23b8d6b70c44af359b951424df1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 == Ic527dbbf40cb847b5e5400f177a635da ) begin
                    If40561e9d6ab97e7dc2c6eca6d0725d8  <= I1487f0027b7d16f4bc85bb00e537cbaf;
                    If6467cc6d4b393b76586f5b65ace1435  <=  0;
                end else begin
                    If40561e9d6ab97e7dc2c6eca6d0725d8  <=  ~I1487f0027b7d16f4bc85bb00e537cbaf + 1;
                    If6467cc6d4b393b76586f5b65ace1435  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 == I44683db6537a0ae1bfdca8b6448c3772 ) begin
                    I630618151200231dda94b3fb59a24829  <= I1a5cdaa10022adf0ffbbc0f58b3e690a;
                    I1e79f24aac8988678a3ac91e9dfa493c  <=  0;
                end else begin
                    I630618151200231dda94b3fb59a24829  <=  ~I1a5cdaa10022adf0ffbbc0f58b3e690a + 1;
                    I1e79f24aac8988678a3ac91e9dfa493c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 == I5a03f223dea2bc87a454b29c3fe6058b ) begin
                    I45948c2ccae2bd2c2fcfe9c75787e2b4  <= I98246759d003e9bc6676ceb2d093a06b;
                    Ie3e87c23a6fbd77afb7a98ba764d937c  <=  0;
                end else begin
                    I45948c2ccae2bd2c2fcfe9c75787e2b4  <=  ~I98246759d003e9bc6676ceb2d093a06b + 1;
                    Ie3e87c23a6fbd77afb7a98ba764d937c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 == I8a7824d737ac024ffd25428f6599c070 ) begin
                    I73048e349b470dbb16b2b3e69aebcb3f  <= Ia3c2dfb3c4a45091be7cfecfad11f3ec;
                    I6406707a5545040df609c67f677e983d  <=  0;
                end else begin
                    I73048e349b470dbb16b2b3e69aebcb3f  <=  ~Ia3c2dfb3c4a45091be7cfecfad11f3ec + 1;
                    I6406707a5545040df609c67f677e983d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1fc521709a1ce2198fd8df5b41d0177 == Ia7e5724b4f05b0b6bdedaf264e797855 ) begin
                    Ic3a706eeb522f64147d4946983a9fcb4  <= I74cda651bcb24472a7697ba017f831a4;
                    I6aacacd072438b5172d5bd0be77c9ff8  <=  0;
                end else begin
                    Ic3a706eeb522f64147d4946983a9fcb4  <=  ~I74cda651bcb24472a7697ba017f831a4 + 1;
                    I6aacacd072438b5172d5bd0be77c9ff8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 == Ic8d1cb210627d8d6e717625ad3dd0fbe ) begin
                    Id8934e8818877e81d701105823366043  <= Id7ba55b14ac0f471142011dc2d57cc4b;
                    Ifea8a5d86f6681180539911cf637e785  <=  0;
                end else begin
                    Id8934e8818877e81d701105823366043  <=  ~Id7ba55b14ac0f471142011dc2d57cc4b + 1;
                    Ifea8a5d86f6681180539911cf637e785  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 == I313adb9858a6a31cce5af3d108459bb8 ) begin
                    Id5fd5653bfa014fa0e956ef4b1d83291  <= I5890643c88c4255a0e5efd45f8af3ee2;
                    I8101cabc2e8401f77a50d561a53b385f  <=  0;
                end else begin
                    Id5fd5653bfa014fa0e956ef4b1d83291  <=  ~I5890643c88c4255a0e5efd45f8af3ee2 + 1;
                    I8101cabc2e8401f77a50d561a53b385f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 == I36dd39ffe6e62b2518e12bb8e544ac20 ) begin
                    I41821f6b5a613fde6539e41a6a0c7b65  <= I4f53e4955e9e506a7169ae810da5dde6;
                    I9574b260963de729540209c0138de41c  <=  0;
                end else begin
                    I41821f6b5a613fde6539e41a6a0c7b65  <=  ~I4f53e4955e9e506a7169ae810da5dde6 + 1;
                    I9574b260963de729540209c0138de41c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 == I94337aa2c4ca0ec7a962962780f21f11 ) begin
                    Ie8d437ed136f7f5971638d1f62ffdf15  <= Ifc7c1ea337b122fb720767f1890f1a6a;
                    I791728546a36e98c0d5c4eb1063082b3  <=  0;
                end else begin
                    Ie8d437ed136f7f5971638d1f62ffdf15  <=  ~Ifc7c1ea337b122fb720767f1890f1a6a + 1;
                    I791728546a36e98c0d5c4eb1063082b3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1bb5511c9cda1a595c45ecde48e9ebc7 == Ib2443922534953e49e1af5343c028fc6 ) begin
                    Iaf46eedc430b55905d73486ac0752c8f  <= Id40d6f3a8dd09678b25b3e579dd5fb68;
                    I338183bc2bdb39e2a3820a768d78ebdc  <=  0;
                end else begin
                    Iaf46eedc430b55905d73486ac0752c8f  <=  ~Id40d6f3a8dd09678b25b3e579dd5fb68 + 1;
                    I338183bc2bdb39e2a3820a768d78ebdc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4a29c37ed36b6e12f1f8e263c92bdbc1 == I08d6c121fbd306f3908a88ce10779ac5 ) begin
                    I32671ef3896bd0b586f13c092dd04b9e  <= I7002830b0a5f40ba2a2fe7a00c7b6d58;
                    I4197bb0d6d0465aeb6fd7f0a8189a368  <=  0;
                end else begin
                    I32671ef3896bd0b586f13c092dd04b9e  <=  ~I7002830b0a5f40ba2a2fe7a00c7b6d58 + 1;
                    I4197bb0d6d0465aeb6fd7f0a8189a368  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4a29c37ed36b6e12f1f8e263c92bdbc1 == I1b947b03d2db27afe8faf78f580c90aa ) begin
                    Ie8bfdf207d647c9f161bdf265a8472b4  <= I3f377e8994959ef8182a08538e393d9a;
                    I8f0d7e1f97b611f6c4a231338aaba68e  <=  0;
                end else begin
                    Ie8bfdf207d647c9f161bdf265a8472b4  <=  ~I3f377e8994959ef8182a08538e393d9a + 1;
                    I8f0d7e1f97b611f6c4a231338aaba68e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4a29c37ed36b6e12f1f8e263c92bdbc1 == I05b4915602c4c635f9e91ff69432ebf2 ) begin
                    Id44fe933294cafff88d133a0ddc1a832  <= I71bf29f3519e3238cec112ef97ce0579;
                    Ie50a86c3b69d3884c72948133083e099  <=  0;
                end else begin
                    Id44fe933294cafff88d133a0ddc1a832  <=  ~I71bf29f3519e3238cec112ef97ce0579 + 1;
                    Ie50a86c3b69d3884c72948133083e099  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4a29c37ed36b6e12f1f8e263c92bdbc1 == Ifdd87b92e70f345ca64fa4e96d732210 ) begin
                    I20c1f8e56a14db0665160ecbb277fb1a  <= Iaa4bc2f51984f383479b597e6cd4c873;
                    I2cf91b227a82701d912cf9e9e1040ddc  <=  0;
                end else begin
                    I20c1f8e56a14db0665160ecbb277fb1a  <=  ~Iaa4bc2f51984f383479b597e6cd4c873 + 1;
                    I2cf91b227a82701d912cf9e9e1040ddc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4bf02a07719402890405fb2e7b679ed9 == I67335037a5b54e1b5bb316cd3519e790 ) begin
                    I7627f96e870f6a3e8abd7ac494bc178c  <= I9066a5cf776f80ebf89bdac1f2edb4ac;
                    I0f50e2edf3586292da17ce7214d37038  <=  0;
                end else begin
                    I7627f96e870f6a3e8abd7ac494bc178c  <=  ~I9066a5cf776f80ebf89bdac1f2edb4ac + 1;
                    I0f50e2edf3586292da17ce7214d37038  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4bf02a07719402890405fb2e7b679ed9 == Ic0feb7035ff8f8962a79aa20f4129bbe ) begin
                    Ia2d3997dce108f85ed64e88780e99efa  <= I7319203d7231bebb6d6e52422cce5ed2;
                    Id7666dd5135e45a1e42f13ffbb8558ed  <=  0;
                end else begin
                    Ia2d3997dce108f85ed64e88780e99efa  <=  ~I7319203d7231bebb6d6e52422cce5ed2 + 1;
                    Id7666dd5135e45a1e42f13ffbb8558ed  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4bf02a07719402890405fb2e7b679ed9 == If11c3d720e491cfc18684f3a23f6b93b ) begin
                    I6a25dc88186816258f1237123ee4968f  <= I4e8309976fd6011d78728cef935dc3c1;
                    I3dbcf0199e35f410c38ab3d9e2cac2ef  <=  0;
                end else begin
                    I6a25dc88186816258f1237123ee4968f  <=  ~I4e8309976fd6011d78728cef935dc3c1 + 1;
                    I3dbcf0199e35f410c38ab3d9e2cac2ef  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4bf02a07719402890405fb2e7b679ed9 == I5d4a36427e26532bca590796e4107dcc ) begin
                    Ia9d61848b5384a8cc63321201174f3d3  <= I5ed502118c175d5bdb4607973554a3a3;
                    I06c6db30fc7e63facd144d0166702e6a  <=  0;
                end else begin
                    Ia9d61848b5384a8cc63321201174f3d3  <=  ~I5ed502118c175d5bdb4607973554a3a3 + 1;
                    I06c6db30fc7e63facd144d0166702e6a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I75bd82990cb60b6d7ccd7aa2982da7aa == Ib0eb8c6ddbbcd4825e8fc5b1c55495b3 ) begin
                    I53ed79856aae53b180f28b47822e89b6  <= If457f80b3d29b60b840f886fa928297c;
                    Id20d5070afe5748b50833f0593777c49  <=  0;
                end else begin
                    I53ed79856aae53b180f28b47822e89b6  <=  ~If457f80b3d29b60b840f886fa928297c + 1;
                    Id20d5070afe5748b50833f0593777c49  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I75bd82990cb60b6d7ccd7aa2982da7aa == I0d5ab203120026f15a1d563bb65fa1ab ) begin
                    I76503bcb779e039edc9acfc03a2d1ee6  <= I7e0f785ec7554540c9a4a413a3afa75f;
                    I3d041f7cf6c679d8d9677445eac96640  <=  0;
                end else begin
                    I76503bcb779e039edc9acfc03a2d1ee6  <=  ~I7e0f785ec7554540c9a4a413a3afa75f + 1;
                    I3d041f7cf6c679d8d9677445eac96640  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I75bd82990cb60b6d7ccd7aa2982da7aa == I35ca485dc9ef601029877a4ee46ed942 ) begin
                    I18ae85d6725cf0ab3b69bedeef651425  <= Id3662bbe1b5191995d1656045fe6b6a6;
                    I51d27603f0a87b78857b8e064182d925  <=  0;
                end else begin
                    I18ae85d6725cf0ab3b69bedeef651425  <=  ~Id3662bbe1b5191995d1656045fe6b6a6 + 1;
                    I51d27603f0a87b78857b8e064182d925  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I75bd82990cb60b6d7ccd7aa2982da7aa == I8c1c4b4851ed06bce6af5b392c75c6b8 ) begin
                    Iaa3bbfc6704e70a55b8e1083c326820f  <= Idf922fab93bc2357ac1f66f73f3ead0b;
                    I9b6d48e71d050b9b0b5c5e7407288103  <=  0;
                end else begin
                    Iaa3bbfc6704e70a55b8e1083c326820f  <=  ~Idf922fab93bc2357ac1f66f73f3ead0b + 1;
                    I9b6d48e71d050b9b0b5c5e7407288103  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia6d3e38249f8a1208540b68f54c46769 == I00fc4e266ce9e790501c78809bfae38e ) begin
                    I8c1c3ee4b57d56ab362672dfeb4e0ae9  <= I780371393ef898aa144c5bc36e74c654;
                    Id05706fe9e0fc4776e0446aacd4c118d  <=  0;
                end else begin
                    I8c1c3ee4b57d56ab362672dfeb4e0ae9  <=  ~I780371393ef898aa144c5bc36e74c654 + 1;
                    Id05706fe9e0fc4776e0446aacd4c118d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia6d3e38249f8a1208540b68f54c46769 == I35fa53ff8ca5fab19b6de45beda84ff2 ) begin
                    Ic8e0765b1cf95f2578a7ec656d027f6e  <= I79696cd10cffa4c0181a2089da6b3262;
                    I2ec61e0e1b707857ca39f532bf970e03  <=  0;
                end else begin
                    Ic8e0765b1cf95f2578a7ec656d027f6e  <=  ~I79696cd10cffa4c0181a2089da6b3262 + 1;
                    I2ec61e0e1b707857ca39f532bf970e03  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia6d3e38249f8a1208540b68f54c46769 == If3c4067202f592fabf77cd76db5575dd ) begin
                    I39eaefaae486119c8741c5e9b7f85bd3  <= I073155ab0359a13b77f730653dcfc08d;
                    Ibd1b4a1010823cc9e4a78a0fcefd7d01  <=  0;
                end else begin
                    I39eaefaae486119c8741c5e9b7f85bd3  <=  ~I073155ab0359a13b77f730653dcfc08d + 1;
                    Ibd1b4a1010823cc9e4a78a0fcefd7d01  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia6d3e38249f8a1208540b68f54c46769 == I64276a920c9ccf7576c15618812fd152 ) begin
                    I6ac8d8000e434fcca222525ac00f9849  <= I1b44f781d81438654f69bb7fbdb94011;
                    I6da2861072f65e35d46d224b982eda7a  <=  0;
                end else begin
                    I6ac8d8000e434fcca222525ac00f9849  <=  ~I1b44f781d81438654f69bb7fbdb94011 + 1;
                    I6da2861072f65e35d46d224b982eda7a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idf548b72357ab28fd956791e84e5d65c == I478a999d16ad8a5266769d1b8caa79db ) begin
                    I114cfd3fe8f5db92b879e0dce592af3b  <= Id68f1a0ec8ff80da3190fe517bd935e3;
                    I860c7e185d38d907c4ed20a64d238dd6  <=  0;
                end else begin
                    I114cfd3fe8f5db92b879e0dce592af3b  <=  ~Id68f1a0ec8ff80da3190fe517bd935e3 + 1;
                    I860c7e185d38d907c4ed20a64d238dd6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idf548b72357ab28fd956791e84e5d65c == I29f2854aec43820204ceb8f3eceed6c9 ) begin
                    I8db1c7f6b5c7c04f71e7fcc18f7b9941  <= I3704464d41956032b779eebe27511815;
                    I76e06fe466c43e4aef0ef860f0274fa8  <=  0;
                end else begin
                    I8db1c7f6b5c7c04f71e7fcc18f7b9941  <=  ~I3704464d41956032b779eebe27511815 + 1;
                    I76e06fe466c43e4aef0ef860f0274fa8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idf548b72357ab28fd956791e84e5d65c == Idf664119a34b4692c0cfaa4c742480f4 ) begin
                    I89e516738a408ccbd495e4f5aeeb38a6  <= Ie6756ee9631791940ffc6fddb223b4d0;
                    I3c00d8a5dd8c99ee527ad4180e469ab7  <=  0;
                end else begin
                    I89e516738a408ccbd495e4f5aeeb38a6  <=  ~Ie6756ee9631791940ffc6fddb223b4d0 + 1;
                    I3c00d8a5dd8c99ee527ad4180e469ab7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idf548b72357ab28fd956791e84e5d65c == Iae32c64d9bf268ccacaec2d40efe70f4 ) begin
                    I0c02b9318bc4f50969f8d486e587a627  <= I085151dfc2e773a7a485f5ef1b7cd6bd;
                    Iba2018bad14888e510fc7f4a4e040ed5  <=  0;
                end else begin
                    I0c02b9318bc4f50969f8d486e587a627  <=  ~I085151dfc2e773a7a485f5ef1b7cd6bd + 1;
                    Iba2018bad14888e510fc7f4a4e040ed5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I50b6f2e0ef2831535ac8c18cd7ca9379 == If30e09a7c080fd91758eacb33912b8d6 ) begin
                    I79224b17e2d1f87175f3118287351e0e  <= I2654e83fff153df7760c341f59a23396;
                    I2e3d469ef08219887c92189ad3759da9  <=  0;
                end else begin
                    I79224b17e2d1f87175f3118287351e0e  <=  ~I2654e83fff153df7760c341f59a23396 + 1;
                    I2e3d469ef08219887c92189ad3759da9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I50b6f2e0ef2831535ac8c18cd7ca9379 == If000ebe4f2ddbec4afb6c0e41abb2f9c ) begin
                    I41ee2f859df1db26618ab9c2c0a57be5  <= Iee3eec7a9d7a3a5c22281545ec143e50;
                    I74628364cf049f0e6de34bd1f9853985  <=  0;
                end else begin
                    I41ee2f859df1db26618ab9c2c0a57be5  <=  ~Iee3eec7a9d7a3a5c22281545ec143e50 + 1;
                    I74628364cf049f0e6de34bd1f9853985  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I50b6f2e0ef2831535ac8c18cd7ca9379 == I714abef2427918d8967e5fff40fd48d7 ) begin
                    I15a667ea371ed0fd464f42fb9ef61766  <= Ied2b9ca07a6d498abada30fb0726df24;
                    Ifec818042c24c8eb96832c782f09ab04  <=  0;
                end else begin
                    I15a667ea371ed0fd464f42fb9ef61766  <=  ~Ied2b9ca07a6d498abada30fb0726df24 + 1;
                    Ifec818042c24c8eb96832c782f09ab04  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I50b6f2e0ef2831535ac8c18cd7ca9379 == I6229267ae259aa8193a90596f8c1d432 ) begin
                    I25c2d3dd7fedd28f0be0e3d8dccddff8  <= If95315702519e7a08386a870e599aab0;
                    I0aa52a892c8969087bf3f158aae7078a  <=  0;
                end else begin
                    I25c2d3dd7fedd28f0be0e3d8dccddff8  <=  ~If95315702519e7a08386a870e599aab0 + 1;
                    I0aa52a892c8969087bf3f158aae7078a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4003a2515229ca8eb6fefa2bef289ca6 == Iaa26fea88e8b3f2ce1d402b48c7a9eff ) begin
                    If22b31d70158d864ca6b0201ffc2b7c3  <= I1091064aef7d915ba8fb6cbded069102;
                    I31b799a3279d7d66b53f4be544498602  <=  0;
                end else begin
                    If22b31d70158d864ca6b0201ffc2b7c3  <=  ~I1091064aef7d915ba8fb6cbded069102 + 1;
                    I31b799a3279d7d66b53f4be544498602  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4003a2515229ca8eb6fefa2bef289ca6 == Idc0f6e44fa41f76f3ddff9628d25c005 ) begin
                    I7950b8505327240095538f60d81834d1  <= I40685c7d2c8be12698f734ec6213b5b4;
                    Ie8e004bf6e301a4ed9d9dcca91b2dc85  <=  0;
                end else begin
                    I7950b8505327240095538f60d81834d1  <=  ~I40685c7d2c8be12698f734ec6213b5b4 + 1;
                    Ie8e004bf6e301a4ed9d9dcca91b2dc85  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4003a2515229ca8eb6fefa2bef289ca6 == I7c14c6e871660c6c830de981c07f6b2d ) begin
                    Ib75297152c09323c7a6f674c93edc01f  <= Icc7775fe34c162006b93662530fd4944;
                    I9995a84609ef3fe477c73f136515ffe9  <=  0;
                end else begin
                    Ib75297152c09323c7a6f674c93edc01f  <=  ~Icc7775fe34c162006b93662530fd4944 + 1;
                    I9995a84609ef3fe477c73f136515ffe9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I4003a2515229ca8eb6fefa2bef289ca6 == Idc5ee83aa6a50531e6de2d9abaa26843 ) begin
                    Ie813deeac800a6b251209a1c8e2adb12  <= I2e6f1a5695ad23b8ca282b344832ee8e;
                    I54e519ab156fdf2054472d4684de064a  <=  0;
                end else begin
                    Ie813deeac800a6b251209a1c8e2adb12  <=  ~I2e6f1a5695ad23b8ca282b344832ee8e + 1;
                    I54e519ab156fdf2054472d4684de064a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I48672f8b83eef8c406694676746469e7 == Ie0ff06499371f17cb8c56c9f0c7ee666 ) begin
                    Iada283b3152a5316b6c7077292ac0a29  <= I016ce894bebdaa7e56af9deb1ccfb3f5;
                    I527950bde49a5c46e818225e41bec4f9  <=  0;
                end else begin
                    Iada283b3152a5316b6c7077292ac0a29  <=  ~I016ce894bebdaa7e56af9deb1ccfb3f5 + 1;
                    I527950bde49a5c46e818225e41bec4f9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I48672f8b83eef8c406694676746469e7 == I59976ed14d4be22603d2d164399389f9 ) begin
                    Ic14e12a907c5d6b7ad2615905a64886d  <= Iad2dd0815c1107160992e5070632f76c;
                    Ieb876e18857117935ca3aecb6a525b1f  <=  0;
                end else begin
                    Ic14e12a907c5d6b7ad2615905a64886d  <=  ~Iad2dd0815c1107160992e5070632f76c + 1;
                    Ieb876e18857117935ca3aecb6a525b1f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I48672f8b83eef8c406694676746469e7 == I9e94cdbd4a445883fb45fb3ed1b05d7b ) begin
                    Ife78b0889c9c7129a3000cca66ae4aa2  <= Iefaba2acd282081b9a0a98ed057ca85e;
                    If22f8fa601e72589b3a5779f23ca7454  <=  0;
                end else begin
                    Ife78b0889c9c7129a3000cca66ae4aa2  <=  ~Iefaba2acd282081b9a0a98ed057ca85e + 1;
                    If22f8fa601e72589b3a5779f23ca7454  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I48672f8b83eef8c406694676746469e7 == I581b4fe258cb92d51ffc1482da718625 ) begin
                    Id926d49513e089a52b17978a9ab84372  <= Id4ef94eb8d5db8810bca4c9d669f0b7f;
                    If222f8f81e40570854a512fe828f9ea9  <=  0;
                end else begin
                    Id926d49513e089a52b17978a9ab84372  <=  ~Id4ef94eb8d5db8810bca4c9d669f0b7f + 1;
                    If222f8f81e40570854a512fe828f9ea9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia14a60c9497c0faf3f1f448ff2abe553 == I19f794db275b2266dd9a91b3b0174329 ) begin
                    I4dfbf2a2c01ce39fea9b756f9b106fc2  <= I04e845e6a5ed71978b636593dd749b12;
                    I6bea78584853c37d7c4993a45668542a  <=  0;
                end else begin
                    I4dfbf2a2c01ce39fea9b756f9b106fc2  <=  ~I04e845e6a5ed71978b636593dd749b12 + 1;
                    I6bea78584853c37d7c4993a45668542a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia14a60c9497c0faf3f1f448ff2abe553 == I7d4b8ac371172cf90b31890df5693875 ) begin
                    Iad7cce628396ce9ffac3ba9dde7ac494  <= I0b2760b437be2cb79382f8d6a7b8969e;
                    Id7cd91008312189123519e44cfb2e141  <=  0;
                end else begin
                    Iad7cce628396ce9ffac3ba9dde7ac494  <=  ~I0b2760b437be2cb79382f8d6a7b8969e + 1;
                    Id7cd91008312189123519e44cfb2e141  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia14a60c9497c0faf3f1f448ff2abe553 == I1f02219120214ac3e5f5279031facc56 ) begin
                    Ib71f9f92515c200bd16591c656d69ee7  <= I1b0fdaeebe5fee6fbb2e13aac5e233a1;
                    Id3c95ac844fe01a85e6251683bb3f9cb  <=  0;
                end else begin
                    Ib71f9f92515c200bd16591c656d69ee7  <=  ~I1b0fdaeebe5fee6fbb2e13aac5e233a1 + 1;
                    Id3c95ac844fe01a85e6251683bb3f9cb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia14a60c9497c0faf3f1f448ff2abe553 == I569a8645fa9f5476d122bccc7f40fd75 ) begin
                    I8e39b301e04135b8ab88d54e7c1e22f7  <= Iee872d17e4a28075be0ad7086c3acc91;
                    I49b96dfb05812ec7b0632bc722d417df  <=  0;
                end else begin
                    I8e39b301e04135b8ab88d54e7c1e22f7  <=  ~Iee872d17e4a28075be0ad7086c3acc91 + 1;
                    I49b96dfb05812ec7b0632bc722d417df  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0ef3962dd323e8ec64c4a881bd4b3044 == Ie620ab2c461442bf7c7ddd962dd65839 ) begin
                    Idadba73fb37b81563818e82af3d89a58  <= I87656ddd4ef8f1ae36c7566d5e7892d8;
                    I89b8ac7adba1c7fe4f04e408857c92bc  <=  0;
                end else begin
                    Idadba73fb37b81563818e82af3d89a58  <=  ~I87656ddd4ef8f1ae36c7566d5e7892d8 + 1;
                    I89b8ac7adba1c7fe4f04e408857c92bc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0ef3962dd323e8ec64c4a881bd4b3044 == I3dc4a3e2c52f2f74aaf1e640543fcecb ) begin
                    Ic19accaf42ef2b61fb52ab3621622ef2  <= I865cd0535644db7f17db1180c85f1744;
                    Ic1a67160ca63763ce6b850bed5371d32  <=  0;
                end else begin
                    Ic19accaf42ef2b61fb52ab3621622ef2  <=  ~I865cd0535644db7f17db1180c85f1744 + 1;
                    Ic1a67160ca63763ce6b850bed5371d32  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0ef3962dd323e8ec64c4a881bd4b3044 == I749c798e403cefc3782b3a63de02e227 ) begin
                    I94f508ac67f07b73b3ff1d5aa5955eea  <= I71d46741fa94df65e1bdf6abff53d2ba;
                    Iaa1ed0cec8df6dec4fb0ef9c57c98d19  <=  0;
                end else begin
                    I94f508ac67f07b73b3ff1d5aa5955eea  <=  ~I71d46741fa94df65e1bdf6abff53d2ba + 1;
                    Iaa1ed0cec8df6dec4fb0ef9c57c98d19  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0ef3962dd323e8ec64c4a881bd4b3044 == I3ce1a50aa7de5d1dae422eed03c450b2 ) begin
                    Ieb8588293562c9c25897044b9e5ed6a4  <= Ic223d7941250d739ce9bb0ae5013646e;
                    I76465e13c5a9ac236635e663e543487c  <=  0;
                end else begin
                    Ieb8588293562c9c25897044b9e5ed6a4  <=  ~Ic223d7941250d739ce9bb0ae5013646e + 1;
                    I76465e13c5a9ac236635e663e543487c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9b64c34e31dab63c03b3de4528d53fe == Id9474b1f0f1ab396654b7048eea873c2 ) begin
                    I671d71d9ca760cc759b96bbacd361f90  <= I1ef9b548b943a1f2012b91c7e0b445f2;
                    Iff18998e317563a12db412950315b397  <=  0;
                end else begin
                    I671d71d9ca760cc759b96bbacd361f90  <=  ~I1ef9b548b943a1f2012b91c7e0b445f2 + 1;
                    Iff18998e317563a12db412950315b397  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9b64c34e31dab63c03b3de4528d53fe == Ib7d69d239aac1a9de86e2f2f1337c5f6 ) begin
                    I3f793de7fcfd045af3970e4ec219128b  <= I88b6d7894d82ff394e89c7471c80dd5b;
                    I279642da9295f410b7482eaedfbcde75  <=  0;
                end else begin
                    I3f793de7fcfd045af3970e4ec219128b  <=  ~I88b6d7894d82ff394e89c7471c80dd5b + 1;
                    I279642da9295f410b7482eaedfbcde75  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9b64c34e31dab63c03b3de4528d53fe == I40a799391b45437a24bf9c7cbc2ec409 ) begin
                    Id49f950b3679093b10f8b64ae89c5558  <= Ia5fc7e1f991f30042b848888a546534b;
                    Iecceba6850d58cd1500bb5129abc8035  <=  0;
                end else begin
                    Id49f950b3679093b10f8b64ae89c5558  <=  ~Ia5fc7e1f991f30042b848888a546534b + 1;
                    Iecceba6850d58cd1500bb5129abc8035  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie9b64c34e31dab63c03b3de4528d53fe == Id81eae2229fec7726aa687d711d1b998 ) begin
                    Ib70c7567e552969a2757c1f48a2468ef  <= If699df4c8261ebce5c5d1aebe062cd61;
                    I6ede97dfb1484ba6fe621c7034e22c0b  <=  0;
                end else begin
                    Ib70c7567e552969a2757c1f48a2468ef  <=  ~If699df4c8261ebce5c5d1aebe062cd61 + 1;
                    I6ede97dfb1484ba6fe621c7034e22c0b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5941476ded9f6dc25d7394f5d133955b == I7bab2b945804593835eb8b63143a3345 ) begin
                    I6dbd0c3ac9f2b3887d87e316b8b40b55  <= I19338369553e96bb2476d80fe84dec3e;
                    I57bf6d033eb5643e96bcdefcfeb76a46  <=  0;
                end else begin
                    I6dbd0c3ac9f2b3887d87e316b8b40b55  <=  ~I19338369553e96bb2476d80fe84dec3e + 1;
                    I57bf6d033eb5643e96bcdefcfeb76a46  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5941476ded9f6dc25d7394f5d133955b == I4e7f07fa261e44488cb5b0903d2e8c5d ) begin
                    I8c309d7fe6aaa8c996e39b8f3dfafef6  <= I9844ff02042cbc04dd5f4179908bbb2d;
                    I5ba33277f07eadbc27835afa96bdc535  <=  0;
                end else begin
                    I8c309d7fe6aaa8c996e39b8f3dfafef6  <=  ~I9844ff02042cbc04dd5f4179908bbb2d + 1;
                    I5ba33277f07eadbc27835afa96bdc535  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5941476ded9f6dc25d7394f5d133955b == I5d69471b78cf5aba461a12cfe6d7d11e ) begin
                    Iefdfd7b1924f8b6049b02576f9948027  <= I89cc6a060b714985b24f724adc782e7b;
                    I256096a960771679c9a7a391448aa711  <=  0;
                end else begin
                    Iefdfd7b1924f8b6049b02576f9948027  <=  ~I89cc6a060b714985b24f724adc782e7b + 1;
                    I256096a960771679c9a7a391448aa711  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5941476ded9f6dc25d7394f5d133955b == Iba0af171e17c12093f5dbde019fff4da ) begin
                    I2c14ee79492962576e12ff1698ac0fe1  <= I39d94ce7fbe37a74404e0043060441ed;
                    I220f38bf301ec4abcd1e07727fc5bae8  <=  0;
                end else begin
                    I2c14ee79492962576e12ff1698ac0fe1  <=  ~I39d94ce7fbe37a74404e0043060441ed + 1;
                    I220f38bf301ec4abcd1e07727fc5bae8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib46c78ff661ee6fb69c704d39235ffe1 == I580c7b678e4f2c08a4d521c335392c07 ) begin
                    I56e90395afb09c7d775111d19856da1d  <= I0a1c9a8d59dbcffd6847f3a65107c407;
                    Id6cabb7608d470ad7dec1951618efa8c  <=  0;
                end else begin
                    I56e90395afb09c7d775111d19856da1d  <=  ~I0a1c9a8d59dbcffd6847f3a65107c407 + 1;
                    Id6cabb7608d470ad7dec1951618efa8c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib46c78ff661ee6fb69c704d39235ffe1 == I8016fc36bc9614afef570a084942081e ) begin
                    I90f0c524f6b98c28d18db952ac40c83e  <= I2328556c467a9e639f2b6ba1d0cb99b7;
                    I30ac677d67ab06a6f5759da2717ef6e2  <=  0;
                end else begin
                    I90f0c524f6b98c28d18db952ac40c83e  <=  ~I2328556c467a9e639f2b6ba1d0cb99b7 + 1;
                    I30ac677d67ab06a6f5759da2717ef6e2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib46c78ff661ee6fb69c704d39235ffe1 == I744066a189658aad33b32468934ca485 ) begin
                    Id50649fc4e9de24fdd9f06499a733b87  <= I5c9d75d6431d69db1abe412e591000a7;
                    If0881734b6b8bb6e3e22823408203887  <=  0;
                end else begin
                    Id50649fc4e9de24fdd9f06499a733b87  <=  ~I5c9d75d6431d69db1abe412e591000a7 + 1;
                    If0881734b6b8bb6e3e22823408203887  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib46c78ff661ee6fb69c704d39235ffe1 == Ic2a5d82d3e19ff84f46d2d71b3d544eb ) begin
                    Ifc988e99b4c4c1ba2d5cf3a76695900d  <= I8dc3dcdefc85b6ff8ecfa09cfc7e69fa;
                    I29502a6df7b40a59cb84f6c1a0d30fbe  <=  0;
                end else begin
                    Ifc988e99b4c4c1ba2d5cf3a76695900d  <=  ~I8dc3dcdefc85b6ff8ecfa09cfc7e69fa + 1;
                    I29502a6df7b40a59cb84f6c1a0d30fbe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iadabc5abc7dfbc1dd747179ad7e37850 == I935a700d902a104974a961beca5ac99a ) begin
                    I53c579c64f0d911fe3fbc43dc3e981de  <= I69f6c909ea6b207c200b154e00e13a05;
                    Ied5d76051c9302e2594e5f1c34dbe8a9  <=  0;
                end else begin
                    I53c579c64f0d911fe3fbc43dc3e981de  <=  ~I69f6c909ea6b207c200b154e00e13a05 + 1;
                    Ied5d76051c9302e2594e5f1c34dbe8a9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iadabc5abc7dfbc1dd747179ad7e37850 == I902f91dfb3bada8a106f46923239c93a ) begin
                    Id729d27d6424495fdb4deb2ffc038f01  <= Id365c9f8f7f97c777bd5da0ce9490511;
                    If6c801f61074108c3342f1c3d0b4a39d  <=  0;
                end else begin
                    Id729d27d6424495fdb4deb2ffc038f01  <=  ~Id365c9f8f7f97c777bd5da0ce9490511 + 1;
                    If6c801f61074108c3342f1c3d0b4a39d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iadabc5abc7dfbc1dd747179ad7e37850 == I4d4f46a02cffbf72298704e8a0504fe2 ) begin
                    I8816c4edb8c7f5fd6e7a3c81013116ce  <= Idf0206d2ad2bdef7db1d30a2d715cc6a;
                    I3f15fe479ccd6715b63db728ffa8b49f  <=  0;
                end else begin
                    I8816c4edb8c7f5fd6e7a3c81013116ce  <=  ~Idf0206d2ad2bdef7db1d30a2d715cc6a + 1;
                    I3f15fe479ccd6715b63db728ffa8b49f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iadabc5abc7dfbc1dd747179ad7e37850 == Ie8fd35237928694738b464d52847c2b6 ) begin
                    I88ba486c5bca54f6c120a654b81e0a90  <= I07d1c54431eed887554a136f15f86d22;
                    Id7e322ddf8565bb59e6377bfc7b3ab36  <=  0;
                end else begin
                    I88ba486c5bca54f6c120a654b81e0a90  <=  ~I07d1c54431eed887554a136f15f86d22 + 1;
                    Id7e322ddf8565bb59e6377bfc7b3ab36  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I97a6b5f0976feceee3a5b5890d4d76a0 == Ib73fc8722db87e7be4b14ce361b79719 ) begin
                    Ie1ba6d92c19ebbc5c994d9da3881f6c9  <= Ic16809a3c82787ed88819fc9e9613f85;
                    I5a325c188a650a75ab298719c0287618  <=  0;
                end else begin
                    Ie1ba6d92c19ebbc5c994d9da3881f6c9  <=  ~Ic16809a3c82787ed88819fc9e9613f85 + 1;
                    I5a325c188a650a75ab298719c0287618  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I97a6b5f0976feceee3a5b5890d4d76a0 == Ifde9664e13fe94aca97da5824ef0c08e ) begin
                    I023278cb7d70d4608259e10c89e97117  <= I1613ae89442495e703a52e65b8a0bf9f;
                    I763f7f930d12bef17e0aa5ed0d6abf96  <=  0;
                end else begin
                    I023278cb7d70d4608259e10c89e97117  <=  ~I1613ae89442495e703a52e65b8a0bf9f + 1;
                    I763f7f930d12bef17e0aa5ed0d6abf96  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I97a6b5f0976feceee3a5b5890d4d76a0 == I3d25580e525216c23557ffa5ed998bab ) begin
                    Ib8c744194310bd59e983e392b828e9b4  <= I6089da825af433e847c0b1bb9ff7d373;
                    I0e34522d1f95f50998246232512bb60c  <=  0;
                end else begin
                    Ib8c744194310bd59e983e392b828e9b4  <=  ~I6089da825af433e847c0b1bb9ff7d373 + 1;
                    I0e34522d1f95f50998246232512bb60c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I97a6b5f0976feceee3a5b5890d4d76a0 == Ia3d21a8d9a8c24b112965d6eb966de8c ) begin
                    Iaa2aba39e0454008fbeff8f9aa87a481  <= I6aa7fccf4e225fa70063fd24dab74e6b;
                    I45b69f889fd15cce35f6812afe0f4894  <=  0;
                end else begin
                    Iaa2aba39e0454008fbeff8f9aa87a481  <=  ~I6aa7fccf4e225fa70063fd24dab74e6b + 1;
                    I45b69f889fd15cce35f6812afe0f4894  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7217d4790fec9797a1eb8cab1ebce71b == I7d7923beddaf4b873ae819914599f02f ) begin
                    I61a43aad15d7a9943f74617f434af306  <= Ibe2a5f680405f233256b6fd806b72ae5;
                    If4db281fdcf771156956dfa30e36b29c  <=  0;
                end else begin
                    I61a43aad15d7a9943f74617f434af306  <=  ~Ibe2a5f680405f233256b6fd806b72ae5 + 1;
                    If4db281fdcf771156956dfa30e36b29c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7217d4790fec9797a1eb8cab1ebce71b == Idc6a066b872fa91ce73e9aa21d668e83 ) begin
                    Ibd8114af3027bd3364395e7b94484272  <= I662d408ffd8fb9f249e531a167161429;
                    Ib312a09daf5e5c38dcd59128256a3ebc  <=  0;
                end else begin
                    Ibd8114af3027bd3364395e7b94484272  <=  ~I662d408ffd8fb9f249e531a167161429 + 1;
                    Ib312a09daf5e5c38dcd59128256a3ebc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7217d4790fec9797a1eb8cab1ebce71b == I5ea37c7893e55ef146fb831d8c09e87f ) begin
                    I49167fd9caea095581855b45b1f85d49  <= Ie95b8a5c2da6c0877d49c646c194f5b7;
                    Iaf3e2d448016a50829b4b0ea6f144b27  <=  0;
                end else begin
                    I49167fd9caea095581855b45b1f85d49  <=  ~Ie95b8a5c2da6c0877d49c646c194f5b7 + 1;
                    Iaf3e2d448016a50829b4b0ea6f144b27  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7217d4790fec9797a1eb8cab1ebce71b == Ic38315ea78c667a1f77a5fe34ac62412 ) begin
                    Ic502f151ee9ee01786e216d90a29403b  <= If940f33461f5e297e158db54f6aad610;
                    Iddbd5820346c3ea47bea79b2ee1ab7e5  <=  0;
                end else begin
                    Ic502f151ee9ee01786e216d90a29403b  <=  ~If940f33461f5e297e158db54f6aad610 + 1;
                    Iddbd5820346c3ea47bea79b2ee1ab7e5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3dd024db4130c105a6817e8a4935de0d == I2b954aae3ff5e2a0ce92a55107a86a46 ) begin
                    I25f89c7f7f11c7e2811913d6254dbc8c  <= I54aa9d4c6333d94970eae97aeb3603fa;
                    I1b024f329d24692f8d143aeeacfaf555  <=  0;
                end else begin
                    I25f89c7f7f11c7e2811913d6254dbc8c  <=  ~I54aa9d4c6333d94970eae97aeb3603fa + 1;
                    I1b024f329d24692f8d143aeeacfaf555  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3dd024db4130c105a6817e8a4935de0d == I958138e39e14c8fc1de83d02091b8f6e ) begin
                    I3f939889c013f740cc63c981d2ff85b2  <= Ib82fc62720e6346e1c05cc33d596447e;
                    I83f200ddde413f07bd296b8602aacdc7  <=  0;
                end else begin
                    I3f939889c013f740cc63c981d2ff85b2  <=  ~Ib82fc62720e6346e1c05cc33d596447e + 1;
                    I83f200ddde413f07bd296b8602aacdc7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3dd024db4130c105a6817e8a4935de0d == Idfd5a9e4c4cbd4ba9828220a7d021d28 ) begin
                    Ib0d2fc4f353a82d37bec9aa19a80475e  <= I24873624848b61f313865e10e77e35c6;
                    Ib4cec30021700f9f02847c2f1e0fc425  <=  0;
                end else begin
                    Ib0d2fc4f353a82d37bec9aa19a80475e  <=  ~I24873624848b61f313865e10e77e35c6 + 1;
                    Ib4cec30021700f9f02847c2f1e0fc425  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iae502e5a5ae518fb7b817afff28b7932 == Ied5041c527b4f04647dc80932b9ce7c4 ) begin
                    I2f19b77e5bb1b22b3cf5b1ace31ee6af  <= Icc3915d8325c22fc172f731553798fef;
                    I3cddf5a4ce875cb4e0c2fce7e36e5200  <=  0;
                end else begin
                    I2f19b77e5bb1b22b3cf5b1ace31ee6af  <=  ~Icc3915d8325c22fc172f731553798fef + 1;
                    I3cddf5a4ce875cb4e0c2fce7e36e5200  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iae502e5a5ae518fb7b817afff28b7932 == If6488c8e84e69a99816842a90c9578c2 ) begin
                    I283f82fd4a9700daca6ff1d16f747a09  <= I93b9837e63103431a0fdaf319a465c90;
                    I9c5d93dc3faea27b0f38898609b41545  <=  0;
                end else begin
                    I283f82fd4a9700daca6ff1d16f747a09  <=  ~I93b9837e63103431a0fdaf319a465c90 + 1;
                    I9c5d93dc3faea27b0f38898609b41545  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iae502e5a5ae518fb7b817afff28b7932 == Ic65f12c4a71f8c3af75f426128b333f9 ) begin
                    I8dc5483fb01a06ad8650e5fd4df30f49  <= I91237af3aa2af551dbbc626bb701215e;
                    I426a2f3c939a72ecff6a6314a19d52cb  <=  0;
                end else begin
                    I8dc5483fb01a06ad8650e5fd4df30f49  <=  ~I91237af3aa2af551dbbc626bb701215e + 1;
                    I426a2f3c939a72ecff6a6314a19d52cb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8b2b1d90204af5b100379ecad20fc0f == Ica6cd8bf97c702ae2541f682cc418a80 ) begin
                    I7e3f6b4bff19a0644c12fa4ef3667d84  <= Ib254d9701567f642d3586641edf85128;
                    I5919e3d3ea27d29a8093c52a6645959e  <=  0;
                end else begin
                    I7e3f6b4bff19a0644c12fa4ef3667d84  <=  ~Ib254d9701567f642d3586641edf85128 + 1;
                    I5919e3d3ea27d29a8093c52a6645959e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8b2b1d90204af5b100379ecad20fc0f == I73054b5829fd26eb2b09dc585f2c62f8 ) begin
                    Idf2371d30bec7ad5dea346a4a48a6e75  <= I25c50067a62d2b3599d15f12f89d384e;
                    I68c4ab26cc7c41ea3f9b8afec502bc42  <=  0;
                end else begin
                    Idf2371d30bec7ad5dea346a4a48a6e75  <=  ~I25c50067a62d2b3599d15f12f89d384e + 1;
                    I68c4ab26cc7c41ea3f9b8afec502bc42  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib8b2b1d90204af5b100379ecad20fc0f == I221be7886d94efc9e1ec553acd79dba4 ) begin
                    Ifd5a3069363cfc42e5a436856eeee708  <= I238be7f0e4a209a6b4201a024c8aed82;
                    Id4ea7f8c016571cc5a0af8327e2f95b9  <=  0;
                end else begin
                    Ifd5a3069363cfc42e5a436856eeee708  <=  ~I238be7f0e4a209a6b4201a024c8aed82 + 1;
                    Id4ea7f8c016571cc5a0af8327e2f95b9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idf0e651d0b13e167df3c0cc40d149c29 == I33557b5dddc36fe3625bf64e016c1c7e ) begin
                    I1a4e12577ac5e87d40bdcb54fe55818b  <= I233f5ddadd45c0df2108ea6c1d634f3c;
                    If6b109772fc17d898d70f75f538a0fdf  <=  0;
                end else begin
                    I1a4e12577ac5e87d40bdcb54fe55818b  <=  ~I233f5ddadd45c0df2108ea6c1d634f3c + 1;
                    If6b109772fc17d898d70f75f538a0fdf  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idf0e651d0b13e167df3c0cc40d149c29 == Ica7d3d482ec7dde7081b68988f76c9b4 ) begin
                    I1f1b6c20910c4f14999da6c9fdb4c349  <= I87a320ddaa1478146ff6e519dc65c40a;
                    I930235d80caaa415247c7fb380b3a134  <=  0;
                end else begin
                    I1f1b6c20910c4f14999da6c9fdb4c349  <=  ~I87a320ddaa1478146ff6e519dc65c40a + 1;
                    I930235d80caaa415247c7fb380b3a134  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Idf0e651d0b13e167df3c0cc40d149c29 == Ibf9561c2c5242296a3b607627e7e7989 ) begin
                    I1b0a200eea98f075f059d2a26b00f833  <= Ibf03d6940c0a38bef038a28b6a7b625d;
                    I324eeb4bf0e552118536fbd641189af1  <=  0;
                end else begin
                    I1b0a200eea98f075f059d2a26b00f833  <=  ~Ibf03d6940c0a38bef038a28b6a7b625d + 1;
                    I324eeb4bf0e552118536fbd641189af1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I89daaca029498d05ca62c095db439eb5 == Id0d621bef47b5c5735a4a999611a1c4a ) begin
                    Ie0dded072843efc1613cfe7136af37da  <= I90942470e2057e50ce4f5745ed68b81c;
                    I839160e07222b1f9f293efe22d68c168  <=  0;
                end else begin
                    Ie0dded072843efc1613cfe7136af37da  <=  ~I90942470e2057e50ce4f5745ed68b81c + 1;
                    I839160e07222b1f9f293efe22d68c168  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I89daaca029498d05ca62c095db439eb5 == I33cee0fcc65354655c9e57b3d43c11f2 ) begin
                    Ia6d6a867ebe63a8926d9affa4c15e376  <= I77fbc3f3b65962b610e39f4b085ecb7e;
                    I5244962685ce36dd805a7dc774c05d31  <=  0;
                end else begin
                    Ia6d6a867ebe63a8926d9affa4c15e376  <=  ~I77fbc3f3b65962b610e39f4b085ecb7e + 1;
                    I5244962685ce36dd805a7dc774c05d31  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I89daaca029498d05ca62c095db439eb5 == I8baad814c6bbc783645f574455b0f2d3 ) begin
                    Iddfc447b0c96056ae6e6434799ea00e9  <= I701845efaf1b02aefa381d4f6b45c401;
                    Ib92300e3d61e8a2bcaf0b2f40d4cb18f  <=  0;
                end else begin
                    Iddfc447b0c96056ae6e6434799ea00e9  <=  ~I701845efaf1b02aefa381d4f6b45c401 + 1;
                    Ib92300e3d61e8a2bcaf0b2f40d4cb18f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I89daaca029498d05ca62c095db439eb5 == Ib23a7e23bc223c7f3e83661811493229 ) begin
                    I36d03daaaaa37229d462f4bf5e521f73  <= Id446ddfd713c6e1592c562cfb123ea8b;
                    Id76c8bf8796c329353836a52e1dd74c3  <=  0;
                end else begin
                    I36d03daaaaa37229d462f4bf5e521f73  <=  ~Id446ddfd713c6e1592c562cfb123ea8b + 1;
                    Id76c8bf8796c329353836a52e1dd74c3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0fe5a34ceda936d0924efdd07fad11e5 == I55e8b1c375d49a1a1f044a4a60073d60 ) begin
                    I91e49319831eeee5dc75eac77ed8f8a3  <= If4f752779d27392e7536565d425bce25;
                    Ibb163802022194494881194dc6b49c2d  <=  0;
                end else begin
                    I91e49319831eeee5dc75eac77ed8f8a3  <=  ~If4f752779d27392e7536565d425bce25 + 1;
                    Ibb163802022194494881194dc6b49c2d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0fe5a34ceda936d0924efdd07fad11e5 == I023853b98208afd9bcb1ff63abb91b2e ) begin
                    I4e9f03752b041491ae2bc40fbd2b8d43  <= If112169057d6293326a56443ac3cf517;
                    Iedb3b8bfd024408f08a2b377956239af  <=  0;
                end else begin
                    I4e9f03752b041491ae2bc40fbd2b8d43  <=  ~If112169057d6293326a56443ac3cf517 + 1;
                    Iedb3b8bfd024408f08a2b377956239af  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0fe5a34ceda936d0924efdd07fad11e5 == Icd656c959fe941e863db11f02d3c514e ) begin
                    I9a71e50dac7ad707a4b0946ebc1fe6d4  <= I78f727f8d85b5d7f0ffa57f02538f939;
                    I6cfe7ce048413c7c959a0eefe967885b  <=  0;
                end else begin
                    I9a71e50dac7ad707a4b0946ebc1fe6d4  <=  ~I78f727f8d85b5d7f0ffa57f02538f939 + 1;
                    I6cfe7ce048413c7c959a0eefe967885b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0fe5a34ceda936d0924efdd07fad11e5 == I06cea262d84c35f3e6a1b6690b82cbf8 ) begin
                    I8220d15825d6bac07d773ff0db2f9795  <= I01ec629f60c17c2251f977205234cd44;
                    I664a362c93dd438aec485063a6f0c7de  <=  0;
                end else begin
                    I8220d15825d6bac07d773ff0db2f9795  <=  ~I01ec629f60c17c2251f977205234cd44 + 1;
                    I664a362c93dd438aec485063a6f0c7de  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7876cbb2b5d8aba3652ec8b218080dff == I1d7bbe81db5320829eb5b29252fc6cf2 ) begin
                    I6b2dc98acc78a1151dd6670ed981d839  <= I23f774adb64807c0edaa9941c75651b6;
                    I9252e19b54173ae2a9d0815dfc46eec2  <=  0;
                end else begin
                    I6b2dc98acc78a1151dd6670ed981d839  <=  ~I23f774adb64807c0edaa9941c75651b6 + 1;
                    I9252e19b54173ae2a9d0815dfc46eec2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7876cbb2b5d8aba3652ec8b218080dff == Iafad27be14640dbdcff055b7e34f6467 ) begin
                    Ie371be4323965591a5786063ba028ce1  <= I2361ef4fd70e4c05b25289d0845564c4;
                    I2ea93b2142eee9f44c8e7bf892bf02ab  <=  0;
                end else begin
                    Ie371be4323965591a5786063ba028ce1  <=  ~I2361ef4fd70e4c05b25289d0845564c4 + 1;
                    I2ea93b2142eee9f44c8e7bf892bf02ab  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7876cbb2b5d8aba3652ec8b218080dff == Idfd58540bb8d1465514c3c843d303825 ) begin
                    Ic4985251ed9f9120d2232ec96949831b  <= Ic3067b434ca17be7bad595e1f9b822c5;
                    I6772834728b2e641c6e3c14cda255ad6  <=  0;
                end else begin
                    Ic4985251ed9f9120d2232ec96949831b  <=  ~Ic3067b434ca17be7bad595e1f9b822c5 + 1;
                    I6772834728b2e641c6e3c14cda255ad6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7876cbb2b5d8aba3652ec8b218080dff == I7c98a5f1ea935e4de159795b5dd795ed ) begin
                    I6015d64c067415fe216d90a5be409e33  <= I3546ddbae9c9db4517802db56cee35f0;
                    Id6a64c33b3beb88abcadc06af18e1858  <=  0;
                end else begin
                    I6015d64c067415fe216d90a5be409e33  <=  ~I3546ddbae9c9db4517802db56cee35f0 + 1;
                    Id6a64c33b3beb88abcadc06af18e1858  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If692ff56ce90d22d7af881599c54df75 == I84b1e71a64cd4d96c44444e337dde784 ) begin
                    If6f304fe091216273270713c6b6e8a6d  <= I35e91092ed503831ed818f36a1ce1537;
                    Ib89f2aee80d36f4e473d1a1046e836dd  <=  0;
                end else begin
                    If6f304fe091216273270713c6b6e8a6d  <=  ~I35e91092ed503831ed818f36a1ce1537 + 1;
                    Ib89f2aee80d36f4e473d1a1046e836dd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If692ff56ce90d22d7af881599c54df75 == I609aef4d51d5d190deea41f71ef0403c ) begin
                    I779ee6daefe3c5c96548dc5e0ba83bd3  <= I973f185cf29e13193abf0108d4faa9d1;
                    I78aeec1644701502f6f71c64341274ab  <=  0;
                end else begin
                    I779ee6daefe3c5c96548dc5e0ba83bd3  <=  ~I973f185cf29e13193abf0108d4faa9d1 + 1;
                    I78aeec1644701502f6f71c64341274ab  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If692ff56ce90d22d7af881599c54df75 == I68a99adfa01586d1ad7bdeb282f11d87 ) begin
                    Ieef21b505cc215387f8930888062b767  <= Iee58b0442a6cccf0990ebb551b47fa92;
                    I9a09fda6e73783a7c9a4582fec8121b4  <=  0;
                end else begin
                    Ieef21b505cc215387f8930888062b767  <=  ~Iee58b0442a6cccf0990ebb551b47fa92 + 1;
                    I9a09fda6e73783a7c9a4582fec8121b4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If692ff56ce90d22d7af881599c54df75 == I1f68aed9a1379bbbd2c531fc0df392fe ) begin
                    Icbabacaecbbac74901402e5e5874328b  <= I2cb3207a5c1b25386ac7eb532955f260;
                    I9db6919efaef0952b84eaf8e71f77777  <=  0;
                end else begin
                    Icbabacaecbbac74901402e5e5874328b  <=  ~I2cb3207a5c1b25386ac7eb532955f260 + 1;
                    I9db6919efaef0952b84eaf8e71f77777  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I18a7a4fe8931c79df3a69223af46c440 == Ib1cbee37b3fad49ab5805647ccf95b7b ) begin
                    I6ec13a161f7f1a0f57e9ba4998474954  <= Icd4f07bc30c66f7f5b431ed97e7ac7b6;
                    I5a4646a8adf0ed43a905fd4ee84d85bd  <=  0;
                end else begin
                    I6ec13a161f7f1a0f57e9ba4998474954  <=  ~Icd4f07bc30c66f7f5b431ed97e7ac7b6 + 1;
                    I5a4646a8adf0ed43a905fd4ee84d85bd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I18a7a4fe8931c79df3a69223af46c440 == Ibbe9c1e2c9f2c0b00e4be25205a824d6 ) begin
                    I71f9823e92c51be2e9a050d01e63902d  <= Ifec6f3a1e10144acb320d5d502ed1ea3;
                    I1e3444ee88dc52881397d266f469b45c  <=  0;
                end else begin
                    I71f9823e92c51be2e9a050d01e63902d  <=  ~Ifec6f3a1e10144acb320d5d502ed1ea3 + 1;
                    I1e3444ee88dc52881397d266f469b45c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I18a7a4fe8931c79df3a69223af46c440 == I6c7e0e56cd76e03261638e924f90377e ) begin
                    Ia0037030d79400734732f061fd81edf6  <= Ic87bff64a597e6d02583041b552328ee;
                    I3c42e969e5e4b99f1f2eaa01419d4ed9  <=  0;
                end else begin
                    Ia0037030d79400734732f061fd81edf6  <=  ~Ic87bff64a597e6d02583041b552328ee + 1;
                    I3c42e969e5e4b99f1f2eaa01419d4ed9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I18a7a4fe8931c79df3a69223af46c440 == I676d7f8a89fbbef4b067d07264ae427c ) begin
                    Id796584e3e7af67536a27f7299b71916  <= I489f21ef8243ef8caa1c29f034c3e2ac;
                    I9210d06734058f76e7a5a470dbe6e74b  <=  0;
                end else begin
                    Id796584e3e7af67536a27f7299b71916  <=  ~I489f21ef8243ef8caa1c29f034c3e2ac + 1;
                    I9210d06734058f76e7a5a470dbe6e74b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I8eec3538b8cc9c046954b6804cc656b0 == Ifcaf093fbbec17632ca0050583df41c4 ) begin
                    Iec938bc1bbad930fade05d74c10989a3  <= I773901563077961acada85962209d68a;
                    I2b35c8fa7c947b3e7691cdcab0c5a7a7  <=  0;
                end else begin
                    Iec938bc1bbad930fade05d74c10989a3  <=  ~I773901563077961acada85962209d68a + 1;
                    I2b35c8fa7c947b3e7691cdcab0c5a7a7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I8eec3538b8cc9c046954b6804cc656b0 == Ia358ae5a96e63f3bb5c6bb34f263c387 ) begin
                    I2a7a7c5eabd1623c1c3d4bd93bf18617  <= Ifbd176fe3e78bc2dc2e0e77ba3ccd2d0;
                    Id58d1af007bb5858499af71a43e6574f  <=  0;
                end else begin
                    I2a7a7c5eabd1623c1c3d4bd93bf18617  <=  ~Ifbd176fe3e78bc2dc2e0e77ba3ccd2d0 + 1;
                    Id58d1af007bb5858499af71a43e6574f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I8eec3538b8cc9c046954b6804cc656b0 == Ib1e4443484bfc289563a8b7d9b1c86b6 ) begin
                    I71cfc7fd85636c5554b9fe9f9ba8e3aa  <= I53f68a4cb81c71ee7bd6f61171b7478d;
                    I12e92aa9c9ca2135f7ba879d82ad615b  <=  0;
                end else begin
                    I71cfc7fd85636c5554b9fe9f9ba8e3aa  <=  ~I53f68a4cb81c71ee7bd6f61171b7478d + 1;
                    I12e92aa9c9ca2135f7ba879d82ad615b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I8eec3538b8cc9c046954b6804cc656b0 == Ib3baee13e51f9fb8c39d04211497e274 ) begin
                    I4c8ae97548bc3dbf3e3621f80c3e0835  <= I7568ec59f1359bedce86dbc6af50df71;
                    If32ea54eb47d27e35a81aa4b9e1f7713  <=  0;
                end else begin
                    I4c8ae97548bc3dbf3e3621f80c3e0835  <=  ~I7568ec59f1359bedce86dbc6af50df71 + 1;
                    If32ea54eb47d27e35a81aa4b9e1f7713  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I653767e659590c1676edf6c25fc0e253 == Ic24de5d8c9148fab7b9dcac9d8996740 ) begin
                    Iaa93c760705c984a0eea90d41a6c049b  <= Id2bf82d6bf0a201f80a58357038a0992;
                    Ib1ddab09d1a726176414e4a877b66e3f  <=  0;
                end else begin
                    Iaa93c760705c984a0eea90d41a6c049b  <=  ~Id2bf82d6bf0a201f80a58357038a0992 + 1;
                    Ib1ddab09d1a726176414e4a877b66e3f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I653767e659590c1676edf6c25fc0e253 == I46489795c1a8e178f1b2d40711655c44 ) begin
                    I2acc73851f8a803e69c0f1865e00f46e  <= I22442354ca2b77306f25839ce6124699;
                    Id3838f634ce2d90a19622185391ba868  <=  0;
                end else begin
                    I2acc73851f8a803e69c0f1865e00f46e  <=  ~I22442354ca2b77306f25839ce6124699 + 1;
                    Id3838f634ce2d90a19622185391ba868  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I653767e659590c1676edf6c25fc0e253 == If39c47fd6b6913ec7946018145d31945 ) begin
                    I928333e9cc75d49fa6f7094e49631123  <= I71a5c2876a07d8edd001ef2d108e59c1;
                    Ia3f429c43f23f4f057abed98cfa94748  <=  0;
                end else begin
                    I928333e9cc75d49fa6f7094e49631123  <=  ~I71a5c2876a07d8edd001ef2d108e59c1 + 1;
                    Ia3f429c43f23f4f057abed98cfa94748  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I653767e659590c1676edf6c25fc0e253 == Ie336a92376f51b145c60f935b8fd0f8c ) begin
                    Idf02dd4b7e8a6958913e6180fec1feee  <= Iaf333aa6b135927cf1ad1f76298ccd63;
                    I62b423a6061215d16871bfdf9a9cdbd2  <=  0;
                end else begin
                    Idf02dd4b7e8a6958913e6180fec1feee  <=  ~Iaf333aa6b135927cf1ad1f76298ccd63 + 1;
                    I62b423a6061215d16871bfdf9a9cdbd2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5ff863be142b92dff89f7916d0d088c1 == Ia6f981e46e3d7ead096d73154e97dca9 ) begin
                    Ib30cc7931858974728d92eb68890449f  <= Ia71cfd8cf9bea4e600ea204e41271c7d;
                    I17f82f6daa8a92f1da5a1952a558ad7e  <=  0;
                end else begin
                    Ib30cc7931858974728d92eb68890449f  <=  ~Ia71cfd8cf9bea4e600ea204e41271c7d + 1;
                    I17f82f6daa8a92f1da5a1952a558ad7e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5ff863be142b92dff89f7916d0d088c1 == If7593819b136ad3db74d793e5a0f18c3 ) begin
                    Ia504dbcee6e5894fed83371bf70b2d44  <= I164b032929ac2b8cf1a6672859639a30;
                    Ie0e9f7c1d69d8930f8452d3618512877  <=  0;
                end else begin
                    Ia504dbcee6e5894fed83371bf70b2d44  <=  ~I164b032929ac2b8cf1a6672859639a30 + 1;
                    Ie0e9f7c1d69d8930f8452d3618512877  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5ff863be142b92dff89f7916d0d088c1 == I0b480fa6fe571ea7d25d13f8f1ba26da ) begin
                    I32b4e50b8acefe1c108d777da565f4ed  <= I2ef0447f5c64fd5c65e23c16069a62ef;
                    Id9de214d84792861772ef396b5b9208f  <=  0;
                end else begin
                    I32b4e50b8acefe1c108d777da565f4ed  <=  ~I2ef0447f5c64fd5c65e23c16069a62ef + 1;
                    Id9de214d84792861772ef396b5b9208f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I5ff863be142b92dff89f7916d0d088c1 == I66ab48b076a0e2006d1f4741e15f3c36 ) begin
                    If9fd1d8c0c13042a6f2d258478b63925  <= Ide7008ee7f1fba156dc6145b3505e553;
                    I027f018e60dda98666458cb69a6e4be2  <=  0;
                end else begin
                    If9fd1d8c0c13042a6f2d258478b63925  <=  ~Ide7008ee7f1fba156dc6145b3505e553 + 1;
                    I027f018e60dda98666458cb69a6e4be2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I49f9fd0e0719be527f2a54814dab83ea == I9e397fd8cfd4ee1b9cd3cccbd4c03005 ) begin
                    Iccb437017198e4421ab51d74aed779f0  <= I129a7ced6bc6f48f20fa552e2519925c;
                    I996821515569c215f3f688d91dee8abe  <=  0;
                end else begin
                    Iccb437017198e4421ab51d74aed779f0  <=  ~I129a7ced6bc6f48f20fa552e2519925c + 1;
                    I996821515569c215f3f688d91dee8abe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I49f9fd0e0719be527f2a54814dab83ea == I177684367c872f5a3df89c0d2bb95434 ) begin
                    Id10bf2bf52a8f1be9eeafcefd6dd5dcb  <= I67123cf825352e52cf0158060ad69a13;
                    I6f617bfa2700fb385d425f6b4581f594  <=  0;
                end else begin
                    Id10bf2bf52a8f1be9eeafcefd6dd5dcb  <=  ~I67123cf825352e52cf0158060ad69a13 + 1;
                    I6f617bfa2700fb385d425f6b4581f594  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I49f9fd0e0719be527f2a54814dab83ea == Icdb37cf629ec16db879e288eba5ef9a9 ) begin
                    Ie590c921147b7252d2605f7712dfe437  <= I09923d784a9f9625a37221f639537941;
                    Id5f8b6b344dc8e629f13e5d157f510cb  <=  0;
                end else begin
                    Ie590c921147b7252d2605f7712dfe437  <=  ~I09923d784a9f9625a37221f639537941 + 1;
                    Id5f8b6b344dc8e629f13e5d157f510cb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I945f2476eb599844cbee0cd89038e392 == I225d035b7f8d13e9895ca60f3da8bf90 ) begin
                    I178ed883c28bbf3e1ab05cb95f62b343  <= I5947be93fdb18bf0ad341fb826c9e6d7;
                    I579a5dc98f16e0c5d52fc7958586a8d5  <=  0;
                end else begin
                    I178ed883c28bbf3e1ab05cb95f62b343  <=  ~I5947be93fdb18bf0ad341fb826c9e6d7 + 1;
                    I579a5dc98f16e0c5d52fc7958586a8d5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I945f2476eb599844cbee0cd89038e392 == Ia3572b856ec1a14e316444c2f15ac9a5 ) begin
                    I01971a175615a422d264805252f91f3b  <= I08621ee033cd49702ad08af4d31eb999;
                    I0f2769698735ab28df30370c3c8b56cc  <=  0;
                end else begin
                    I01971a175615a422d264805252f91f3b  <=  ~I08621ee033cd49702ad08af4d31eb999 + 1;
                    I0f2769698735ab28df30370c3c8b56cc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I945f2476eb599844cbee0cd89038e392 == I2c927c7ee3628a78f48c6099d2036959 ) begin
                    Ie770c4567f35b40c46ccbda059e6d3a8  <= Id5eca60b22d3835119571fe4b1a03479;
                    I9fbc79fd7be52757770dce6e04749b4f  <=  0;
                end else begin
                    Ie770c4567f35b40c46ccbda059e6d3a8  <=  ~Id5eca60b22d3835119571fe4b1a03479 + 1;
                    I9fbc79fd7be52757770dce6e04749b4f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied0c5f8a9243cd9d93672ad6cc907d21 == I578551b6331fffa97a6d05652e406e3f ) begin
                    I25975702f0b9c0baf586fe471676dfea  <= I7267ba2b9cb511a48a3a7044e854f7da;
                    Idfe33235c2f93ac311da89ba63e0f1c5  <=  0;
                end else begin
                    I25975702f0b9c0baf586fe471676dfea  <=  ~I7267ba2b9cb511a48a3a7044e854f7da + 1;
                    Idfe33235c2f93ac311da89ba63e0f1c5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied0c5f8a9243cd9d93672ad6cc907d21 == I6f301798efb2c67ea363df40f2fe340f ) begin
                    Id2ef737d910326394b68eaa0833bfccb  <= I5893fa21ec8bbdcea9677cc12fc4057a;
                    Ic46d706f6be34cb4133a4128567837d3  <=  0;
                end else begin
                    Id2ef737d910326394b68eaa0833bfccb  <=  ~I5893fa21ec8bbdcea9677cc12fc4057a + 1;
                    Ic46d706f6be34cb4133a4128567837d3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied0c5f8a9243cd9d93672ad6cc907d21 == I744d142b9316b9f8937563c1023882e6 ) begin
                    I577cd1f9ad512ec10f5008165f2e4a74  <= I564896fe01ec799a0fbe790473753559;
                    Ibb3c635f2e62a63c9bdb150b3cda7155  <=  0;
                end else begin
                    I577cd1f9ad512ec10f5008165f2e4a74  <=  ~I564896fe01ec799a0fbe790473753559 + 1;
                    Ibb3c635f2e62a63c9bdb150b3cda7155  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9134c7f579723c7615af60b4344efe76 == Id7fa5f9fb6059439297f246cb228cc02 ) begin
                    I1de8f87eb39276e073f5804b1df3b67a  <= If279ab7c515c4039c8272b913c2fa107;
                    I7bdfb2d2b7dd18fc7c0d43b708fb1e35  <=  0;
                end else begin
                    I1de8f87eb39276e073f5804b1df3b67a  <=  ~If279ab7c515c4039c8272b913c2fa107 + 1;
                    I7bdfb2d2b7dd18fc7c0d43b708fb1e35  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9134c7f579723c7615af60b4344efe76 == I18e9dd5583f3ac91451a4e75f0d5d474 ) begin
                    I7f8e7928e6caeac14f787d7e0b6a47df  <= Ib61705ff5820f531eb17c40ed05f6ec3;
                    I42a1cd616514a1c7384d07095e6b2d70  <=  0;
                end else begin
                    I7f8e7928e6caeac14f787d7e0b6a47df  <=  ~Ib61705ff5820f531eb17c40ed05f6ec3 + 1;
                    I42a1cd616514a1c7384d07095e6b2d70  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9134c7f579723c7615af60b4344efe76 == I64afac5bd1ea7a2ab696e630cc3ad162 ) begin
                    Ia7048aa3f949b0b2e54ab900efe01131  <= I50149e5de41ca2998c4e8cc4b19e166b;
                    I19a91106f189ef43ee50edab49d297c1  <=  0;
                end else begin
                    Ia7048aa3f949b0b2e54ab900efe01131  <=  ~I50149e5de41ca2998c4e8cc4b19e166b + 1;
                    I19a91106f189ef43ee50edab49d297c1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 == I0b3bfd6ce482cfb20d461862a0bf8f61 ) begin
                    I1fcbb73d165eab038c745fac370fd68f  <= Id40cac3272643f3f91b73c6aa1740f3b;
                    I90088e4928092e62e193039faf154240  <=  0;
                end else begin
                    I1fcbb73d165eab038c745fac370fd68f  <=  ~Id40cac3272643f3f91b73c6aa1740f3b + 1;
                    I90088e4928092e62e193039faf154240  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 == I16119df9372ce61c0c8600ddba36e607 ) begin
                    Ia822cd52015d599bc45ae7338b4e88e1  <= Ic63eee2d700493c41ee2d186ff7111b9;
                    Ic0fed8f997e03bcca119270589f8bf0a  <=  0;
                end else begin
                    Ia822cd52015d599bc45ae7338b4e88e1  <=  ~Ic63eee2d700493c41ee2d186ff7111b9 + 1;
                    Ic0fed8f997e03bcca119270589f8bf0a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 == I0957a6c9a87bc89dd9748491807837af ) begin
                    I56b85e2d5a7259eb50fa983b92d8b160  <= I51de42598e0df4a76cf7b02c61ae9550;
                    I3ba811abe28766d976a2afd02c22fc76  <=  0;
                end else begin
                    I56b85e2d5a7259eb50fa983b92d8b160  <=  ~I51de42598e0df4a76cf7b02c61ae9550 + 1;
                    I3ba811abe28766d976a2afd02c22fc76  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 == I12f8c91d67e31e11033d5b3b266c659b ) begin
                    I1d23632f8e8f66a30b4ef6c76aae3ece  <= Ia89a1a58f6327ee3c105cae860942171;
                    I66463d17d0fcb691e727568e4d55ae43  <=  0;
                end else begin
                    I1d23632f8e8f66a30b4ef6c76aae3ece  <=  ~Ia89a1a58f6327ee3c105cae860942171 + 1;
                    I66463d17d0fcb691e727568e4d55ae43  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie92388a9d1e71d73c07ed86e9bf6c887 == I690b96154d7717bf62eeb740b10ce6d5 ) begin
                    Ib578de11f0407cfeb0dac68bd5fbf7a0  <= Ib149a5872e31cd5df77b66298b4aad12;
                    Icf73bfd92fe6265b8e7d9b2439573a96  <=  0;
                end else begin
                    Ib578de11f0407cfeb0dac68bd5fbf7a0  <=  ~Ib149a5872e31cd5df77b66298b4aad12 + 1;
                    Icf73bfd92fe6265b8e7d9b2439573a96  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 == I25b3993479d7cc172ba6a480628b9188 ) begin
                    I08879fb80c58de5fb2bf547ce013c67f  <= Iaa16c14572ad0442eb3c58a97bef5ada;
                    I7c3f7076072ee81960c8b0187648eb41  <=  0;
                end else begin
                    I08879fb80c58de5fb2bf547ce013c67f  <=  ~Iaa16c14572ad0442eb3c58a97bef5ada + 1;
                    I7c3f7076072ee81960c8b0187648eb41  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 == I7f3a220cdbf5bf1737690e1719f888e5 ) begin
                    I8f7c4c602b7de5d9a401d3933a7e50a8  <= I88d5d48e05b1c9a6d8060f58917e3834;
                    I68ccb34c409f89f1a2872d64f85e3245  <=  0;
                end else begin
                    I8f7c4c602b7de5d9a401d3933a7e50a8  <=  ~I88d5d48e05b1c9a6d8060f58917e3834 + 1;
                    I68ccb34c409f89f1a2872d64f85e3245  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 == I8d068dee7478a9f899c8145ef6d824a5 ) begin
                    I2ab4cc1ef6b743cda8765a22e28fd7a7  <= I4269e18c2df4d39c683ffb7d01a08322;
                    I069661eba4d8f68a4e5c78e99e9355e8  <=  0;
                end else begin
                    I2ab4cc1ef6b743cda8765a22e28fd7a7  <=  ~I4269e18c2df4d39c683ffb7d01a08322 + 1;
                    I069661eba4d8f68a4e5c78e99e9355e8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 == I2286af8d6007a7da5c745d75f407b5d9 ) begin
                    Idc58a89f7d8ee884b198b6e4752ec58f  <= Ia29017fa9327fdaa7c10b2797f8aa6ec;
                    I6cc756f9cb1020c8045872d628b771f8  <=  0;
                end else begin
                    Idc58a89f7d8ee884b198b6e4752ec58f  <=  ~Ia29017fa9327fdaa7c10b2797f8aa6ec + 1;
                    I6cc756f9cb1020c8045872d628b771f8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I6804fecdf59233c6cf14409bf2f1e430 == I214f77e05ac2ce4b94d4c5e53675717d ) begin
                    If9c0f4c64c7648e509077df16c14b7a1  <= Ia142ac799256541fe33f898a6a31dd71;
                    I95494fb67de54f6055f54c7568106488  <=  0;
                end else begin
                    If9c0f4c64c7648e509077df16c14b7a1  <=  ~Ia142ac799256541fe33f898a6a31dd71 + 1;
                    I95494fb67de54f6055f54c7568106488  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9e777a342bf53eaba0280737ae404bc1 == I8fc900d4110bc862ad7287255dddf2f0 ) begin
                    I8cc434418203702ad5a21eb4f0340dc5  <= I4c039794243933a9bb7ad6db7eda6a87;
                    Ibbfab9efcd61f23b09e371554c0778b0  <=  0;
                end else begin
                    I8cc434418203702ad5a21eb4f0340dc5  <=  ~I4c039794243933a9bb7ad6db7eda6a87 + 1;
                    Ibbfab9efcd61f23b09e371554c0778b0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9e777a342bf53eaba0280737ae404bc1 == If609e068414eed49fbe97f86e2546768 ) begin
                    Iee9d96f800fc848f3c4b6b6901a72623  <= I0debb3ed4f9540c162cd525588e0ae3f;
                    Ibb2a246712268d6d8a0ad0354b8e611f  <=  0;
                end else begin
                    Iee9d96f800fc848f3c4b6b6901a72623  <=  ~I0debb3ed4f9540c162cd525588e0ae3f + 1;
                    Ibb2a246712268d6d8a0ad0354b8e611f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9e777a342bf53eaba0280737ae404bc1 == I69177c754e87bc42401bccf54b770358 ) begin
                    I989036e56c9c7386279e83ae83ad4f7d  <= I681eed68ee814fb18fd794207d9266e1;
                    Ie9f5d2f06f60d7f436118f2c92695107  <=  0;
                end else begin
                    I989036e56c9c7386279e83ae83ad4f7d  <=  ~I681eed68ee814fb18fd794207d9266e1 + 1;
                    Ie9f5d2f06f60d7f436118f2c92695107  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9e777a342bf53eaba0280737ae404bc1 == I3b121702ca62507c2afda1ed93183499 ) begin
                    Icf23ca0439c76198fe647a0b785d9503  <= Ic260784b8910f5a0483afee9b68efb31;
                    I0ee25f335a84b7a190ccd690fccc1fce  <=  0;
                end else begin
                    Icf23ca0439c76198fe647a0b785d9503  <=  ~Ic260784b8910f5a0483afee9b68efb31 + 1;
                    I0ee25f335a84b7a190ccd690fccc1fce  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9e777a342bf53eaba0280737ae404bc1 == Id979aeb39d36400b85386a8e96ca5a35 ) begin
                    I406bddf2c4a4b6e6aedb86d72f14994f  <= I22cd2d30a7684002cacca4deae4c95a0;
                    Ica83129589b16c7392387bcddd9e81e9  <=  0;
                end else begin
                    I406bddf2c4a4b6e6aedb86d72f14994f  <=  ~I22cd2d30a7684002cacca4deae4c95a0 + 1;
                    Ica83129589b16c7392387bcddd9e81e9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied53820aab06b5c3423b1d878c71948f == I61ca2dba668792ee6a83850e2f118eb0 ) begin
                    I5331e97930599788b1df06992c5e4a5c  <= I136b4136d582f9fad21f90297cfafea3;
                    I91fc1c1758eb8c136744c1ef47785b49  <=  0;
                end else begin
                    I5331e97930599788b1df06992c5e4a5c  <=  ~I136b4136d582f9fad21f90297cfafea3 + 1;
                    I91fc1c1758eb8c136744c1ef47785b49  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied53820aab06b5c3423b1d878c71948f == I7e7f1d73e81031a38992b4f9a3f90717 ) begin
                    I98577e71126ac9bdbe4359101d4d48d7  <= Id8d6be9677d3b0ceca26b3b671757c2c;
                    I2bede76feb8d499cef693a3cc0bb95f4  <=  0;
                end else begin
                    I98577e71126ac9bdbe4359101d4d48d7  <=  ~Id8d6be9677d3b0ceca26b3b671757c2c + 1;
                    I2bede76feb8d499cef693a3cc0bb95f4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied53820aab06b5c3423b1d878c71948f == I029dbf330bab56469b88cbd602e8e16b ) begin
                    I696f551b6f96d0f7d27eb685bd374229  <= I6a93f928c104ea211dcc8a461506327d;
                    Ia0d9b7bd503ddeeefe9d0646c1f4e6d8  <=  0;
                end else begin
                    I696f551b6f96d0f7d27eb685bd374229  <=  ~I6a93f928c104ea211dcc8a461506327d + 1;
                    Ia0d9b7bd503ddeeefe9d0646c1f4e6d8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied53820aab06b5c3423b1d878c71948f == I47ddb6cfe64c5addb3900e193094ac8f ) begin
                    I1aa256ab19406597846ff353b65224cb  <= I240da147648bec33195a5f5c273fc6f4;
                    I2af1f93bd1d85a66028ef0add7a69962  <=  0;
                end else begin
                    I1aa256ab19406597846ff353b65224cb  <=  ~I240da147648bec33195a5f5c273fc6f4 + 1;
                    I2af1f93bd1d85a66028ef0add7a69962  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied53820aab06b5c3423b1d878c71948f == Ibdf7e609b7e42c57450d9d9fdd610881 ) begin
                    I00f1b24291a0e8496e13fe076e377cb8  <= I55494d0e8454e3cbb4158559e0d29984;
                    Icc568348313201d6814f92694d7db06f  <=  0;
                end else begin
                    I00f1b24291a0e8496e13fe076e377cb8  <=  ~I55494d0e8454e3cbb4158559e0d29984 + 1;
                    Icc568348313201d6814f92694d7db06f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24cceded372d782c67b33f3a78b16045 == Ia096e8920afb814330e53778c955f8b0 ) begin
                    Ie6f40dc356120aeb6cfa7a3fb5fae8cc  <= Ied3cc579b3cf126081acf8e1117007cf;
                    Iba815b719f813a245efb2627660634ff  <=  0;
                end else begin
                    Ie6f40dc356120aeb6cfa7a3fb5fae8cc  <=  ~Ied3cc579b3cf126081acf8e1117007cf + 1;
                    Iba815b719f813a245efb2627660634ff  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24cceded372d782c67b33f3a78b16045 == I365fd3d16d984516e33a7b68338d0384 ) begin
                    I67e23e6286edc4e01a7ebdace62ce56d  <= I76140bdc374dd6031097575fd231b468;
                    Id67d39730eb990c4b125cfa772e27e3a  <=  0;
                end else begin
                    I67e23e6286edc4e01a7ebdace62ce56d  <=  ~I76140bdc374dd6031097575fd231b468 + 1;
                    Id67d39730eb990c4b125cfa772e27e3a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24cceded372d782c67b33f3a78b16045 == I5e86c33e58b50627d7e69a4200525e05 ) begin
                    Id2c7c6d20146edcca65120c025e25a0a  <= I650345d21e5c2e7a9bf1810630161089;
                    Ib09008d80ae9d6708371c0c40f157656  <=  0;
                end else begin
                    Id2c7c6d20146edcca65120c025e25a0a  <=  ~I650345d21e5c2e7a9bf1810630161089 + 1;
                    Ib09008d80ae9d6708371c0c40f157656  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2e78d36bca5bfb016af674c343f9c041 == I52ef2681091d643e4ed026581feeb3f2 ) begin
                    Ida1e2d8b0e45e14c4c669c8b9d6947f5  <= Ie852635f073dc918e7b1075ffad46f24;
                    Id61b17db82e540f939ed8a4c3b596278  <=  0;
                end else begin
                    Ida1e2d8b0e45e14c4c669c8b9d6947f5  <=  ~Ie852635f073dc918e7b1075ffad46f24 + 1;
                    Id61b17db82e540f939ed8a4c3b596278  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2e78d36bca5bfb016af674c343f9c041 == I0e30717ed1e983e1c5af25037d5cfca3 ) begin
                    I1fd443d00410d0577eef9f1f26e64700  <= I9ec80c14eb5f0f305e1a9e6107a6001e;
                    I24868694c2523bb657da19c2e84ec8ef  <=  0;
                end else begin
                    I1fd443d00410d0577eef9f1f26e64700  <=  ~I9ec80c14eb5f0f305e1a9e6107a6001e + 1;
                    I24868694c2523bb657da19c2e84ec8ef  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I2e78d36bca5bfb016af674c343f9c041 == I640e720e6aaa2f8e14b5dacd51cc6e66 ) begin
                    I9ea760f08ba7b84fcaad929a3669450d  <= I80ba56447ab19b33610c23105b0b1637;
                    I9dcf88e53c655bce8190c5e85f5ca777  <=  0;
                end else begin
                    I9ea760f08ba7b84fcaad929a3669450d  <=  ~I80ba56447ab19b33610c23105b0b1637 + 1;
                    I9dcf88e53c655bce8190c5e85f5ca777  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I17a9a995de58643dbbfb78604f26198b == I81f4ac1f01d8170f427ee5ef89e8bd78 ) begin
                    Ia522420603dbde92a49da297554ede5e  <= Ib9132d9fa7180c3fcbacb7c570d6b0f2;
                    Ib881ec4b6a6de42dfcb2be830ca39ac8  <=  0;
                end else begin
                    Ia522420603dbde92a49da297554ede5e  <=  ~Ib9132d9fa7180c3fcbacb7c570d6b0f2 + 1;
                    Ib881ec4b6a6de42dfcb2be830ca39ac8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I17a9a995de58643dbbfb78604f26198b == I8319f97640191977a9b89e7639aee739 ) begin
                    I9be575cacaafcc13a0306545be56a04d  <= I01621f113f636a9caf9b5ca0bb20ef77;
                    Ifd2ece02d5ffb0a50d8b151a8fa8e703  <=  0;
                end else begin
                    I9be575cacaafcc13a0306545be56a04d  <=  ~I01621f113f636a9caf9b5ca0bb20ef77 + 1;
                    Ifd2ece02d5ffb0a50d8b151a8fa8e703  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I17a9a995de58643dbbfb78604f26198b == I21add24f8eed563787b8567fe43947f8 ) begin
                    Ieb9a03ad2c7c7df356477e8b4224ebd9  <= I3eeddb549c6e1f07469c0e0dca68be92;
                    I7da3a787760c42ef510ece8234c020a8  <=  0;
                end else begin
                    Ieb9a03ad2c7c7df356477e8b4224ebd9  <=  ~I3eeddb549c6e1f07469c0e0dca68be92 + 1;
                    I7da3a787760c42ef510ece8234c020a8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iad642c4c62766e8f8bd5a1e9e73bdc80 == I1a772b29d533c44422332cf291d27253 ) begin
                    If7f263cb2fb7fd35682d44c42639bab6  <= Ibe664dd203ed4162abcd36eb8d57bfa6;
                    I2204fa0d852e56e843393b3959f3df72  <=  0;
                end else begin
                    If7f263cb2fb7fd35682d44c42639bab6  <=  ~Ibe664dd203ed4162abcd36eb8d57bfa6 + 1;
                    I2204fa0d852e56e843393b3959f3df72  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iad642c4c62766e8f8bd5a1e9e73bdc80 == I8ec002e0ccc2cee9a210b987bf1cccc7 ) begin
                    I5046227e18f800785f8ddfb4a89b1bea  <= Ia66176893fe306ecfb415d948c50486d;
                    Iaee3ca649d20dd29363781e8dcae17c0  <=  0;
                end else begin
                    I5046227e18f800785f8ddfb4a89b1bea  <=  ~Ia66176893fe306ecfb415d948c50486d + 1;
                    Iaee3ca649d20dd29363781e8dcae17c0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iad642c4c62766e8f8bd5a1e9e73bdc80 == Ia13212b613a21e983b097fe0adbe59ec ) begin
                    I73feb8438775bf3faffed6895b6a4638  <= I8bd4210dcbfc1956381b460fd9ef789b;
                    Id8bb7c6409e383793af592892caf23e4  <=  0;
                end else begin
                    I73feb8438775bf3faffed6895b6a4638  <=  ~I8bd4210dcbfc1956381b460fd9ef789b + 1;
                    Id8bb7c6409e383793af592892caf23e4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96f92481be1ac6cf985b8ab387d326bf == Ieeddfaf876af8120f779286b4f60f767 ) begin
                    I6a423d4e11a97d84120a475db8fabca1  <= I1ba6328ea9cb7cebcce47d5407d0eae7;
                    I96c6b861bfaad7c411db93f1318d6b87  <=  0;
                end else begin
                    I6a423d4e11a97d84120a475db8fabca1  <=  ~I1ba6328ea9cb7cebcce47d5407d0eae7 + 1;
                    I96c6b861bfaad7c411db93f1318d6b87  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96f92481be1ac6cf985b8ab387d326bf == If1912201b852f91e8aa0c73439ca7022 ) begin
                    I2098616787bd728bc4af6be5ee094bae  <= I9e79c17bd782bb7981b4a3623baf96a1;
                    I76eb400ed4d1502f7f1864d9556948ad  <=  0;
                end else begin
                    I2098616787bd728bc4af6be5ee094bae  <=  ~I9e79c17bd782bb7981b4a3623baf96a1 + 1;
                    I76eb400ed4d1502f7f1864d9556948ad  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96f92481be1ac6cf985b8ab387d326bf == I0995a527d1b13090cf68b771d591c041 ) begin
                    Id9ef21a12edf48e574256ea34fcde992  <= I7c6f64d73ff9c6e7f2ed69713e056a2b;
                    I02155a5c26345ff00d18cec6e2f01592  <=  0;
                end else begin
                    Id9ef21a12edf48e574256ea34fcde992  <=  ~I7c6f64d73ff9c6e7f2ed69713e056a2b + 1;
                    I02155a5c26345ff00d18cec6e2f01592  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I96f92481be1ac6cf985b8ab387d326bf == I04bb94f5e9927cb7efa70e68658862d3 ) begin
                    I31ab57596896201ff52990b0641b9511  <= I00b962a9bf04b62244591051d2dfdbbd;
                    I91e6dcd9fa2efd055125878ab38de3fd  <=  0;
                end else begin
                    I31ab57596896201ff52990b0641b9511  <=  ~I00b962a9bf04b62244591051d2dfdbbd + 1;
                    I91e6dcd9fa2efd055125878ab38de3fd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie03c09039ccafb427153d2347c1caea8 == I7594f22f889c391838f987765ad478e7 ) begin
                    Ib3dd33a163b0c8153edb4fcc90a453f2  <= I3a660b57588325989319701026f658e6;
                    If561e078b234a0be8c0b8ade8f5ec0f1  <=  0;
                end else begin
                    Ib3dd33a163b0c8153edb4fcc90a453f2  <=  ~I3a660b57588325989319701026f658e6 + 1;
                    If561e078b234a0be8c0b8ade8f5ec0f1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie03c09039ccafb427153d2347c1caea8 == I93a25759f720769b941088884bb6db59 ) begin
                    I28496a34b2ee033767fd64f631426b23  <= Ibae27cccf3f64e8653c1e244e940e421;
                    I0ef01533d6494ce8f092d54c5fb0865e  <=  0;
                end else begin
                    I28496a34b2ee033767fd64f631426b23  <=  ~Ibae27cccf3f64e8653c1e244e940e421 + 1;
                    I0ef01533d6494ce8f092d54c5fb0865e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie03c09039ccafb427153d2347c1caea8 == Id518694e3b3a268e7168c17250bfab52 ) begin
                    I0a4ef7fac369df46d1a4b094d7687645  <= I27b89a5001312b2aa48fe385d8a52063;
                    I782b73148fd7ed7f9d734baf42b8b5d0  <=  0;
                end else begin
                    I0a4ef7fac369df46d1a4b094d7687645  <=  ~I27b89a5001312b2aa48fe385d8a52063 + 1;
                    I782b73148fd7ed7f9d734baf42b8b5d0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie03c09039ccafb427153d2347c1caea8 == Ieaf2b41941b840b3ade630e721e6367a ) begin
                    Ie7944f3e2adfac325808f8711c0eedcd  <= Ic6a7476db711a812d146331c562ca7c9;
                    I2099d6f614a5f7432f6331b1bf56c31c  <=  0;
                end else begin
                    Ie7944f3e2adfac325808f8711c0eedcd  <=  ~Ic6a7476db711a812d146331c562ca7c9 + 1;
                    I2099d6f614a5f7432f6331b1bf56c31c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie7381a8294b4cdf669b9c57cfe4012b5 == I01a2be56c727d7ca0c5059e8d34919cb ) begin
                    I58cecb5376f675339028440f0671b0b7  <= I01ca07fe91b5f1edf87300b3583e77c5;
                    Ia8c9228b5d23c91ac06450ab1296dc65  <=  0;
                end else begin
                    I58cecb5376f675339028440f0671b0b7  <=  ~I01ca07fe91b5f1edf87300b3583e77c5 + 1;
                    Ia8c9228b5d23c91ac06450ab1296dc65  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie7381a8294b4cdf669b9c57cfe4012b5 == I605682c90ff448b91a2e1a82a3cb0c08 ) begin
                    I62f85c1602819e586d9656ba42d263c3  <= I6da707fd74249175d1f68dccb66390c0;
                    I4b76ea8b5d4ed8ccd8ec532889dd6d4b  <=  0;
                end else begin
                    I62f85c1602819e586d9656ba42d263c3  <=  ~I6da707fd74249175d1f68dccb66390c0 + 1;
                    I4b76ea8b5d4ed8ccd8ec532889dd6d4b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie7381a8294b4cdf669b9c57cfe4012b5 == I0a075b833950927c58d8f55264947f00 ) begin
                    I79585885950084095d2ce4a31aa73e4c  <= I0ae62aae426b75b06d95c46baf33f08e;
                    Ifff6d20dcf891c78ad12a304ca757c95  <=  0;
                end else begin
                    I79585885950084095d2ce4a31aa73e4c  <=  ~I0ae62aae426b75b06d95c46baf33f08e + 1;
                    Ifff6d20dcf891c78ad12a304ca757c95  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie7381a8294b4cdf669b9c57cfe4012b5 == I3b699342f0100a2d56c7013da055fdd6 ) begin
                    Ic3af09106eada35f1d786ed60e314ea5  <= Iec512b5870f295a50921e7e0289a7d35;
                    I0dbefebca7ff055a6e9dce2a2c37bd69  <=  0;
                end else begin
                    Ic3af09106eada35f1d786ed60e314ea5  <=  ~Iec512b5870f295a50921e7e0289a7d35 + 1;
                    I0dbefebca7ff055a6e9dce2a2c37bd69  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61c9e3f8e42f869f4c9c1386325100b3 == Ic223e47525ca27261b7db8c1afddadc9 ) begin
                    I81e374d671edb31d060875cdfdcd61c7  <= I3aac84acd9d78070472b1cbc745c80a7;
                    I8aadd755861e90ac12047f259091ad85  <=  0;
                end else begin
                    I81e374d671edb31d060875cdfdcd61c7  <=  ~I3aac84acd9d78070472b1cbc745c80a7 + 1;
                    I8aadd755861e90ac12047f259091ad85  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61c9e3f8e42f869f4c9c1386325100b3 == Ibb5c74ed3a37c5e244e537e8b8d403fb ) begin
                    I1e22ea5ecaf87499b7106246a824a547  <= Ibbb900f56de318bf6e65b49791835ef4;
                    Ia7d21a17d62e7bfb00b83b244201e941  <=  0;
                end else begin
                    I1e22ea5ecaf87499b7106246a824a547  <=  ~Ibbb900f56de318bf6e65b49791835ef4 + 1;
                    Ia7d21a17d62e7bfb00b83b244201e941  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61c9e3f8e42f869f4c9c1386325100b3 == I5915ba867f798193c35a4af58e8cabf6 ) begin
                    I0e46eb0f32c91384b07c7b1ba84caf98  <= I2c2ac1e722fba72c759f1d37b88a9a10;
                    I6c63fab8059cc3f0c02b0dff5a8cacf9  <=  0;
                end else begin
                    I0e46eb0f32c91384b07c7b1ba84caf98  <=  ~I2c2ac1e722fba72c759f1d37b88a9a10 + 1;
                    I6c63fab8059cc3f0c02b0dff5a8cacf9  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I61c9e3f8e42f869f4c9c1386325100b3 == I73ce6acb5ca8a57906440578f4ae15aa ) begin
                    I562b5f77aedd91f0cb3df00387c7956a  <= Ida0a18f1b79aff4ddf0e8f7e27794674;
                    I8744fea2c7de33b5308dc9a2828647d4  <=  0;
                end else begin
                    I562b5f77aedd91f0cb3df00387c7956a  <=  ~Ida0a18f1b79aff4ddf0e8f7e27794674 + 1;
                    I8744fea2c7de33b5308dc9a2828647d4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24c5b2de59eb1f43fe1efe687231c4b7 == I9cea4e30593a1275f4450adb25b5c5cb ) begin
                    Id819e47f502c18dca8d1e804d346c1ea  <= I9f2029db42c5a968b370587c958c8929;
                    I04c99b4d0c54b23a72b698753510a4f3  <=  0;
                end else begin
                    Id819e47f502c18dca8d1e804d346c1ea  <=  ~I9f2029db42c5a968b370587c958c8929 + 1;
                    I04c99b4d0c54b23a72b698753510a4f3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24c5b2de59eb1f43fe1efe687231c4b7 == I3dacee8649adfc1a8b2092f5af3cada6 ) begin
                    Ie0586f4b015fd32777d24c2d9856b27f  <= If5755f4f61a89d91a91188c17ff5dc5a;
                    I5de86a27849e73b21e4c40e9e8515033  <=  0;
                end else begin
                    Ie0586f4b015fd32777d24c2d9856b27f  <=  ~If5755f4f61a89d91a91188c17ff5dc5a + 1;
                    I5de86a27849e73b21e4c40e9e8515033  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24c5b2de59eb1f43fe1efe687231c4b7 == I00537a49036c970d6df97b3917de104e ) begin
                    Ic28248b41552d2537d0478c23e33e0f3  <= I4419d97c3174ee4610eb6ee9c06cb256;
                    I185257f76b2886cd845e50a01ef5b05b  <=  0;
                end else begin
                    Ic28248b41552d2537d0478c23e33e0f3  <=  ~I4419d97c3174ee4610eb6ee9c06cb256 + 1;
                    I185257f76b2886cd845e50a01ef5b05b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I43d43acde5f831fc32b7bf5f10b9b3a9 == If6ce1f97c23f1d1bf23c283ce37682ce ) begin
                    I3463cbe0d16b14aa670fda6a0d34e255  <= Ia964f83676273055e20a2f63c8fffa0d;
                    I1a2c7b5505f4124f945a28565eed6013  <=  0;
                end else begin
                    I3463cbe0d16b14aa670fda6a0d34e255  <=  ~Ia964f83676273055e20a2f63c8fffa0d + 1;
                    I1a2c7b5505f4124f945a28565eed6013  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I43d43acde5f831fc32b7bf5f10b9b3a9 == Ieae92b67815d507df906e1be71d6346b ) begin
                    I0aac7a09d9253385d34e87bfbb216a79  <= Iab4fbc811e87df1d1f5821ea732b6a93;
                    I771d417f6226b04ef016d0943bbc4584  <=  0;
                end else begin
                    I0aac7a09d9253385d34e87bfbb216a79  <=  ~Iab4fbc811e87df1d1f5821ea732b6a93 + 1;
                    I771d417f6226b04ef016d0943bbc4584  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I43d43acde5f831fc32b7bf5f10b9b3a9 == I1af89e1ec1210d4d3dafc0927b62afe5 ) begin
                    I305967a657db8531d1ae309fa3e3b98f  <= I4fbefbb10724b0844c95e85495d4a87f;
                    Icb0a73f2dd46e2195d5efd34fba3a985  <=  0;
                end else begin
                    I305967a657db8531d1ae309fa3e3b98f  <=  ~I4fbefbb10724b0844c95e85495d4a87f + 1;
                    Icb0a73f2dd46e2195d5efd34fba3a985  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib06e93161fc8ca3be232f4261b04feb1 == Ic264e7826b90e379048b094875eeb921 ) begin
                    I0524108ee49eec5fa7861bed35e4ea3c  <= I717217d0b5a526f04c7f5ab0835dd5c7;
                    Ia992f7eacefc028526ab4f105e244e02  <=  0;
                end else begin
                    I0524108ee49eec5fa7861bed35e4ea3c  <=  ~I717217d0b5a526f04c7f5ab0835dd5c7 + 1;
                    Ia992f7eacefc028526ab4f105e244e02  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib06e93161fc8ca3be232f4261b04feb1 == Iea6d4bb1137e579b1605a16c578cbd7d ) begin
                    Iced1e0b874918a1c66e28752e340a51b  <= I235937b643e8f2848116dc76c43f47a7;
                    I85454620b6568bb7fde468a2e9a5fb42  <=  0;
                end else begin
                    Iced1e0b874918a1c66e28752e340a51b  <=  ~I235937b643e8f2848116dc76c43f47a7 + 1;
                    I85454620b6568bb7fde468a2e9a5fb42  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib06e93161fc8ca3be232f4261b04feb1 == I706d85c9d83bcfc5a2204a67e5c1f84e ) begin
                    I670e910f74fafccaa9f1a8279fd6ebb6  <= I7481f17d659cce5b4c72a68a9f6be67f;
                    I87557ef641a7b209d4d210498bb15271  <=  0;
                end else begin
                    I670e910f74fafccaa9f1a8279fd6ebb6  <=  ~I7481f17d659cce5b4c72a68a9f6be67f + 1;
                    I87557ef641a7b209d4d210498bb15271  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia0dd00f83afc805036f2c6a0e38f725e == I6e832b004d0dddf4c3edb682669acf7a ) begin
                    I02fe6b32b2405fb94afd5d7abbaf0195  <= I5715c21c80992a61bff8aabc3f80415b;
                    I28d1125b647b953f2a19ecd6edd8e450  <=  0;
                end else begin
                    I02fe6b32b2405fb94afd5d7abbaf0195  <=  ~I5715c21c80992a61bff8aabc3f80415b + 1;
                    I28d1125b647b953f2a19ecd6edd8e450  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia0dd00f83afc805036f2c6a0e38f725e == Id0f69c70b38b7483a19e32d5982bb4b5 ) begin
                    I5f5304e4b132f816c87248d3ca954164  <= I434e3216a615eb46be5c26ef914b9cd2;
                    I4a8aa3010248f0bdd3e31822bf2fe0a1  <=  0;
                end else begin
                    I5f5304e4b132f816c87248d3ca954164  <=  ~I434e3216a615eb46be5c26ef914b9cd2 + 1;
                    I4a8aa3010248f0bdd3e31822bf2fe0a1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia0dd00f83afc805036f2c6a0e38f725e == I9cb245dceba82553db23cb15854f59f1 ) begin
                    I0ecebe47e1a9ede33c3995945a6ee760  <= I918326ac0a744d234d74e2c08cf41eb4;
                    Ie1966fd5b564dd6eccfc458e9c6aca2a  <=  0;
                end else begin
                    I0ecebe47e1a9ede33c3995945a6ee760  <=  ~I918326ac0a744d234d74e2c08cf41eb4 + 1;
                    Ie1966fd5b564dd6eccfc458e9c6aca2a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 == I978d0157f7403d2f35fa648271f4fbd9 ) begin
                    If425109071b5310e097d2174625b6383  <= I966706d314f4c0a7ec842dd699d34926;
                    I8ad51753f106d0a30cc79bd08e799348  <=  0;
                end else begin
                    If425109071b5310e097d2174625b6383  <=  ~I966706d314f4c0a7ec842dd699d34926 + 1;
                    I8ad51753f106d0a30cc79bd08e799348  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 == I70e5f31e8c4f1aa9a9aa21c28ba20d08 ) begin
                    Ic0f324c7ba05a7cfae9d70b62e30f94b  <= I5a7d246d88ef12e999f4bdee40e5a585;
                    I1c3bf915a6b62d22d04b8c8d92a72a73  <=  0;
                end else begin
                    Ic0f324c7ba05a7cfae9d70b62e30f94b  <=  ~I5a7d246d88ef12e999f4bdee40e5a585 + 1;
                    I1c3bf915a6b62d22d04b8c8d92a72a73  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 == I3cf2040a93a0184f619ce941c4f910d0 ) begin
                    I35631cbe926290974c90ddeb9b07f231  <= Ic2dfaf65c4e17a8dcd55f766c314d6ef;
                    Ie557629e9d52e5fa7435b4fb19e5276f  <=  0;
                end else begin
                    I35631cbe926290974c90ddeb9b07f231  <=  ~Ic2dfaf65c4e17a8dcd55f766c314d6ef + 1;
                    Ie557629e9d52e5fa7435b4fb19e5276f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 == I3278841178f87a4d0ccdf8316c3fb689 ) begin
                    Iceae425f37f3b1194a2ef5cd46d1b6eb  <= I151831ba6bd0e162275c84815e3c0f12;
                    I38fc977bb1d52cbc5e02a6733f6a8190  <=  0;
                end else begin
                    Iceae425f37f3b1194a2ef5cd46d1b6eb  <=  ~I151831ba6bd0e162275c84815e3c0f12 + 1;
                    I38fc977bb1d52cbc5e02a6733f6a8190  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib0a0f924fe3757a1e0aade7017ad9277 == I73d0e5f3635c5a2c3f1824c578c07658 ) begin
                    I4faa2187d970078870078c3eff180b4a  <= I5a8f1675234ebed14d719344b530bbd7;
                    If84914aaabb020baad2b222f27c9ad38  <=  0;
                end else begin
                    I4faa2187d970078870078c3eff180b4a  <=  ~I5a8f1675234ebed14d719344b530bbd7 + 1;
                    If84914aaabb020baad2b222f27c9ad38  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1ca949071d734d230cdb8adda46c9d79 == Id1b7ef639fcb74c8fa47fd7ef0cbe96c ) begin
                    Iec2860f518edf688a9b1b2736ae00835  <= I95dce76a8d0e729d40fb3f573cfc06ad;
                    I54c457a658721fa7de175432b340532e  <=  0;
                end else begin
                    Iec2860f518edf688a9b1b2736ae00835  <=  ~I95dce76a8d0e729d40fb3f573cfc06ad + 1;
                    I54c457a658721fa7de175432b340532e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1ca949071d734d230cdb8adda46c9d79 == I1c83edeea3cd4c32bae64594a2f8b256 ) begin
                    I20e7b48527e4456874d59e50c723c6a5  <= I6c26c7918254426c18f2e747c91438c5;
                    I9036f6cf74a2aecd827c7239da13db70  <=  0;
                end else begin
                    I20e7b48527e4456874d59e50c723c6a5  <=  ~I6c26c7918254426c18f2e747c91438c5 + 1;
                    I9036f6cf74a2aecd827c7239da13db70  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1ca949071d734d230cdb8adda46c9d79 == I0b930276a1887380da03c22aa8fb9adb ) begin
                    Idd60af0dbb02680e11c1b1734f23b895  <= I0414ead2472e42da8a271cb0bd1debf4;
                    I8825e2665dcee58925a5106a9cbce9ca  <=  0;
                end else begin
                    Idd60af0dbb02680e11c1b1734f23b895  <=  ~I0414ead2472e42da8a271cb0bd1debf4 + 1;
                    I8825e2665dcee58925a5106a9cbce9ca  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1ca949071d734d230cdb8adda46c9d79 == I63ec886123f0ff76bfa46c2d6b2c5760 ) begin
                    I79cfbb5d5e920bc8cece60565ee0c5c2  <= Ic6a6f5090470a76ddb7315c022ddc104;
                    Ic3311c2f88a7ae151999b2de86d82dfc  <=  0;
                end else begin
                    I79cfbb5d5e920bc8cece60565ee0c5c2  <=  ~Ic6a6f5090470a76ddb7315c022ddc104 + 1;
                    Ic3311c2f88a7ae151999b2de86d82dfc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I1ca949071d734d230cdb8adda46c9d79 == I32bf44d4f4df42cb664e75ccef06fb34 ) begin
                    Id765a3f659dcdf01cfe23cafdf066f92  <= I2a00ee56a5aa639f45eb3b1bdcffe81c;
                    I3ef7eddb92284b28f97feea52f489aff  <=  0;
                end else begin
                    Id765a3f659dcdf01cfe23cafdf066f92  <=  ~I2a00ee56a5aa639f45eb3b1bdcffe81c + 1;
                    I3ef7eddb92284b28f97feea52f489aff  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40170922c652fa7fa42abc6f580b5e3d == Iadc0319541fc978cd0efbdf5b3af7078 ) begin
                    If370aaa56b4ba3eee873c99a86577c3d  <= Ibceb2b824cd4bc10bb06ee8adc693bd1;
                    I68728d0cbb3a84370006277186a0829d  <=  0;
                end else begin
                    If370aaa56b4ba3eee873c99a86577c3d  <=  ~Ibceb2b824cd4bc10bb06ee8adc693bd1 + 1;
                    I68728d0cbb3a84370006277186a0829d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40170922c652fa7fa42abc6f580b5e3d == I9f4036502b40315cfa7d8bb9b83b5806 ) begin
                    I4508376202467dc1bebc69757bd5f95a  <= Ia8b9f373fe68ac4cbca35e04376e3cca;
                    If5bdbdfa73406a6a9d426920f51fbc73  <=  0;
                end else begin
                    I4508376202467dc1bebc69757bd5f95a  <=  ~Ia8b9f373fe68ac4cbca35e04376e3cca + 1;
                    If5bdbdfa73406a6a9d426920f51fbc73  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40170922c652fa7fa42abc6f580b5e3d == I91dd649eab4a8eb0f8d97553560d3b7e ) begin
                    Ibf115f80ad72df8599073c05ac58e028  <= I5d1a89e85f6609b469e73e15aeffcbc4;
                    Ibd3179c01665a17f9c232196648de8d5  <=  0;
                end else begin
                    Ibf115f80ad72df8599073c05ac58e028  <=  ~I5d1a89e85f6609b469e73e15aeffcbc4 + 1;
                    Ibd3179c01665a17f9c232196648de8d5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40170922c652fa7fa42abc6f580b5e3d == Iee09e9c54961c380ff7e1758c84d663e ) begin
                    I27960a9d3923d053d466955c660a91ca  <= I677fe06bad241bc8dd6a65a97f6db520;
                    I42c2c03a158ed79ea91ea6b9f9a6f243  <=  0;
                end else begin
                    I27960a9d3923d053d466955c660a91ca  <=  ~I677fe06bad241bc8dd6a65a97f6db520 + 1;
                    I42c2c03a158ed79ea91ea6b9f9a6f243  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I40170922c652fa7fa42abc6f580b5e3d == Iaec27722c40c7cb0c0baaee4d30adc72 ) begin
                    I7c52711e3b71823dd47861341d22adc3  <= If3c0f892fd71eb0ed8d1f70b4b33450b;
                    Iec064c18b262b95bd6412b1e50e4b5ef  <=  0;
                end else begin
                    I7c52711e3b71823dd47861341d22adc3  <=  ~If3c0f892fd71eb0ed8d1f70b4b33450b + 1;
                    Iec064c18b262b95bd6412b1e50e4b5ef  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 == I5fe79d8695d426ba54609af4b38bf2dd ) begin
                    I547ea6a130740e4b0bb85f6c9d3a6549  <= Ic65f0f75f56bf85122a89cdf07e98152;
                    I0470f0fd133851c1241c654abc19992a  <=  0;
                end else begin
                    I547ea6a130740e4b0bb85f6c9d3a6549  <=  ~Ic65f0f75f56bf85122a89cdf07e98152 + 1;
                    I0470f0fd133851c1241c654abc19992a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 == I8a2b1e09c6f852b0aa4e599e7ef42187 ) begin
                    I0ec19c18ef7da4793427a00a652a9a35  <= I41d22bafaf58e4a6de04640864653a16;
                    I550661edfa7a7b440d43c0840aeed8fe  <=  0;
                end else begin
                    I0ec19c18ef7da4793427a00a652a9a35  <=  ~I41d22bafaf58e4a6de04640864653a16 + 1;
                    I550661edfa7a7b440d43c0840aeed8fe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 == Ie1f415cbb2d3e1d46f2e0e4201fe7ba0 ) begin
                    I640d147f241267ccc89f9ab132d724f8  <= I06a46b86f6edede0f5f72658a19910b7;
                    I2f01145e1b41f2f7103c5247bb548a6b  <=  0;
                end else begin
                    I640d147f241267ccc89f9ab132d724f8  <=  ~I06a46b86f6edede0f5f72658a19910b7 + 1;
                    I2f01145e1b41f2f7103c5247bb548a6b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 == I46a75678565a43e0da6b6dc55686c4c8 ) begin
                    I3507152877484394769c12879ce0aed0  <= I8591d0399594adacfeb006c5195c2c71;
                    I34d143e9a6f936b83863a5ebdf8afc43  <=  0;
                end else begin
                    I3507152877484394769c12879ce0aed0  <=  ~I8591d0399594adacfeb006c5195c2c71 + 1;
                    I34d143e9a6f936b83863a5ebdf8afc43  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib1ad0b531ac9028971d68f533e7ae566 == I200bec7d713bc7f05dc3931f20523763 ) begin
                    I382f86490f568ead2dcf51e8bc6989f8  <= Id90588b5f82cd32e801fbea04d24e4a5;
                    Id2f831bc219ca3f43c5c4d69f6724e64  <=  0;
                end else begin
                    I382f86490f568ead2dcf51e8bc6989f8  <=  ~Id90588b5f82cd32e801fbea04d24e4a5 + 1;
                    Id2f831bc219ca3f43c5c4d69f6724e64  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0ab0170c7ceffbb58377b65d2ad92093 == I978b7018cd38c7c4f0b6199cc46d258c ) begin
                    I953178c54a672474dda2f48c70ec21a7  <= Ib642d757fae818cd6d713ffb6ce18fc1;
                    Ib708fd61ab7016190a2a7156439201cf  <=  0;
                end else begin
                    I953178c54a672474dda2f48c70ec21a7  <=  ~Ib642d757fae818cd6d713ffb6ce18fc1 + 1;
                    Ib708fd61ab7016190a2a7156439201cf  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0ab0170c7ceffbb58377b65d2ad92093 == I9d298dcd244445c8a047a1ac056fb6a6 ) begin
                    I13b43982093e885ae7bb04a2b61e4eaa  <= Id76bff2a12cf792e52ccc463647334c0;
                    I6a2e574a2d27e40faff379b6c26ae51b  <=  0;
                end else begin
                    I13b43982093e885ae7bb04a2b61e4eaa  <=  ~Id76bff2a12cf792e52ccc463647334c0 + 1;
                    I6a2e574a2d27e40faff379b6c26ae51b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I0ab0170c7ceffbb58377b65d2ad92093 == Ib5de0226d215418202f2cff36b573daa ) begin
                    I3d7491ac28a4adafbc138d17f08c9111  <= I92ffa890ed6d83d4fc543504e4d421c1;
                    I4be2286baca2745e981a0d153c0f5c42  <=  0;
                end else begin
                    I3d7491ac28a4adafbc138d17f08c9111  <=  ~I92ffa890ed6d83d4fc543504e4d421c1 + 1;
                    I4be2286baca2745e981a0d153c0f5c42  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ac68f228a93bbf4aa4a559b1364e42e == I58e42ededb36d8aaf022e7b42a8fb36c ) begin
                    I3e0ca15752add87cc01981e7d89d53f2  <= Ifc4a65edeaf630b3d29437bcd6c20121;
                    Ib9643265dc8c283d7b0c7afdb19101fd  <=  0;
                end else begin
                    I3e0ca15752add87cc01981e7d89d53f2  <=  ~Ifc4a65edeaf630b3d29437bcd6c20121 + 1;
                    Ib9643265dc8c283d7b0c7afdb19101fd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ac68f228a93bbf4aa4a559b1364e42e == I8017904689642a7e3d82c34839403614 ) begin
                    Id1b152deea3ee894ed5a4c6ff10a6fda  <= Id57a11f56fc223501a9b68b8b05ebd3e;
                    I78d7637bbd13c620434d3619e615114c  <=  0;
                end else begin
                    Id1b152deea3ee894ed5a4c6ff10a6fda  <=  ~Id57a11f56fc223501a9b68b8b05ebd3e + 1;
                    I78d7637bbd13c620434d3619e615114c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ac68f228a93bbf4aa4a559b1364e42e == I773d6a848aa20abe6d1ebf8f7d6dad85 ) begin
                    I7df9cc0e3ad69985fe9a3c8f2dec1de3  <= I522ba8bfc1949337e8befe82cc1e86e6;
                    I358ee555d9955cdee436375ff898f4d6  <=  0;
                end else begin
                    I7df9cc0e3ad69985fe9a3c8f2dec1de3  <=  ~I522ba8bfc1949337e8befe82cc1e86e6 + 1;
                    I358ee555d9955cdee436375ff898f4d6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I375c5f7eac92d853e85e0606011f3fb0 == I8bafb2d0a6bf186c179ee07ed51a2e33 ) begin
                    I52910c0c2d26095c965d32b85e850d92  <= I7153e27c44ebbc2f04e9ba03cf09b5e1;
                    Ic3961c918c81b14d964e96892b95f00b  <=  0;
                end else begin
                    I52910c0c2d26095c965d32b85e850d92  <=  ~I7153e27c44ebbc2f04e9ba03cf09b5e1 + 1;
                    Ic3961c918c81b14d964e96892b95f00b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I375c5f7eac92d853e85e0606011f3fb0 == I63d8a99e826b0d6a5051fb454f15f44a ) begin
                    I93fd4b4f7d01ec59834f3054fc2eddfd  <= Id15e4b4f186ec863f12a54acd8ef8963;
                    I580e98d4bec3eeeb1642baa425a96099  <=  0;
                end else begin
                    I93fd4b4f7d01ec59834f3054fc2eddfd  <=  ~Id15e4b4f186ec863f12a54acd8ef8963 + 1;
                    I580e98d4bec3eeeb1642baa425a96099  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I375c5f7eac92d853e85e0606011f3fb0 == I0b831c8e1d7187024eb93f980cb04f61 ) begin
                    I481b6feb1f1ced501a157b06a4782e05  <= I95c77eec7575cd7aa93a36f31ea635a2;
                    I4cec0a54301908b3f58166a9b0ef1eb5  <=  0;
                end else begin
                    I481b6feb1f1ced501a157b06a4782e05  <=  ~I95c77eec7575cd7aa93a36f31ea635a2 + 1;
                    I4cec0a54301908b3f58166a9b0ef1eb5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I94f9b1f2e63748c21ec7222c9641366a == I17867f12563819dd7b89f9079fb0a385 ) begin
                    Ie99b8f3190ee307e743255156b7f7f90  <= I3c8114dbe0658cc2889c787f1366abfa;
                    Ib7f7c88d83d207bac3daba4658342879  <=  0;
                end else begin
                    Ie99b8f3190ee307e743255156b7f7f90  <=  ~I3c8114dbe0658cc2889c787f1366abfa + 1;
                    Ib7f7c88d83d207bac3daba4658342879  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I94f9b1f2e63748c21ec7222c9641366a == I2a2b4eaef143deb9e61110334dc5c2ea ) begin
                    Iac858597facbc0025a4760eac49531fe  <= Ieacf971e9e10fb73c7df9f1da8372f30;
                    I371401ca0c589a1b8fa816beed36ab0c  <=  0;
                end else begin
                    Iac858597facbc0025a4760eac49531fe  <=  ~Ieacf971e9e10fb73c7df9f1da8372f30 + 1;
                    I371401ca0c589a1b8fa816beed36ab0c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I94f9b1f2e63748c21ec7222c9641366a == Ieb02d465c1ac76962dd663067ebcd445 ) begin
                    I18c2833554a5b358578e7b6901c91c0c  <= I35de1b03ea865f2c6381ce73e03dc220;
                    I81f561f223b916600ebc572c05dedde5  <=  0;
                end else begin
                    I18c2833554a5b358578e7b6901c91c0c  <=  ~I35de1b03ea865f2c6381ce73e03dc220 + 1;
                    I81f561f223b916600ebc572c05dedde5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I55500c1d85c4970932be67cc5cd2e023 == I6ad4bc4bc7c0f005307199814893faee ) begin
                    I0cc6945a47b3ffadd1e52e3f71c9728d  <= Idec12e02904ea98c7580919584f2dba1;
                    I7ee36d73f8c69e5e017f4616094d992f  <=  0;
                end else begin
                    I0cc6945a47b3ffadd1e52e3f71c9728d  <=  ~Idec12e02904ea98c7580919584f2dba1 + 1;
                    I7ee36d73f8c69e5e017f4616094d992f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I55500c1d85c4970932be67cc5cd2e023 == If9a814db74759469b79411ed7038c860 ) begin
                    If2807866c5d481cd31c69b67ec537a4f  <= Ia370c83631a2c1bbf39c7264deafafb5;
                    I706d7d2238c5882491d479df0cc40c3e  <=  0;
                end else begin
                    If2807866c5d481cd31c69b67ec537a4f  <=  ~Ia370c83631a2c1bbf39c7264deafafb5 + 1;
                    I706d7d2238c5882491d479df0cc40c3e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I55500c1d85c4970932be67cc5cd2e023 == I3d0f05a6136e0c14536830bc53a5333d ) begin
                    Ib24d495a86e15d9c8b2c8d360445e511  <= I05b4a07dfc0d2695eae34bea4c1c6565;
                    Ie28bec241cb36d75c1f2ad846dc5c7d6  <=  0;
                end else begin
                    Ib24d495a86e15d9c8b2c8d360445e511  <=  ~I05b4a07dfc0d2695eae34bea4c1c6565 + 1;
                    Ie28bec241cb36d75c1f2ad846dc5c7d6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I55500c1d85c4970932be67cc5cd2e023 == I1f168715063587b7dfb01e0fefbca615 ) begin
                    Iad2cdac80bc26a0c50335c6467921c94  <= If1ecdc27e3419dd1434e403f237c2b58;
                    I9fe8aa4f9f74c1f004e5bb536e902ea2  <=  0;
                end else begin
                    Iad2cdac80bc26a0c50335c6467921c94  <=  ~If1ecdc27e3419dd1434e403f237c2b58 + 1;
                    I9fe8aa4f9f74c1f004e5bb536e902ea2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I36b487cd1a57a3a503e587fdefbb19e4 == Ida3cc6922fe4edded7f2e59b909d6d72 ) begin
                    I18c93f107d0520171864b789ae9707b9  <= I039c552777d0fb40bebcdd2d4a3394c2;
                    I444003b27464f275311d07ae7d4fe016  <=  0;
                end else begin
                    I18c93f107d0520171864b789ae9707b9  <=  ~I039c552777d0fb40bebcdd2d4a3394c2 + 1;
                    I444003b27464f275311d07ae7d4fe016  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I36b487cd1a57a3a503e587fdefbb19e4 == Ic2b81c5409d555402164dd12ae7decc4 ) begin
                    Ifd40aae90a89d2420e43fe4ee533a1a2  <= Iaa52fb63184514b6d754bcc896235150;
                    Ibbe636e1e98bbd4cd97dca56d769d269  <=  0;
                end else begin
                    Ifd40aae90a89d2420e43fe4ee533a1a2  <=  ~Iaa52fb63184514b6d754bcc896235150 + 1;
                    Ibbe636e1e98bbd4cd97dca56d769d269  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I36b487cd1a57a3a503e587fdefbb19e4 == I8edabaa27753c6f70325108c9c1b12b6 ) begin
                    If46a176f32240b03ae959e9ad889fc2c  <= Ied9781e625c1fa8741853dd6b8b3a9e7;
                    Ib195ccbfb4411bd3aaece336a5aed65b  <=  0;
                end else begin
                    If46a176f32240b03ae959e9ad889fc2c  <=  ~Ied9781e625c1fa8741853dd6b8b3a9e7 + 1;
                    Ib195ccbfb4411bd3aaece336a5aed65b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I36b487cd1a57a3a503e587fdefbb19e4 == Ie58289ff961fc431fbf10f78fda337ab ) begin
                    I5e7b386298be05835cd24554966cdedc  <= I767272262e9d2e85dba1aa93f578f25c;
                    Ieafb75c62922cdb3acd95a9614a86efc  <=  0;
                end else begin
                    I5e7b386298be05835cd24554966cdedc  <=  ~I767272262e9d2e85dba1aa93f578f25c + 1;
                    Ieafb75c62922cdb3acd95a9614a86efc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icb5350e8c55a2adb370078a7575e28f8 == I3ee219716889ea93423603105de22c6c ) begin
                    I5258d2bd4ae07dcfe7e022b046800856  <= Ib3b4cd6d8ab17869a2278552c02635c8;
                    I5d7018ab259e054ecb48a238f3c03208  <=  0;
                end else begin
                    I5258d2bd4ae07dcfe7e022b046800856  <=  ~Ib3b4cd6d8ab17869a2278552c02635c8 + 1;
                    I5d7018ab259e054ecb48a238f3c03208  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icb5350e8c55a2adb370078a7575e28f8 == I957518cfe822b5afcc1f7153e07e26c4 ) begin
                    I14da6601ba08fd3e9a2bcdd20bb43536  <= Ie7a5cb2ecb3fce35825785b9bca6b3bd;
                    Iedabb09ffcf910c4dbed2f142dc96df0  <=  0;
                end else begin
                    I14da6601ba08fd3e9a2bcdd20bb43536  <=  ~Ie7a5cb2ecb3fce35825785b9bca6b3bd + 1;
                    Iedabb09ffcf910c4dbed2f142dc96df0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icb5350e8c55a2adb370078a7575e28f8 == Id8fb66bc4afa4f7f7f4ca0d7ce3f5543 ) begin
                    I76bbfed1a115c2f503531682cd171185  <= Ib9a0f8efd3dad427f247ce90fdfb94a4;
                    I07b84cae4f002659d68f5c1746416e70  <=  0;
                end else begin
                    I76bbfed1a115c2f503531682cd171185  <=  ~Ib9a0f8efd3dad427f247ce90fdfb94a4 + 1;
                    I07b84cae4f002659d68f5c1746416e70  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Icb5350e8c55a2adb370078a7575e28f8 == I3beb0bdc4242c12a068f7aec11bf022a ) begin
                    I64f37f25618c6bf5b35e863e3be05a3e  <= I69a221a1bd95a588aa74b9bed0357762;
                    Iba31516a82e9d2a5ad1a1c89dfb6af70  <=  0;
                end else begin
                    I64f37f25618c6bf5b35e863e3be05a3e  <=  ~I69a221a1bd95a588aa74b9bed0357762 + 1;
                    Iba31516a82e9d2a5ad1a1c89dfb6af70  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I8a7a31327c9e4cbd88ce39fea8971caf == I629a5a30684270d00605b4fc02eab693 ) begin
                    Iba3b847497a7572624a3a1f172b47d3e  <= I64f125cf2ca6a6da8a9cdae9e246c24a;
                    If5c42feaf3d586e1f2285b0f3e3a2d39  <=  0;
                end else begin
                    Iba3b847497a7572624a3a1f172b47d3e  <=  ~I64f125cf2ca6a6da8a9cdae9e246c24a + 1;
                    If5c42feaf3d586e1f2285b0f3e3a2d39  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I8a7a31327c9e4cbd88ce39fea8971caf == I32aa431be1c47b8c52c3b3f6d371f439 ) begin
                    Ic9885fd472d244d4810bc9ff0971dc65  <= Ifac9dd60dd6c543aa94b39c599f0819a;
                    I3f15f6722f339c32bf1dfa41b5b24648  <=  0;
                end else begin
                    Ic9885fd472d244d4810bc9ff0971dc65  <=  ~Ifac9dd60dd6c543aa94b39c599f0819a + 1;
                    I3f15f6722f339c32bf1dfa41b5b24648  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I8a7a31327c9e4cbd88ce39fea8971caf == I88d8124a68d50e1730a87914ed6b2a55 ) begin
                    I5753bb74c9d925b91c0173bcc320af36  <= Icf062382a1e462571569ccee75b0a3ee;
                    I74d5d4a25b6ceba088652dbad9c35bae  <=  0;
                end else begin
                    I5753bb74c9d925b91c0173bcc320af36  <=  ~Icf062382a1e462571569ccee75b0a3ee + 1;
                    I74d5d4a25b6ceba088652dbad9c35bae  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I8a7a31327c9e4cbd88ce39fea8971caf == I474bd0d0a044aae82cfb1afbd3d40f74 ) begin
                    I66cf73ce0a93f90287df52adb628716d  <= Ieed8b94295bed265961c4f52c3379914;
                    I1e3e7019425109b26d4ebc7522074e33  <=  0;
                end else begin
                    I66cf73ce0a93f90287df52adb628716d  <=  ~Ieed8b94295bed265961c4f52c3379914 + 1;
                    I1e3e7019425109b26d4ebc7522074e33  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied069655ed3775819d0bcb722d6d0488 == I2bcfe7aeef8f2b772605c9ad10a289ea ) begin
                    I84a477263ea86f2014d28e9ec928fa1b  <= I165eabcdde76821fdc308ff7a8c6d2ea;
                    I4f0d4baa740b2f9bea59f4653cc9e8fc  <=  0;
                end else begin
                    I84a477263ea86f2014d28e9ec928fa1b  <=  ~I165eabcdde76821fdc308ff7a8c6d2ea + 1;
                    I4f0d4baa740b2f9bea59f4653cc9e8fc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied069655ed3775819d0bcb722d6d0488 == Id4a7c3a22060cfcaff64e2a3980dea91 ) begin
                    Idda9e2f9a5e24406700b04e6035dafc7  <= I8b3542a6d64d6a7ebba4124bc6702f3e;
                    I2df393a2d764f120433f310797abb2c3  <=  0;
                end else begin
                    Idda9e2f9a5e24406700b04e6035dafc7  <=  ~I8b3542a6d64d6a7ebba4124bc6702f3e + 1;
                    I2df393a2d764f120433f310797abb2c3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied069655ed3775819d0bcb722d6d0488 == I6085d7398ccd685c1a60a21e4a15a606 ) begin
                    I694ec5f3a1e7cfc02c1af8369064967c  <= I7b68afec199be705d766c169f1ece981;
                    Ib9a2e4c37430ad33531f318a313d4646  <=  0;
                end else begin
                    I694ec5f3a1e7cfc02c1af8369064967c  <=  ~I7b68afec199be705d766c169f1ece981 + 1;
                    Ib9a2e4c37430ad33531f318a313d4646  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ied069655ed3775819d0bcb722d6d0488 == I203cd1948326fb3fa3dc14423bf3f992 ) begin
                    Id0c6285ee3789c104e483a5626b5827d  <= I4b6c8226ef2bc20dbd31d242bdb98b8c;
                    Ide344589b18aa0332a7114424956b65b  <=  0;
                end else begin
                    Id0c6285ee3789c104e483a5626b5827d  <=  ~I4b6c8226ef2bc20dbd31d242bdb98b8c + 1;
                    Ide344589b18aa0332a7114424956b65b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I78a5fc80d42e8db1b56cce5f4c97e325 == I67412169057453e2fb39c3b0760039c0 ) begin
                    If9bc7b1498733ed921b51cb613c2cf53  <= Ic3b4a86f22caf5b6103d52b6c9d2a991;
                    I789b8e58762f722bc0e86e17c2655965  <=  0;
                end else begin
                    If9bc7b1498733ed921b51cb613c2cf53  <=  ~Ic3b4a86f22caf5b6103d52b6c9d2a991 + 1;
                    I789b8e58762f722bc0e86e17c2655965  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I78a5fc80d42e8db1b56cce5f4c97e325 == I520d93aaf6b72a2ec7c23ae4e253aa07 ) begin
                    Ieeda4b6b301d662ab9be9f6b979bb1f1  <= Ia37592b207086f63e2d94e3d7d26c740;
                    I243898aa7700f57974ea2834df469f48  <=  0;
                end else begin
                    Ieeda4b6b301d662ab9be9f6b979bb1f1  <=  ~Ia37592b207086f63e2d94e3d7d26c740 + 1;
                    I243898aa7700f57974ea2834df469f48  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I78a5fc80d42e8db1b56cce5f4c97e325 == I34a77904a4a75d2907acd173bf27800c ) begin
                    Icad98c93196218a7dbd25af042b4a32d  <= Id0d786026e3ab0ddbffbc20e4d409857;
                    Ic65d6b89fc082438b9956504f30a5483  <=  0;
                end else begin
                    Icad98c93196218a7dbd25af042b4a32d  <=  ~Id0d786026e3ab0ddbffbc20e4d409857 + 1;
                    Ic65d6b89fc082438b9956504f30a5483  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I78a5fc80d42e8db1b56cce5f4c97e325 == I7a4ea8ffce8d52bb241553a681408dec ) begin
                    I408e198b0eeade8b94c27ab7e04a8776  <= I333837f976cfc7f90ab0a6dcd8c1ce79;
                    Ibdcf7926e0b7412e4a56d2ae15a4e892  <=  0;
                end else begin
                    I408e198b0eeade8b94c27ab7e04a8776  <=  ~I333837f976cfc7f90ab0a6dcd8c1ce79 + 1;
                    Ibdcf7926e0b7412e4a56d2ae15a4e892  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3ade7e345432319c1a9c91d4068b3ec9 == I8e89fb1ed1d604bbf0177e0c61da6e94 ) begin
                    I24b90526a93dc177a5d23b61d20f8797  <= Id115b4708a49dcfd167e79ef6993e371;
                    Ie552917ecc454608adca6dbc4d9153ad  <=  0;
                end else begin
                    I24b90526a93dc177a5d23b61d20f8797  <=  ~Id115b4708a49dcfd167e79ef6993e371 + 1;
                    Ie552917ecc454608adca6dbc4d9153ad  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3ade7e345432319c1a9c91d4068b3ec9 == I5d2148b5809cd169c41663caa441c464 ) begin
                    I4da324410e88d8c9738949c287e7bff9  <= I666da645400344644e848ee6f7592d3c;
                    If3b234f8485412e76e5cc497b7c3a6f7  <=  0;
                end else begin
                    I4da324410e88d8c9738949c287e7bff9  <=  ~I666da645400344644e848ee6f7592d3c + 1;
                    If3b234f8485412e76e5cc497b7c3a6f7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3ade7e345432319c1a9c91d4068b3ec9 == I5bb0ab59e3468a9a95b65bfe58acd6a5 ) begin
                    Ie24b89ee61bddac2f2bbf1b8b5dd437f  <= Ibafeadd691eee03f855ed657c01022c9;
                    I67c58e4de1a3413b77529f5374201308  <=  0;
                end else begin
                    Ie24b89ee61bddac2f2bbf1b8b5dd437f  <=  ~Ibafeadd691eee03f855ed657c01022c9 + 1;
                    I67c58e4de1a3413b77529f5374201308  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3ade7e345432319c1a9c91d4068b3ec9 == I3e9c216d05b6a9c1040616a42af371ff ) begin
                    I27b99df87eefd6fcd484ec321bb73dc7  <= I10ec5c43a3fb65273053063001307280;
                    I9ad9a905418216c83643eae11965f330  <=  0;
                end else begin
                    I27b99df87eefd6fcd484ec321bb73dc7  <=  ~I10ec5c43a3fb65273053063001307280 + 1;
                    I9ad9a905418216c83643eae11965f330  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I88aed46f6dad7a81006562a720670654 == I4902647240aca7d98844546130944322 ) begin
                    Iaac7f8ca30f4e74e1ae5016a222673d7  <= I05c778eb3588bdaccf714ba456f534c2;
                    I2f3232289260297dfb0cb36e42e459be  <=  0;
                end else begin
                    Iaac7f8ca30f4e74e1ae5016a222673d7  <=  ~I05c778eb3588bdaccf714ba456f534c2 + 1;
                    I2f3232289260297dfb0cb36e42e459be  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I88aed46f6dad7a81006562a720670654 == Ia4c22694be7c5db34c1b875db1e91ff3 ) begin
                    Id3076c8e12f28723096148d8cf91a13d  <= Icd11e8d97a6ac6c0a73e8adee1f98c4e;
                    I58525519bd3b6773ec9ebabdf2764f69  <=  0;
                end else begin
                    Id3076c8e12f28723096148d8cf91a13d  <=  ~Icd11e8d97a6ac6c0a73e8adee1f98c4e + 1;
                    I58525519bd3b6773ec9ebabdf2764f69  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I88aed46f6dad7a81006562a720670654 == I0760280d5f5f23d9e06752908f0bbd96 ) begin
                    Ib2e36c2d0a51f5b953b9f368f11bb295  <= If07c2223d4262e22cca9b77c3ed5ee01;
                    I0e369759d6a2e5df5cd4fe6765ef8436  <=  0;
                end else begin
                    Ib2e36c2d0a51f5b953b9f368f11bb295  <=  ~If07c2223d4262e22cca9b77c3ed5ee01 + 1;
                    I0e369759d6a2e5df5cd4fe6765ef8436  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I88aed46f6dad7a81006562a720670654 == Ic807e0ddc985cffca6a389b468aeae49 ) begin
                    I9ef5138c78fee50aeb2568def8bc62a0  <= If0c8ce0ff66fe2806448f1c819d58ec8;
                    If155fcdeb6ebdce7305bf57a5e8fc426  <=  0;
                end else begin
                    I9ef5138c78fee50aeb2568def8bc62a0  <=  ~If0c8ce0ff66fe2806448f1c819d58ec8 + 1;
                    If155fcdeb6ebdce7305bf57a5e8fc426  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I79e574dc9c7e18b695c9a2619b71b995 == I9e3643f805ebd6623b9ab7ab41c41ec2 ) begin
                    Ic1cac944a0ed80e5b6e3821e8451045d  <= Iccdc2371dfd9fda3e506adc2b1681ba3;
                    I53e38457ad9a8a8244c9a2dd06034f60  <=  0;
                end else begin
                    Ic1cac944a0ed80e5b6e3821e8451045d  <=  ~Iccdc2371dfd9fda3e506adc2b1681ba3 + 1;
                    I53e38457ad9a8a8244c9a2dd06034f60  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I79e574dc9c7e18b695c9a2619b71b995 == I0dcf2ac5c06f517ea62c1ccd5acd9298 ) begin
                    I915f18e8333d52f6ec4162fe35317d17  <= I26e61dca9d045c4661b97afe346152c8;
                    I0cdf5ba9765cb28f2718129218794ec3  <=  0;
                end else begin
                    I915f18e8333d52f6ec4162fe35317d17  <=  ~I26e61dca9d045c4661b97afe346152c8 + 1;
                    I0cdf5ba9765cb28f2718129218794ec3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I79e574dc9c7e18b695c9a2619b71b995 == I26879becf6ee094c9b8b4969c9377af7 ) begin
                    Idbcf9e41a431a42028cc99d6be0c46da  <= Id488d650b86f5def0668f4a1ef841b6a;
                    Ic8e633425dff5441ceaa669bdd924077  <=  0;
                end else begin
                    Idbcf9e41a431a42028cc99d6be0c46da  <=  ~Id488d650b86f5def0668f4a1ef841b6a + 1;
                    Ic8e633425dff5441ceaa669bdd924077  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I79e574dc9c7e18b695c9a2619b71b995 == I3daa291236c162f58fdb9587a880dddb ) begin
                    Ic46dd35355bcd4470886fbd416b3c75c  <= I479365266255d2228ecd86c350e8d38b;
                    Ie7efb37f21bcddfe6cb7969533bbaca7  <=  0;
                end else begin
                    Ic46dd35355bcd4470886fbd416b3c75c  <=  ~I479365266255d2228ecd86c350e8d38b + 1;
                    Ie7efb37f21bcddfe6cb7969533bbaca7  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I800ef583bec1d46d3d4ffdea6b312ef9 == I2e150157b54bedd2bc6d31435e29af0e ) begin
                    I0765c8beae32257c6c37dabd94cbab7c  <= I08d9c488fd85db45344e649699196263;
                    Ie5a9f440574d20f6047c0ce556bc8477  <=  0;
                end else begin
                    I0765c8beae32257c6c37dabd94cbab7c  <=  ~I08d9c488fd85db45344e649699196263 + 1;
                    Ie5a9f440574d20f6047c0ce556bc8477  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I800ef583bec1d46d3d4ffdea6b312ef9 == If392bba16edcc39c846dc23bdf59f976 ) begin
                    Ibc002286423e5ddf50b8ea25ea1b3377  <= Icde86d0ead44385b07e9a29057417417;
                    I8fb0748ba8138a9188a557fcf752a055  <=  0;
                end else begin
                    Ibc002286423e5ddf50b8ea25ea1b3377  <=  ~Icde86d0ead44385b07e9a29057417417 + 1;
                    I8fb0748ba8138a9188a557fcf752a055  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I800ef583bec1d46d3d4ffdea6b312ef9 == Id0838a2f54127e6e86536294821b8fd2 ) begin
                    I714b85ebaccb1e11d16d53cf6bcf65b9  <= I21feecd24d912ef3d0aec0e375958f3f;
                    If6261c7d9d9c1b95edf08322eac2332e  <=  0;
                end else begin
                    I714b85ebaccb1e11d16d53cf6bcf65b9  <=  ~I21feecd24d912ef3d0aec0e375958f3f + 1;
                    If6261c7d9d9c1b95edf08322eac2332e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I800ef583bec1d46d3d4ffdea6b312ef9 == I3d11d3dc5ad053fd7a82b00d4ab4b180 ) begin
                    I864ca16e4e93b435a94fb012d995c7e5  <= I59f419b3bc183a5fe743be3878fac587;
                    Ib9f5522d41ddd9087096bb10ce7f5e23  <=  0;
                end else begin
                    I864ca16e4e93b435a94fb012d995c7e5  <=  ~I59f419b3bc183a5fe743be3878fac587 + 1;
                    Ib9f5522d41ddd9087096bb10ce7f5e23  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56cc5cd6d0a5a4e4601fd48e838fdaf3 == I1f67b8b8a325071662e006b730b1cc8a ) begin
                    I227ef7de18494a9f62b2e8cf37687840  <= Ib0804d8bdda49ecd0024300eed52be53;
                    I686a59acf3c8d19e90c2060b7db4be8f  <=  0;
                end else begin
                    I227ef7de18494a9f62b2e8cf37687840  <=  ~Ib0804d8bdda49ecd0024300eed52be53 + 1;
                    I686a59acf3c8d19e90c2060b7db4be8f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56cc5cd6d0a5a4e4601fd48e838fdaf3 == Icd7c05e9200f346555aa6b82827ad164 ) begin
                    I535a78cff546aed9fbd1d79827d56fe6  <= I37b0efdee34647a5111d698a5a80f367;
                    I73ba52dc87f86c76035540575994a224  <=  0;
                end else begin
                    I535a78cff546aed9fbd1d79827d56fe6  <=  ~I37b0efdee34647a5111d698a5a80f367 + 1;
                    I73ba52dc87f86c76035540575994a224  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56cc5cd6d0a5a4e4601fd48e838fdaf3 == Id136b4b678027d89c31614cd5baa6282 ) begin
                    I90cf52bd1332ea1b955e8c193b670218  <= Id382a04e94d0749d0858041bdc5861be;
                    I5947a59182e394e4b2f84b68ffd7bccc  <=  0;
                end else begin
                    I90cf52bd1332ea1b955e8c193b670218  <=  ~Id382a04e94d0749d0858041bdc5861be + 1;
                    I5947a59182e394e4b2f84b68ffd7bccc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56cc5cd6d0a5a4e4601fd48e838fdaf3 == I08dad437a9b452f65231279ae25ab7e1 ) begin
                    If7dc2cec6ded3b32d42281d08e871513  <= I368be992a21201268c41506396dcdcf6;
                    I006c14dc1c5be7dd3c5e1e5dcce08c21  <=  0;
                end else begin
                    If7dc2cec6ded3b32d42281d08e871513  <=  ~I368be992a21201268c41506396dcdcf6 + 1;
                    I006c14dc1c5be7dd3c5e1e5dcce08c21  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I21047a3955b8b89bdb9013d571b2bd0d == Ief01dd5ab84a9f9b05e48b07e0d1ed54 ) begin
                    Iee43875ccb00a79e67acbd3e12cb516d  <= I603a008893b5196d9f273b47a9d63144;
                    Iee841700cb259de93cbbfb47e828e1f4  <=  0;
                end else begin
                    Iee43875ccb00a79e67acbd3e12cb516d  <=  ~I603a008893b5196d9f273b47a9d63144 + 1;
                    Iee841700cb259de93cbbfb47e828e1f4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I21047a3955b8b89bdb9013d571b2bd0d == Iba8886370777ea357fd7c1e13bf03cd2 ) begin
                    I7aaad9fdd239670e028a896695c01216  <= Ie70d3a768bc09ddff6ac68aaba7d9f2c;
                    I71e36dabaef7951e59fc8b08da50003d  <=  0;
                end else begin
                    I7aaad9fdd239670e028a896695c01216  <=  ~Ie70d3a768bc09ddff6ac68aaba7d9f2c + 1;
                    I71e36dabaef7951e59fc8b08da50003d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I21047a3955b8b89bdb9013d571b2bd0d == I9e1e97a64e15a82443cc946178c11d52 ) begin
                    I4a992ed2550a3c5b346158ffe18c255d  <= Ifb8bd837ada3d8ed5116db29da82d2a9;
                    I323df8d18a73cd3947512f8a2c41b323  <=  0;
                end else begin
                    I4a992ed2550a3c5b346158ffe18c255d  <=  ~Ifb8bd837ada3d8ed5116db29da82d2a9 + 1;
                    I323df8d18a73cd3947512f8a2c41b323  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I21047a3955b8b89bdb9013d571b2bd0d == Ib830e17254cac0158be2b443e3dd4d43 ) begin
                    Ib2eb28843cf201e8c6f8900b7029d42d  <= I978b93d46e20cb3eda70e5a976d62348;
                    I30604b84bad8b4bba6d340cf020ca901  <=  0;
                end else begin
                    Ib2eb28843cf201e8c6f8900b7029d42d  <=  ~I978b93d46e20cb3eda70e5a976d62348 + 1;
                    I30604b84bad8b4bba6d340cf020ca901  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56eb529a34b484cd20e29958cd6878eb == I819741033c6737000bcf4a07a78e0938 ) begin
                    Ic9a5b2c8aee24c3fbc7e92b8fdaed5dc  <= Ib404040d4fb58f47f245184c3be01789;
                    Ib436620d6352c9ad5fa1d1fb5083de7a  <=  0;
                end else begin
                    Ic9a5b2c8aee24c3fbc7e92b8fdaed5dc  <=  ~Ib404040d4fb58f47f245184c3be01789 + 1;
                    Ib436620d6352c9ad5fa1d1fb5083de7a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56eb529a34b484cd20e29958cd6878eb == Ief41b57c092906a598c1cdcfea9b1062 ) begin
                    I6996efa8115f38da03518dcb7dd42a4d  <= I9c664265c53ebffaad097b70ff3cbbce;
                    I0722db2c7497d82a0ee09a109f698250  <=  0;
                end else begin
                    I6996efa8115f38da03518dcb7dd42a4d  <=  ~I9c664265c53ebffaad097b70ff3cbbce + 1;
                    I0722db2c7497d82a0ee09a109f698250  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56eb529a34b484cd20e29958cd6878eb == Ibea5db121c78f1b6d5288231ef59d04b ) begin
                    I1c4bf7954b4bd5f4e9c176a3ae1fc28a  <= I781306c6b1ce0741d9c2fa06865f7a19;
                    I34fe1fee7604351d37636552ecb32d8d  <=  0;
                end else begin
                    I1c4bf7954b4bd5f4e9c176a3ae1fc28a  <=  ~I781306c6b1ce0741d9c2fa06865f7a19 + 1;
                    I34fe1fee7604351d37636552ecb32d8d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I56eb529a34b484cd20e29958cd6878eb == If9d3ee7956572ceb26e7d60077de7e00 ) begin
                    I55d0fd8eda9c128cacdebab55a8dda5b  <= I16fa2e3dc0b3eddbc72811b51d6ac8ed;
                    Ie9ca773a78e9592fc49a7c590a3afee1  <=  0;
                end else begin
                    I55d0fd8eda9c128cacdebab55a8dda5b  <=  ~I16fa2e3dc0b3eddbc72811b51d6ac8ed + 1;
                    Ie9ca773a78e9592fc49a7c590a3afee1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I74588df6399af2c1112e3fa557e89e17 == I46fa901f3606f4d2ef11e13cdf029826 ) begin
                    I02fcd92b426929f24b9a8c063a56c0ed  <= Ia6f232495726806d01b702b0e248b2f2;
                    I023b8de48fefb0b45bed81ada503d779  <=  0;
                end else begin
                    I02fcd92b426929f24b9a8c063a56c0ed  <=  ~Ia6f232495726806d01b702b0e248b2f2 + 1;
                    I023b8de48fefb0b45bed81ada503d779  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I74588df6399af2c1112e3fa557e89e17 == I9918607fc0fdd746a6830800696a9439 ) begin
                    I3202a0ce45afe072eb955cd6e0789cd6  <= I66b3734060600caa45d699508c5083d2;
                    Id0ac1f9bcd5fa52b3b0536f0c831d504  <=  0;
                end else begin
                    I3202a0ce45afe072eb955cd6e0789cd6  <=  ~I66b3734060600caa45d699508c5083d2 + 1;
                    Id0ac1f9bcd5fa52b3b0536f0c831d504  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I74588df6399af2c1112e3fa557e89e17 == Iac50ab3381392442d8e7f18bd9ecacd8 ) begin
                    I06c82466a2ca646abb62bcaad3d63748  <= I85fae6b23d086235a94a0162e2fb5310;
                    Ic5c3ce39ad2fd88b6a26e639e390155d  <=  0;
                end else begin
                    I06c82466a2ca646abb62bcaad3d63748  <=  ~I85fae6b23d086235a94a0162e2fb5310 + 1;
                    Ic5c3ce39ad2fd88b6a26e639e390155d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I74588df6399af2c1112e3fa557e89e17 == Ie8bd9deffa3345851a9ff645b5bd1ddf ) begin
                    I23af695cf96a03638f0c1ef719d8d530  <= I8d6443d1be42203cb834345ae7e5aff5;
                    I80a34c662ed81f7d38d3055d470a1d1d  <=  0;
                end else begin
                    I23af695cf96a03638f0c1ef719d8d530  <=  ~I8d6443d1be42203cb834345ae7e5aff5 + 1;
                    I80a34c662ed81f7d38d3055d470a1d1d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic8eae1a92f46db040eb22d726c3a0e6d == Ia7d6b9edd50a4046aab863855f9491ee ) begin
                    Ie20b7fc4110631c1da7de4c7f38e2581  <= I717332b7f76e9caf9351f1aa69b72a12;
                    I0552127e741bcac86d4ef3994bf8830a  <=  0;
                end else begin
                    Ie20b7fc4110631c1da7de4c7f38e2581  <=  ~I717332b7f76e9caf9351f1aa69b72a12 + 1;
                    I0552127e741bcac86d4ef3994bf8830a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic8eae1a92f46db040eb22d726c3a0e6d == If8c22f4e0850faaa35f617a99c827f84 ) begin
                    Ic6983ef65e0de21992fa0b90ddbdce9d  <= Ieebd34db071409288f489129b70ab599;
                    Idef88c7c7169dae7b6d14e0edb17f47d  <=  0;
                end else begin
                    Ic6983ef65e0de21992fa0b90ddbdce9d  <=  ~Ieebd34db071409288f489129b70ab599 + 1;
                    Idef88c7c7169dae7b6d14e0edb17f47d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic8eae1a92f46db040eb22d726c3a0e6d == Iee22d62b28aee7dfc6c9304c92214e55 ) begin
                    Ie7c2317cef621a89ad24c8b5bc79a39c  <= I917c874137d64a9a495335c8f8ef5374;
                    I6f2e27ee85aad612520efe0e53f05aac  <=  0;
                end else begin
                    Ie7c2317cef621a89ad24c8b5bc79a39c  <=  ~I917c874137d64a9a495335c8f8ef5374 + 1;
                    I6f2e27ee85aad612520efe0e53f05aac  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ic8eae1a92f46db040eb22d726c3a0e6d == Idd235ad7cda4d67de5992f50db3b8de3 ) begin
                    Ic58955d8604cb1a6a20a199372d44774  <= I15fb4fb838d4a614c468f7d49261bda3;
                    Ia9afdb2578f40035f59aabad30a7e156  <=  0;
                end else begin
                    Ic58955d8604cb1a6a20a199372d44774  <=  ~I15fb4fb838d4a614c468f7d49261bda3 + 1;
                    Ia9afdb2578f40035f59aabad30a7e156  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I854a15bc7e9728b01c9a1960f6248dc9 == I6bb6fc0f5773f1386ac5af0688f224db ) begin
                    I8198473d2a666821cdf398dcf1b0fdc1  <= I2eb093d2a38ba8cf4be47d1d7f54ecc4;
                    I3c07ba2d2d09f45d52fbfe66bc54975f  <=  0;
                end else begin
                    I8198473d2a666821cdf398dcf1b0fdc1  <=  ~I2eb093d2a38ba8cf4be47d1d7f54ecc4 + 1;
                    I3c07ba2d2d09f45d52fbfe66bc54975f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I854a15bc7e9728b01c9a1960f6248dc9 == If44d50ac2bf54fad8236b3fcd9484792 ) begin
                    Ic60bdcbc8a55bc760e52c37aa3030001  <= I8f9affdc5cda0fecc35dd15fc5aeb244;
                    I77a2d8cfbb2e6f050545e2865b514205  <=  0;
                end else begin
                    Ic60bdcbc8a55bc760e52c37aa3030001  <=  ~I8f9affdc5cda0fecc35dd15fc5aeb244 + 1;
                    I77a2d8cfbb2e6f050545e2865b514205  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I854a15bc7e9728b01c9a1960f6248dc9 == I9039a46d1a19d43e6c1cb3f0c162efb1 ) begin
                    I987cca9a9fcbe4b617a7e524476431be  <= I615a443d49d1479338d033d2a2cab51f;
                    If126c59dab3d743d2451279fc184182d  <=  0;
                end else begin
                    I987cca9a9fcbe4b617a7e524476431be  <=  ~I615a443d49d1479338d033d2a2cab51f + 1;
                    If126c59dab3d743d2451279fc184182d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I854a15bc7e9728b01c9a1960f6248dc9 == Ib3c48b1a31a7198cc8d4fdd10d0c2db8 ) begin
                    I765c7209f3c7173362057fdb60aab732  <= I0635a3270a9653ca0f23c116fd5b2f97;
                    If745dbf2f0d756857eff51da036067fe  <=  0;
                end else begin
                    I765c7209f3c7173362057fdb60aab732  <=  ~I0635a3270a9653ca0f23c116fd5b2f97 + 1;
                    If745dbf2f0d756857eff51da036067fe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iae332cfd000fd0529684ab787041b5dc == If37efa97b30f1c80267e986fc90f759b ) begin
                    I2c117c8ea4060a5094453cc6140c9bb6  <= I93a7c75ebce8fbf4c613b4d11dc98b72;
                    I22231ac2204ad703262885231f7451e8  <=  0;
                end else begin
                    I2c117c8ea4060a5094453cc6140c9bb6  <=  ~I93a7c75ebce8fbf4c613b4d11dc98b72 + 1;
                    I22231ac2204ad703262885231f7451e8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iae332cfd000fd0529684ab787041b5dc == I42e35cda79f11acac889996660ec32ab ) begin
                    I56a6be4115d52bd49fc003b164fbcdb0  <= I39334aa9d55bcc001ece37ce2a6c329c;
                    I4e1e119c87f56b39ec6ddab9b160430d  <=  0;
                end else begin
                    I56a6be4115d52bd49fc003b164fbcdb0  <=  ~I39334aa9d55bcc001ece37ce2a6c329c + 1;
                    I4e1e119c87f56b39ec6ddab9b160430d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iae332cfd000fd0529684ab787041b5dc == I0ac3076614fbc543f41c76c6be389a37 ) begin
                    Ib834a7e4f3a491e351e2e49d809d2448  <= I07e328d23da9383a296ecb03679ec74b;
                    I9d9cc96988bd0af2b2c8682af3779794  <=  0;
                end else begin
                    Ib834a7e4f3a491e351e2e49d809d2448  <=  ~I07e328d23da9383a296ecb03679ec74b + 1;
                    I9d9cc96988bd0af2b2c8682af3779794  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iae332cfd000fd0529684ab787041b5dc == Iefae454b50cfb5b83c8016d5826e7670 ) begin
                    Ifdcb28209b39b8d99c2eb00a72921a75  <= I8a6e1eace6152af5c98c415804cb60fa;
                    I027210d36e2ae38a39746ac6fde3129a  <=  0;
                end else begin
                    Ifdcb28209b39b8d99c2eb00a72921a75  <=  ~I8a6e1eace6152af5c98c415804cb60fa + 1;
                    I027210d36e2ae38a39746ac6fde3129a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I70148fe95244eebf7f0ec953703398de == I86cd5db563b397776c52a89f0b44e442 ) begin
                    Id721a94e50637fa39c5bf6124ecfae6f  <= I6ed4d6c350e8691b3a12ab51419cfa65;
                    I28e32abf786d964b95d72bc17425a90f  <=  0;
                end else begin
                    Id721a94e50637fa39c5bf6124ecfae6f  <=  ~I6ed4d6c350e8691b3a12ab51419cfa65 + 1;
                    I28e32abf786d964b95d72bc17425a90f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I70148fe95244eebf7f0ec953703398de == Ibbf7f6c104c9f3163fc8d6b8a33ff5fe ) begin
                    I72ee7b62c165dc693cc6b5185970f7f5  <= Ie2b9ed680dac51ac866cb830ca17ef84;
                    Id29266756e91fa3c40480f9cf22f1671  <=  0;
                end else begin
                    I72ee7b62c165dc693cc6b5185970f7f5  <=  ~Ie2b9ed680dac51ac866cb830ca17ef84 + 1;
                    Id29266756e91fa3c40480f9cf22f1671  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I70148fe95244eebf7f0ec953703398de == Ife8ac54e4431329086b20d2111eb4f28 ) begin
                    I564ae36637e0cd6a8a06289e95823572  <= Ie439b520bbb0c8b29a5ecea167acb1c9;
                    Iad31d6f7d366c849222593883210e817  <=  0;
                end else begin
                    I564ae36637e0cd6a8a06289e95823572  <=  ~Ie439b520bbb0c8b29a5ecea167acb1c9 + 1;
                    Iad31d6f7d366c849222593883210e817  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I70148fe95244eebf7f0ec953703398de == I38c2a0e463853ac84b1f4e5c92f44243 ) begin
                    I085e99650c86078bf02f1b2aed141add  <= I9f8ef3295578acf5b0a42d074a15a70b;
                    I495d2cfe02637adf0bde6dd48201cedc  <=  0;
                end else begin
                    I085e99650c86078bf02f1b2aed141add  <=  ~I9f8ef3295578acf5b0a42d074a15a70b + 1;
                    I495d2cfe02637adf0bde6dd48201cedc  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24ee2d953e65fefdc73b3d3c4c0ddd05 == Ib73515d47a61e4a795005e8ae6bb2968 ) begin
                    Ie4e63cba44dee9885eeae32cc844c3f5  <= Ief01b06341d489e36ee344fd52084ccf;
                    I544225b6c571710d59f804f082f475c8  <=  0;
                end else begin
                    Ie4e63cba44dee9885eeae32cc844c3f5  <=  ~Ief01b06341d489e36ee344fd52084ccf + 1;
                    I544225b6c571710d59f804f082f475c8  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24ee2d953e65fefdc73b3d3c4c0ddd05 == I48b52a0f686c64c91c6ef4b1ca47593f ) begin
                    Ic054b062712da78ddd4a148bafeb1a0d  <= I3b72a085b104e17dca3d8b2824f84e97;
                    I6f7ff2aeffdfe5bd4090ecd655ff5aa2  <=  0;
                end else begin
                    Ic054b062712da78ddd4a148bafeb1a0d  <=  ~I3b72a085b104e17dca3d8b2824f84e97 + 1;
                    I6f7ff2aeffdfe5bd4090ecd655ff5aa2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24ee2d953e65fefdc73b3d3c4c0ddd05 == I9ed8d0fadbdab4e176b2d03549e41c91 ) begin
                    I81b01fc018ad1c79ec03a123763e95d9  <= I5e1f41e23887493db1d723e1e2cbd996;
                    I1783da96203ac6a00cd2e8f2dfe1ac34  <=  0;
                end else begin
                    I81b01fc018ad1c79ec03a123763e95d9  <=  ~I5e1f41e23887493db1d723e1e2cbd996 + 1;
                    I1783da96203ac6a00cd2e8f2dfe1ac34  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24ee2d953e65fefdc73b3d3c4c0ddd05 == Ibed24a9317d456b1a27bf71649c9a751 ) begin
                    I1d38ff144c3dcfe4c04778e50a044d5e  <= I0e6f4c7bdc39bd22833f3d9fcfa55f1d;
                    I00ae9e980c05d6d55570d92582a80410  <=  0;
                end else begin
                    I1d38ff144c3dcfe4c04778e50a044d5e  <=  ~I0e6f4c7bdc39bd22833f3d9fcfa55f1d + 1;
                    I00ae9e980c05d6d55570d92582a80410  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3a5f8eec283fd4f682b5d0f909b051c == If6b0b5b913b2f16e0354a62459f87487 ) begin
                    I2e31a90886f87907d19d0c034caeee9c  <= Ie346802a8898b4b075be289e062b462c;
                    I86282458466a079a1063e068011d58eb  <=  0;
                end else begin
                    I2e31a90886f87907d19d0c034caeee9c  <=  ~Ie346802a8898b4b075be289e062b462c + 1;
                    I86282458466a079a1063e068011d58eb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3a5f8eec283fd4f682b5d0f909b051c == I6cf5556c5887ad4d2f85b26aefe2aabf ) begin
                    I7c48130cd79566b1f1e30b7c709ee5cb  <= I82ea6f21706a97166ef11af548e80392;
                    I7dcde2729bcd8e63b86dcac06325887b  <=  0;
                end else begin
                    I7c48130cd79566b1f1e30b7c709ee5cb  <=  ~I82ea6f21706a97166ef11af548e80392 + 1;
                    I7dcde2729bcd8e63b86dcac06325887b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3a5f8eec283fd4f682b5d0f909b051c == I4fa8769d910cc70e158a0b649ce1e1d4 ) begin
                    I3868c6ed60d1f0ef9d3ad98e91931acf  <= I5f38764f6ecc2dcd1fdd5316102f1f82;
                    I31ca3f6f5d61b73718bbd9c19f7fd53b  <=  0;
                end else begin
                    I3868c6ed60d1f0ef9d3ad98e91931acf  <=  ~I5f38764f6ecc2dcd1fdd5316102f1f82 + 1;
                    I31ca3f6f5d61b73718bbd9c19f7fd53b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie3a5f8eec283fd4f682b5d0f909b051c == If25316f70adbd92abb74b4338c63d7d0 ) begin
                    I7fa57873a108e5894f837bdf45979b8d  <= Id4034bf7a0e92a6c92d0187e00d3df99;
                    Ie01688869a15f6b506bc3fbdea78b6b0  <=  0;
                end else begin
                    I7fa57873a108e5894f837bdf45979b8d  <=  ~Id4034bf7a0e92a6c92d0187e00d3df99 + 1;
                    Ie01688869a15f6b506bc3fbdea78b6b0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I781d986d7fd6c2fec3a8cf3f29545174 == I38b3f467871a1646a7694cc6433b5c8b ) begin
                    I59d4025a86d065a84741dafb86b50cbd  <= I44692fd63388c57268ea9035a7e4c3ef;
                    Iff748fa3440e5d0f80969f64b10eca98  <=  0;
                end else begin
                    I59d4025a86d065a84741dafb86b50cbd  <=  ~I44692fd63388c57268ea9035a7e4c3ef + 1;
                    Iff748fa3440e5d0f80969f64b10eca98  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I781d986d7fd6c2fec3a8cf3f29545174 == I0c7ee025ebd05956c96fd50885d627c6 ) begin
                    Ib28a3fb3dcdea36c883c88b017fefa56  <= I0c2892a34e5236f1366959eadfd83825;
                    I85018196561b6ef22994dfff7e3a8b80  <=  0;
                end else begin
                    Ib28a3fb3dcdea36c883c88b017fefa56  <=  ~I0c2892a34e5236f1366959eadfd83825 + 1;
                    I85018196561b6ef22994dfff7e3a8b80  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I781d986d7fd6c2fec3a8cf3f29545174 == I680660d6ba504eb445d2588ecfa046bf ) begin
                    I91e4dca55e1a5d1d8ddee5c3bd1048bc  <= Iccef2754044e7066e191bc5e1a3805f1;
                    Ifff25101d23e8e0ac43d5f0507a34217  <=  0;
                end else begin
                    I91e4dca55e1a5d1d8ddee5c3bd1048bc  <=  ~Iccef2754044e7066e191bc5e1a3805f1 + 1;
                    Ifff25101d23e8e0ac43d5f0507a34217  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib4db8131350f8605e00907234aff901d == Ia861785bea48073ffcabfd97a16890de ) begin
                    I55dd62b8ff91323075533e896207c1e5  <= I8ace46f1c56cfb3f4773324e0f8cae58;
                    I261ed926e2e82b283ac24970f546a5fe  <=  0;
                end else begin
                    I55dd62b8ff91323075533e896207c1e5  <=  ~I8ace46f1c56cfb3f4773324e0f8cae58 + 1;
                    I261ed926e2e82b283ac24970f546a5fe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib4db8131350f8605e00907234aff901d == I8619e41804844cd4d98818cb8387c3a7 ) begin
                    Ia30ca84355bb976cd045e969b2862856  <= I94ec0139bd827ef5dce2c5ee9eb9aded;
                    Ibf081c14165822b88553a913ba320016  <=  0;
                end else begin
                    Ia30ca84355bb976cd045e969b2862856  <=  ~I94ec0139bd827ef5dce2c5ee9eb9aded + 1;
                    Ibf081c14165822b88553a913ba320016  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib4db8131350f8605e00907234aff901d == If916ac75b729dfffab3cf6b0029197ce ) begin
                    Ifa1359651fd7e160301261bdbb81b02c  <= Ied62b116607c549ff5918d5b95e2118f;
                    I595bd58339ea7427b88385a62835aab6  <=  0;
                end else begin
                    Ifa1359651fd7e160301261bdbb81b02c  <=  ~Ied62b116607c549ff5918d5b95e2118f + 1;
                    I595bd58339ea7427b88385a62835aab6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie093f0750b60d3aed75705637933f34c == Id4f85daa963c656cff69ca2a821247fa ) begin
                    I0b465f693268f6f56f52d41165bf66ef  <= I9efa5796297bc922bc5fe17f8319a515;
                    I41b82d4c805471097a0dd4f85615f990  <=  0;
                end else begin
                    I0b465f693268f6f56f52d41165bf66ef  <=  ~I9efa5796297bc922bc5fe17f8319a515 + 1;
                    I41b82d4c805471097a0dd4f85615f990  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie093f0750b60d3aed75705637933f34c == Ic39575e662d7843dcd7418a7e8cc4a75 ) begin
                    I3deffa3a53b31688f28dfbfa66571d0c  <= Ifa6908d8fda29713d7c1bbaa69b72b53;
                    Ie07ed8367e7b83324c539bddcb3b1dfd  <=  0;
                end else begin
                    I3deffa3a53b31688f28dfbfa66571d0c  <=  ~Ifa6908d8fda29713d7c1bbaa69b72b53 + 1;
                    Ie07ed8367e7b83324c539bddcb3b1dfd  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ie093f0750b60d3aed75705637933f34c == I7c445b4e53ebe960faa00a46e00d66b4 ) begin
                    Id40c9857a5bb6c8cdc616fe68d8dc39d  <= Ieb46857229186ce0391cddb2d30f434e;
                    I67ba6804ea940c34c7c588832272581e  <=  0;
                end else begin
                    Id40c9857a5bb6c8cdc616fe68d8dc39d  <=  ~Ieb46857229186ce0391cddb2d30f434e + 1;
                    I67ba6804ea940c34c7c588832272581e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id2fba7c1b3dc7a75a5e0d90494d56962 == Iede71af4d6ced16d85e2576f035cc712 ) begin
                    I26754124b13858a3b925cddca5cd8c5b  <= I67fa03f808026b38ca5b4e71e21588bf;
                    Ifb2d4794b0630c3cdecb6cd2d2b1b384  <=  0;
                end else begin
                    I26754124b13858a3b925cddca5cd8c5b  <=  ~I67fa03f808026b38ca5b4e71e21588bf + 1;
                    Ifb2d4794b0630c3cdecb6cd2d2b1b384  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id2fba7c1b3dc7a75a5e0d90494d56962 == Ifffbd3dc45d11e43be5de5a276300bd4 ) begin
                    I2ebc1a7d32a5457de4d35b6bb25507d1  <= I70938dfe09b0da9d87dafed6af3fa05c;
                    I9c6dda8e9e0d7e69032a1fb40684c87c  <=  0;
                end else begin
                    I2ebc1a7d32a5457de4d35b6bb25507d1  <=  ~I70938dfe09b0da9d87dafed6af3fa05c + 1;
                    I9c6dda8e9e0d7e69032a1fb40684c87c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Id2fba7c1b3dc7a75a5e0d90494d56962 == Ib7be21d644d545e6671098d3d8622fe0 ) begin
                    I77bf5b03fa300d1dbf8df5ca4acbed14  <= Iff30a4e14b6282e9ef92e7f58230b516;
                    Ie7d857b468dedb6b7a73fe918332ff1d  <=  0;
                end else begin
                    I77bf5b03fa300d1dbf8df5ca4acbed14  <=  ~Iff30a4e14b6282e9ef92e7f58230b516 + 1;
                    Ie7d857b468dedb6b7a73fe918332ff1d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ecee74c445711a376133636ef414666 == I1bcc55c2c22b349f421eac34341487c4 ) begin
                    I6c1c1e404f92fc80495e8e5d187934a6  <= I43e0faf8070869ab0528a7a4a5cdc103;
                    I34662a12c505be8abbe01cb690d117d5  <=  0;
                end else begin
                    I6c1c1e404f92fc80495e8e5d187934a6  <=  ~I43e0faf8070869ab0528a7a4a5cdc103 + 1;
                    I34662a12c505be8abbe01cb690d117d5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ecee74c445711a376133636ef414666 == I5117b588204bc017b2a94a6e1097df82 ) begin
                    I126a2b15cdc34d88d17ebacb3681625f  <= Ib2f0333fac7701ae4a5589d54005b8f3;
                    Idc13433074453a726e7a35789d7d27d2  <=  0;
                end else begin
                    I126a2b15cdc34d88d17ebacb3681625f  <=  ~Ib2f0333fac7701ae4a5589d54005b8f3 + 1;
                    Idc13433074453a726e7a35789d7d27d2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ecee74c445711a376133636ef414666 == I7c6e35ef749c858168d55bcabea9078b ) begin
                    I9c5ec8e21febe3ebe00c53ac8b21d1f1  <= Ie4e1491da700923e81b2c1a246e528b1;
                    Id16d40761b18218d4270c00db6d4eca2  <=  0;
                end else begin
                    I9c5ec8e21febe3ebe00c53ac8b21d1f1  <=  ~Ie4e1491da700923e81b2c1a246e528b1 + 1;
                    Id16d40761b18218d4270c00db6d4eca2  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ecee74c445711a376133636ef414666 == I84a9bd349a6cd85859437ad4f9e70693 ) begin
                    If27eaa7cc4d1b5d2b7a962b48f0919df  <= Ie8602467de2ece2013878a6b8d3129a1;
                    Ifac93c987a8fb9726d85b77a2e4c8bba  <=  0;
                end else begin
                    If27eaa7cc4d1b5d2b7a962b48f0919df  <=  ~Ie8602467de2ece2013878a6b8d3129a1 + 1;
                    Ifac93c987a8fb9726d85b77a2e4c8bba  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifb3cf6b88835d27220df837682c4dc93 == I27b66137a39cb30b8059289cf98f8a19 ) begin
                    Ic15f443512d68537f9764a3ba88334f6  <= I85c93c62f79b1703cb6928f96737cf27;
                    Id742302a78483bbb2852b002262ed33d  <=  0;
                end else begin
                    Ic15f443512d68537f9764a3ba88334f6  <=  ~I85c93c62f79b1703cb6928f96737cf27 + 1;
                    Id742302a78483bbb2852b002262ed33d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifb3cf6b88835d27220df837682c4dc93 == I89b31cd7510ff82f89398b8682f040f7 ) begin
                    I47b266262fb5a98f66706f460f1248e6  <= I3dc816ee6c2a818b32f6d4e1228704bf;
                    I2f87df8d48fe83aa0ce493d69aaa3d88  <=  0;
                end else begin
                    I47b266262fb5a98f66706f460f1248e6  <=  ~I3dc816ee6c2a818b32f6d4e1228704bf + 1;
                    I2f87df8d48fe83aa0ce493d69aaa3d88  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifb3cf6b88835d27220df837682c4dc93 == I801f6e47b9e4f6b6acfaf6f8369ea217 ) begin
                    Id301f31702270a4f8e9964e3a75e3d62  <= Id34d83701e815c01359bc5cd1b9c993c;
                    Ic4bb880cb9f8d5a6d1cbbdf7cd205470  <=  0;
                end else begin
                    Id301f31702270a4f8e9964e3a75e3d62  <=  ~Id34d83701e815c01359bc5cd1b9c993c + 1;
                    Ic4bb880cb9f8d5a6d1cbbdf7cd205470  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ifb3cf6b88835d27220df837682c4dc93 == I6f7db7eb1e5bc6d08ea9059ef7c31949 ) begin
                    I097ba3ae5a0232ae6aa35478635640b3  <= I0a20e3e26261ba558d681346649cf0b3;
                    I369ea36c9da8f4c9b93ee70f8d4c149f  <=  0;
                end else begin
                    I097ba3ae5a0232ae6aa35478635640b3  <=  ~I0a20e3e26261ba558d681346649cf0b3 + 1;
                    I369ea36c9da8f4c9b93ee70f8d4c149f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I386fbb3bd550891d682e137044e8773a == Idd01178431a1c4a53be45095dc897c33 ) begin
                    I3b65eb49005aee57f61279c5a172d158  <= I331c6e8dbe2ea1e2232f82766926d0e6;
                    I17f6c250d2d07a58ddde6d232a1ab5de  <=  0;
                end else begin
                    I3b65eb49005aee57f61279c5a172d158  <=  ~I331c6e8dbe2ea1e2232f82766926d0e6 + 1;
                    I17f6c250d2d07a58ddde6d232a1ab5de  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I386fbb3bd550891d682e137044e8773a == I64ae03b30dd467619e71498ce8126df4 ) begin
                    I8573059885be4373531275502affd59d  <= Ie27046fd2751357e4a81dc62086f00be;
                    Iba5b23512434eb51ec8679a798273551  <=  0;
                end else begin
                    I8573059885be4373531275502affd59d  <=  ~Ie27046fd2751357e4a81dc62086f00be + 1;
                    Iba5b23512434eb51ec8679a798273551  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I386fbb3bd550891d682e137044e8773a == I36eba1bdcf4eac1c5c4b458515ed3f6e ) begin
                    I627f9d9ac0c07ded7306fd14773fbee4  <= I0897ceba8201bc14a49ab30318183875;
                    I91a06282a09b01980f2e7be4ecd3a982  <=  0;
                end else begin
                    I627f9d9ac0c07ded7306fd14773fbee4  <=  ~I0897ceba8201bc14a49ab30318183875 + 1;
                    I91a06282a09b01980f2e7be4ecd3a982  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I386fbb3bd550891d682e137044e8773a == Ibb1a5ae8240913132795df9605e82ce8 ) begin
                    Ib559f45098803b21622fa96ade885abc  <= Ie7b15aa8ce2492bfb433894efeb967f3;
                    I1b928fa95275de94960b3e2b4d67338b  <=  0;
                end else begin
                    Ib559f45098803b21622fa96ade885abc  <=  ~Ie7b15aa8ce2492bfb433894efeb967f3 + 1;
                    I1b928fa95275de94960b3e2b4d67338b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7ede7d2e1c2730b3b71340b11e880f5b == I597865149cd8d3e173f8aed514cec357 ) begin
                    I10e294379879538ecbf65fd423e7355d  <= I255add08e982f701508a98db221e617d;
                    I6488c30acdb3b47d4d4ee7b5947abdfe  <=  0;
                end else begin
                    I10e294379879538ecbf65fd423e7355d  <=  ~I255add08e982f701508a98db221e617d + 1;
                    I6488c30acdb3b47d4d4ee7b5947abdfe  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7ede7d2e1c2730b3b71340b11e880f5b == I667f0a049c87ac48820b60b2346de1c4 ) begin
                    Ice861034cd3b2f3847f325dbc9f52d08  <= If7ca4919fa1449f38777f742ee1fb875;
                    I29a436013f98b750df592eb7d26d0d1e  <=  0;
                end else begin
                    Ice861034cd3b2f3847f325dbc9f52d08  <=  ~If7ca4919fa1449f38777f742ee1fb875 + 1;
                    I29a436013f98b750df592eb7d26d0d1e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7ede7d2e1c2730b3b71340b11e880f5b == Ieb1c4ec26a969a2c1cb60e0d1c67b5cf ) begin
                    If201eea7e0023bb17fe41dbb4b5ec076  <= I24cafcb5b9825321c54e84827a662fdc;
                    I6fb12e6f50ffa6e94c9d43a22681702c  <=  0;
                end else begin
                    If201eea7e0023bb17fe41dbb4b5ec076  <=  ~I24cafcb5b9825321c54e84827a662fdc + 1;
                    I6fb12e6f50ffa6e94c9d43a22681702c  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I7ede7d2e1c2730b3b71340b11e880f5b == Id3293a3ac3bb53134fade82ddb8aace1 ) begin
                    Ib15f9bf401d734008d6a2b9a00c572d1  <= I3ede71cb7cb39774aedb9889240a2462;
                    Ib3f42f17505d5c091c8c924bbc26d117  <=  0;
                end else begin
                    Ib15f9bf401d734008d6a2b9a00c572d1  <=  ~I3ede71cb7cb39774aedb9889240a2462 + 1;
                    Ib3f42f17505d5c091c8c924bbc26d117  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64c65fad4a7d958d625c783626808175 == If7ed4187de370efdc1b9798bb6b05232 ) begin
                    I581f4e137ec21e639eec32a1675f4750  <= I24da9598a6840d3ba7b12fe4f638219b;
                    Ia4c22a118187d5b2dd154a4371dc06d1  <=  0;
                end else begin
                    I581f4e137ec21e639eec32a1675f4750  <=  ~I24da9598a6840d3ba7b12fe4f638219b + 1;
                    Ia4c22a118187d5b2dd154a4371dc06d1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64c65fad4a7d958d625c783626808175 == Iefc40b941a682059aca6ac8abffe1cfb ) begin
                    Ib7ff7b93c88fc8d9bcd915f0c678acff  <= I0358ca8833007cec4ce5047db32ab7a3;
                    I1a87822c50f6a0ac5a5e96021ad49fb3  <=  0;
                end else begin
                    Ib7ff7b93c88fc8d9bcd915f0c678acff  <=  ~I0358ca8833007cec4ce5047db32ab7a3 + 1;
                    I1a87822c50f6a0ac5a5e96021ad49fb3  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64c65fad4a7d958d625c783626808175 == I746ebc4b00c09f116eb087dfed4bf89a ) begin
                    I34dc9dff97e78a2d711f75675944b0d1  <= I85b5354463c1c15f91ed67292da912c1;
                    I6addbc7c163ce97b3482277e76c5feaa  <=  0;
                end else begin
                    I34dc9dff97e78a2d711f75675944b0d1  <=  ~I85b5354463c1c15f91ed67292da912c1 + 1;
                    I6addbc7c163ce97b3482277e76c5feaa  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I64c65fad4a7d958d625c783626808175 == I69683a0683ab00462065f6c3069fb6f3 ) begin
                    I8bc35065fe56bb75e6595937aaf9ef2a  <= Ie93731739ace44811198d0fd95b04a6a;
                    I124c4374f19808abbdc401a3b85aec67  <=  0;
                end else begin
                    I8bc35065fe56bb75e6595937aaf9ef2a  <=  ~Ie93731739ace44811198d0fd95b04a6a + 1;
                    I124c4374f19808abbdc401a3b85aec67  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib2e0cd0a2b51c3a265bdd20834c0ed2d == I183ad57174d779bab96973fc5ba5efd9 ) begin
                    I1822ab8ed690d872380ef820dc4282fe  <= I464926faf4e005ad491b0bf93a365e07;
                    I162653d33938a4553978b08df208228b  <=  0;
                end else begin
                    I1822ab8ed690d872380ef820dc4282fe  <=  ~I464926faf4e005ad491b0bf93a365e07 + 1;
                    I162653d33938a4553978b08df208228b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib2e0cd0a2b51c3a265bdd20834c0ed2d == Ic4e5558ac995583236747a83b3f54f33 ) begin
                    I1a1965726584c6c91a7e20de63f0fce3  <= Icdaaccfead6f2d5ac2ce19caf1104d57;
                    I291a3bbec5669b8958c0ded154af1f89  <=  0;
                end else begin
                    I1a1965726584c6c91a7e20de63f0fce3  <=  ~Icdaaccfead6f2d5ac2ce19caf1104d57 + 1;
                    I291a3bbec5669b8958c0ded154af1f89  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib2e0cd0a2b51c3a265bdd20834c0ed2d == I12899b73e235f01bce4137c479f6b300 ) begin
                    I08c5dcac6674c1671b85d07a55a005b0  <= I916d6f9429f2b0cc1bd6fb900484cde5;
                    I53a1d11cce6e036ba3a23dcc29d1cc3e  <=  0;
                end else begin
                    I08c5dcac6674c1671b85d07a55a005b0  <=  ~I916d6f9429f2b0cc1bd6fb900484cde5 + 1;
                    I53a1d11cce6e036ba3a23dcc29d1cc3e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ib2e0cd0a2b51c3a265bdd20834c0ed2d == I8dc3438a0d2b1c000f2b581f9a7ee588 ) begin
                    I40d67287bf525ab2696c30755d6babd5  <= I0142f9b3d361a0d88522f1c5f54aca84;
                    I5fda5f3c582bb88cb7de87298d15194a  <=  0;
                end else begin
                    I40d67287bf525ab2696c30755d6babd5  <=  ~I0142f9b3d361a0d88522f1c5f54aca84 + 1;
                    I5fda5f3c582bb88cb7de87298d15194a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I67be0b66c8d0680eb23290a4b3885af3 == Ia589b25714c687f50bfa26ead5cfae55 ) begin
                    I60dc8e5b6204e3a5fa32e79c5cceae94  <= Ie6871983b4f81b5321519647e628bd0e;
                    Id3933d661bcebbc3584c9e437c96c89d  <=  0;
                end else begin
                    I60dc8e5b6204e3a5fa32e79c5cceae94  <=  ~Ie6871983b4f81b5321519647e628bd0e + 1;
                    Id3933d661bcebbc3584c9e437c96c89d  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I67be0b66c8d0680eb23290a4b3885af3 == I7e4263d478638c2f3127394328deea11 ) begin
                    I0074b447046d75787aa872d8167171aa  <= I17d7be125df22153fc1ed051d4e0770a;
                    I0d38a30070a5ae3e879c357c3dde88ea  <=  0;
                end else begin
                    I0074b447046d75787aa872d8167171aa  <=  ~I17d7be125df22153fc1ed051d4e0770a + 1;
                    I0d38a30070a5ae3e879c357c3dde88ea  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I67be0b66c8d0680eb23290a4b3885af3 == I1c432aa61cf7d02567ef990929a15696 ) begin
                    I384965816ec3b915b9b623ad68fcc4c9  <= I50b13959e06243e54fad2088eaf65aa7;
                    I928993ece796543b23fb83df8c250845  <=  0;
                end else begin
                    I384965816ec3b915b9b623ad68fcc4c9  <=  ~I50b13959e06243e54fad2088eaf65aa7 + 1;
                    I928993ece796543b23fb83df8c250845  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I67be0b66c8d0680eb23290a4b3885af3 == I64531ff978fb8892605f2b0dd8422873 ) begin
                    Ic0e2656bee7174384f7f952dbb9da619  <= I7a423d609b492f73d5a322849b4b1cce;
                    I226f8490438d72f58c43377c8e60fc34  <=  0;
                end else begin
                    Ic0e2656bee7174384f7f952dbb9da619  <=  ~I7a423d609b492f73d5a322849b4b1cce + 1;
                    I226f8490438d72f58c43377c8e60fc34  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I01148401f7d058614dc1ae6ed3c8bd94 == Ib8c44be17e150cbd0b49d41c060f95f1 ) begin
                    I4cc3b0546ddc14d78da59e4981a77b58  <= Iefec67e214d1868670a34a7297d4a1c8;
                    Idaefaba16ce80e24f16df683cc83d759  <=  0;
                end else begin
                    I4cc3b0546ddc14d78da59e4981a77b58  <=  ~Iefec67e214d1868670a34a7297d4a1c8 + 1;
                    Idaefaba16ce80e24f16df683cc83d759  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I01148401f7d058614dc1ae6ed3c8bd94 == Ic45b89f2b51ee014d9a0fb19a7ed7619 ) begin
                    I7b680caf7d0d94114fae1d96ba374e68  <= Iae7da7fdc002b635ce4285d6916d8156;
                    If1da75cd8208f606c1b121f441685cbb  <=  0;
                end else begin
                    I7b680caf7d0d94114fae1d96ba374e68  <=  ~Iae7da7fdc002b635ce4285d6916d8156 + 1;
                    If1da75cd8208f606c1b121f441685cbb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I01148401f7d058614dc1ae6ed3c8bd94 == I338e32162153b4ed5d991c44c38aca27 ) begin
                    I7f8986a922c03b6afb5786cd2e1d5288  <= Ic561e44b2caeae84df6720f1afa3e8f6;
                    Ib63f66960a3981879aad950588ea14be  <=  0;
                end else begin
                    I7f8986a922c03b6afb5786cd2e1d5288  <=  ~Ic561e44b2caeae84df6720f1afa3e8f6 + 1;
                    Ib63f66960a3981879aad950588ea14be  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I01148401f7d058614dc1ae6ed3c8bd94 == I06c60ff1b8b447112b28f71eb9e3944d ) begin
                    Ie7814643e3833736c0f54b39f91fe792  <= I5be062f5b52e104ca67e615ce75a7c80;
                    Ia2c2ecedc809186e3f9224a9aa4bf385  <=  0;
                end else begin
                    Ie7814643e3833736c0f54b39f91fe792  <=  ~I5be062f5b52e104ca67e615ce75a7c80 + 1;
                    Ia2c2ecedc809186e3f9224a9aa4bf385  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3394319c370daf6102be00d938d55769 == Ic2cc5a2da05052c4a68cadde2745b44e ) begin
                    Id1f0c95b85ee041818da4fd9b5466c7d  <= Iecdde23e34c34ee0055be41f44959a19;
                    I1fc189d6e8a90cc0033c6e690916de83  <=  0;
                end else begin
                    Id1f0c95b85ee041818da4fd9b5466c7d  <=  ~Iecdde23e34c34ee0055be41f44959a19 + 1;
                    I1fc189d6e8a90cc0033c6e690916de83  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3394319c370daf6102be00d938d55769 == I8073ab2d9dc1d68d0bb4694ff206995f ) begin
                    Iefa8421c0c908de69fccffbe22f40911  <= Ibe09be9cad0e56d5403868d072d7d628;
                    I7fa18d2c7159b9fda8957384ebca5700  <=  0;
                end else begin
                    Iefa8421c0c908de69fccffbe22f40911  <=  ~Ibe09be9cad0e56d5403868d072d7d628 + 1;
                    I7fa18d2c7159b9fda8957384ebca5700  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3394319c370daf6102be00d938d55769 == I6aec90f4d15da8590fe767c4facfe19b ) begin
                    I4319bf1bbb31debc7f58157b75025134  <= I464e1f3c13acaf466afb354a9b35ba0a;
                    I7ea0274f5b34aac64a17fa9171201a5a  <=  0;
                end else begin
                    I4319bf1bbb31debc7f58157b75025134  <=  ~I464e1f3c13acaf466afb354a9b35ba0a + 1;
                    I7ea0274f5b34aac64a17fa9171201a5a  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3394319c370daf6102be00d938d55769 == I39a8cf4c424841d2b367cb3a1207fe03 ) begin
                    I4a349021efeeda16b646979a959bff6e  <= I160a465c22073a53510e8a4c489c3321;
                    I8d26db6f54d068f798e2951701aebed1  <=  0;
                end else begin
                    I4a349021efeeda16b646979a959bff6e  <=  ~I160a465c22073a53510e8a4c489c3321 + 1;
                    I8d26db6f54d068f798e2951701aebed1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24d6a334dd15ccdea558f32cd029e6d1 == I031f3e2575360f675bed8e87a71755d7 ) begin
                    Iaae0c136077ecc36fc382a76abd550e7  <= I9e86d3e49827861b24f4fbeb308ad3a4;
                    I8fb8a6e1ab4647e8e1dda4da8b3ef3c6  <=  0;
                end else begin
                    Iaae0c136077ecc36fc382a76abd550e7  <=  ~I9e86d3e49827861b24f4fbeb308ad3a4 + 1;
                    I8fb8a6e1ab4647e8e1dda4da8b3ef3c6  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24d6a334dd15ccdea558f32cd029e6d1 == I40feba64660df64a02c3df651a2ca26c ) begin
                    I4a442564148493664046e7b38cc6cfe4  <= Ib96b7d796e20967e89a47e01bf424e59;
                    Ie4821dad77dec0567d64f7c1de7710af  <=  0;
                end else begin
                    I4a442564148493664046e7b38cc6cfe4  <=  ~Ib96b7d796e20967e89a47e01bf424e59 + 1;
                    Ie4821dad77dec0567d64f7c1de7710af  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24d6a334dd15ccdea558f32cd029e6d1 == I985f121a0212a4d64ca4a47c1c210b40 ) begin
                    I12cc5eec3de8ceb3ca084194d430d9a5  <= I565e666f6ba14b4c25e0dd402a3266e1;
                    Ic4d741a90fcc86f31eb3567d028eb27f  <=  0;
                end else begin
                    I12cc5eec3de8ceb3ca084194d430d9a5  <=  ~I565e666f6ba14b4c25e0dd402a3266e1 + 1;
                    Ic4d741a90fcc86f31eb3567d028eb27f  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I24d6a334dd15ccdea558f32cd029e6d1 == Id4ce64c9f467d1b1c4bc9099ab855db2 ) begin
                    I56db71b7df11c35080cbaee80c389c59  <= I97e8bac5becd5128bc70f3bb48f73e6c;
                    I1d2641b8888a0f7b4b78cae16779da75  <=  0;
                end else begin
                    I56db71b7df11c35080cbaee80c389c59  <=  ~I97e8bac5becd5128bc70f3bb48f73e6c + 1;
                    I1d2641b8888a0f7b4b78cae16779da75  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a41f68bca2d7edd1f5738c4fda8e73c == I01c6d49bf9698d7621a545481b129692 ) begin
                    Ifd1431230378775456efa4bdd5bfc397  <= Iced39475c6e5e3d8f36d2a5c5a80f146;
                    I48badf0536ab133751d4be1e0450fd81  <=  0;
                end else begin
                    Ifd1431230378775456efa4bdd5bfc397  <=  ~Iced39475c6e5e3d8f36d2a5c5a80f146 + 1;
                    I48badf0536ab133751d4be1e0450fd81  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a41f68bca2d7edd1f5738c4fda8e73c == I73164ee0df8db9282850f1b325afc7ae ) begin
                    I6f0cef6d870e38e5ba192463a3920818  <= Idcbd423c2b963c1f693dea2ddf428195;
                    I043ba9e5157ad18a4e466df0540b79ba  <=  0;
                end else begin
                    I6f0cef6d870e38e5ba192463a3920818  <=  ~Idcbd423c2b963c1f693dea2ddf428195 + 1;
                    I043ba9e5157ad18a4e466df0540b79ba  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a41f68bca2d7edd1f5738c4fda8e73c == Ic985d004f7feb36aaa6415dc7365e617 ) begin
                    I3ee87c05f23571b687611fdce84a1b91  <= If1640e294bdcc51ee12fca5b3a33be6d;
                    Ib9760b69084b2d4a3a93126e5da0f20b  <=  0;
                end else begin
                    I3ee87c05f23571b687611fdce84a1b91  <=  ~If1640e294bdcc51ee12fca5b3a33be6d + 1;
                    Ib9760b69084b2d4a3a93126e5da0f20b  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I3a41f68bca2d7edd1f5738c4fda8e73c == Ia09ac88781a570aead25d43447ff9afc ) begin
                    Ide521f7523b897bb6fb747202f730ac5  <= I4754c6c355e632d2ed1336b5a88c3b46;
                    I4978a011cb09d68ac2850e1f515d7e88  <=  0;
                end else begin
                    Ide521f7523b897bb6fb747202f730ac5  <=  ~I4754c6c355e632d2ed1336b5a88c3b46 + 1;
                    I4978a011cb09d68ac2850e1f515d7e88  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ef1784d165492f3482d14f475732451 == I17cb6dfd1374c74d63862703fa6665ce ) begin
                    I314b64e5fbbc14807fd7fe3c7bca101f  <= I1634d703ad5d6e58a97b13ef957bdbec;
                    Ib09ea18232dfca23f3f139438e6cb800  <=  0;
                end else begin
                    I314b64e5fbbc14807fd7fe3c7bca101f  <=  ~I1634d703ad5d6e58a97b13ef957bdbec + 1;
                    Ib09ea18232dfca23f3f139438e6cb800  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ef1784d165492f3482d14f475732451 == I6c05d39d4c7a50f019474562f741e591 ) begin
                    Id5ad2e12b160bc6a9f96f2524f849c8e  <= I804e1e6a01edeb780b0159ecae707b71;
                    If29c61ebd2b452efe995c212a76a77a0  <=  0;
                end else begin
                    Id5ad2e12b160bc6a9f96f2524f849c8e  <=  ~I804e1e6a01edeb780b0159ecae707b71 + 1;
                    If29c61ebd2b452efe995c212a76a77a0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ef1784d165492f3482d14f475732451 == I413638a340bf1e686e718453f1b243b6 ) begin
                    I2b2bf6d4e879b8f53b02f94f1e964344  <= Iea3c0f3c3c3017fe87a3b01647189fe0;
                    I60fa2e2b5dd8b0a99612d2f2f6c5c740  <=  0;
                end else begin
                    I2b2bf6d4e879b8f53b02f94f1e964344  <=  ~Iea3c0f3c3c3017fe87a3b01647189fe0 + 1;
                    I60fa2e2b5dd8b0a99612d2f2f6c5c740  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9ef1784d165492f3482d14f475732451 == I904a05d4a23c6d15438654f937811877 ) begin
                    Ic60cb038b4b90d8035059b1e06f8d765  <= I756b7d7e6bd3e71afa472e7e4727264a;
                    Ifc9b6cc64f5bf8bc685911bb28884a0e  <=  0;
                end else begin
                    Ic60cb038b4b90d8035059b1e06f8d765  <=  ~I756b7d7e6bd3e71afa472e7e4727264a + 1;
                    Ifc9b6cc64f5bf8bc685911bb28884a0e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9d9378337a77515a4e8d04fb88938808 == Iab36b17e472fde9a92c4dc5ebb75ca6c ) begin
                    I707e2d6d9807076bfc91417fb9e198e6  <= Ifbeae0a2acf80eda6ffd050d3bb07eb3;
                    I1aeaa36994ba29298931735d5a1237e0  <=  0;
                end else begin
                    I707e2d6d9807076bfc91417fb9e198e6  <=  ~Ifbeae0a2acf80eda6ffd050d3bb07eb3 + 1;
                    I1aeaa36994ba29298931735d5a1237e0  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9d9378337a77515a4e8d04fb88938808 == I4d265ef808b1e19fb1dcef26a6dd4204 ) begin
                    I49f5797b92e17562e6dfde42c20c7a37  <= I990ab4dcb70ee860c2c40f306ef314d3;
                    I415ed6a9802acf39be10b220ddb3ff66  <=  0;
                end else begin
                    I49f5797b92e17562e6dfde42c20c7a37  <=  ~I990ab4dcb70ee860c2c40f306ef314d3 + 1;
                    I415ed6a9802acf39be10b220ddb3ff66  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9d9378337a77515a4e8d04fb88938808 == I535542d9580a449d24a712ef814d5e58 ) begin
                    I0a9f0274dc61d574c40e0e2048fb0b9e  <= Ib131087ea9ccc4bd161c3f9ac2c72303;
                    I1c06321ed28c991ad2aa8a3725769dee  <=  0;
                end else begin
                    I0a9f0274dc61d574c40e0e2048fb0b9e  <=  ~Ib131087ea9ccc4bd161c3f9ac2c72303 + 1;
                    I1c06321ed28c991ad2aa8a3725769dee  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (I9d9378337a77515a4e8d04fb88938808 == I82298047310dc4da0ea3762c6a48e07f ) begin
                    I53ae3de5769255a9e69a2ae690d44ba9  <= I9a967ac9d11583faaa783984229aeb2c;
                    I198d5b5bf8f39f9bd6b2f4c993fd58ca  <=  0;
                end else begin
                    I53ae3de5769255a9e69a2ae690d44ba9  <=  ~I9a967ac9d11583faaa783984229aeb2c + 1;
                    I198d5b5bf8f39f9bd6b2f4c993fd58ca  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If0e20ef9aa69b77ae0e58ca3dfc9998f == I761dfdefbc96fec3c2ac79f0a1de18b7 ) begin
                    I1390f0ff082dbff11a64cdfcbe1b681d  <= Ib9921dfcf121e5f4ac4d8be83a868210;
                    I3bf64d0a85c83de954a286e6afa8f727  <=  0;
                end else begin
                    I1390f0ff082dbff11a64cdfcbe1b681d  <=  ~Ib9921dfcf121e5f4ac4d8be83a868210 + 1;
                    I3bf64d0a85c83de954a286e6afa8f727  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If0e20ef9aa69b77ae0e58ca3dfc9998f == Ib68e4d694df8e44519916724104f7962 ) begin
                    Id2f8816659d3881ee1b1d14668a53a08  <= If22d8fd45caed08b2c7cee8b7349700f;
                    I897c7fc822d490f69b531a8f749815f4  <=  0;
                end else begin
                    Id2f8816659d3881ee1b1d14668a53a08  <=  ~If22d8fd45caed08b2c7cee8b7349700f + 1;
                    I897c7fc822d490f69b531a8f749815f4  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If0e20ef9aa69b77ae0e58ca3dfc9998f == I3284ce21b5d114a7127917f8b261b21a ) begin
                    I286bacc5a8a77b89cb99dbb00962555b  <= Iabf029e67c7f827faf17b6518cd1bfa3;
                    I6c7cb10db83156b49d46fab38d0f9fc5  <=  0;
                end else begin
                    I286bacc5a8a77b89cb99dbb00962555b  <=  ~Iabf029e67c7f827faf17b6518cd1bfa3 + 1;
                    I6c7cb10db83156b49d46fab38d0f9fc5  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (If0e20ef9aa69b77ae0e58ca3dfc9998f == I30b857065185101e8e4cb0270e747cae ) begin
                    Icda8e8a6ba7607752ed282114a542b67  <= Iaeab83001c6285630e3404ae67227f46;
                    Ie47af3b071351ec683abe28b7fe2b642  <=  0;
                end else begin
                    Icda8e8a6ba7607752ed282114a542b67  <=  ~Iaeab83001c6285630e3404ae67227f46 + 1;
                    Ie47af3b071351ec683abe28b7fe2b642  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iec2cb48bb1b58f268bf164d5e8a8120f == If9be63889327fc1b68abc628c9a0a78d ) begin
                    I2da4a59f9a6bd71af95790a75b172df0  <= I53ac6d02d2bfc9aca9469148753070a7;
                    If2dd4df3af6446c05da4afdaa7e92cab  <=  0;
                end else begin
                    I2da4a59f9a6bd71af95790a75b172df0  <=  ~I53ac6d02d2bfc9aca9469148753070a7 + 1;
                    If2dd4df3af6446c05da4afdaa7e92cab  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iec2cb48bb1b58f268bf164d5e8a8120f == If0c3ec1e3a80a23b2506621ec2d9f02a ) begin
                    I1bcf01b7fde13919f5d7c4df4483e61c  <= I61992979f60b26d313efd1dc23bb54ab;
                    Iabf085ea078abe8748810e81a6d03cac  <=  0;
                end else begin
                    I1bcf01b7fde13919f5d7c4df4483e61c  <=  ~I61992979f60b26d313efd1dc23bb54ab + 1;
                    Iabf085ea078abe8748810e81a6d03cac  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iec2cb48bb1b58f268bf164d5e8a8120f == I2842882109b7ef022421ab185471ab33 ) begin
                    Id5f000c37734979d057f7887739a5615  <= I8b46b3f0835310114208963de7ac8e97;
                    Ia2ae348906a599a4d327ff1419315afb  <=  0;
                end else begin
                    Id5f000c37734979d057f7887739a5615  <=  ~I8b46b3f0835310114208963de7ac8e97 + 1;
                    Ia2ae348906a599a4d327ff1419315afb  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Iec2cb48bb1b58f268bf164d5e8a8120f == Iecb13253abbfb0a891a4e526f05841f3 ) begin
                    Ibccd7142ba951dadbeca13178458bb3a  <= Icda26ba6f5c7f77a80776b2c1bbc975d;
                    I18df34aea04ea7dc99fc918892bf8f0e  <=  0;
                end else begin
                    Ibccd7142ba951dadbeca13178458bb3a  <=  ~Icda26ba6f5c7f77a80776b2c1bbc975d + 1;
                    I18df34aea04ea7dc99fc918892bf8f0e  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia4ae7c98720d43a604f28dfc5dd67d50 == I899cefdf3938be01e93d011e046c1e49 ) begin
                    Ic1fe6b93bc8d517686ba430d3d1fe7ab  <= I0863565b3ae88137a2384750436f9e19;
                    I910749abcd809e1c730f27fb5e1ddab1  <=  0;
                end else begin
                    Ic1fe6b93bc8d517686ba430d3d1fe7ab  <=  ~I0863565b3ae88137a2384750436f9e19 + 1;
                    I910749abcd809e1c730f27fb5e1ddab1  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia4ae7c98720d43a604f28dfc5dd67d50 == Ib96a9bf253b178aa920a63c8493932fb ) begin
                    Ib1c8d1d733e91f052f6d6824e734b1e3  <= Id646110f8d09cd47dc7695e05f73efc6;
                    Iae95ea2f32f53a5060c0199c8196d681  <=  0;
                end else begin
                    Ib1c8d1d733e91f052f6d6824e734b1e3  <=  ~Id646110f8d09cd47dc7695e05f73efc6 + 1;
                    Iae95ea2f32f53a5060c0199c8196d681  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia4ae7c98720d43a604f28dfc5dd67d50 == I5f534382562a3394100cdadb3ad1e0be ) begin
                    I08348d0a177e264af1a4769422878a06  <= I5999eef2304e579a3d47e4f15ba336e1;
                    I8c3d927ec93e73c5bca489a2f2b43f55  <=  0;
                end else begin
                    I08348d0a177e264af1a4769422878a06  <=  ~I5999eef2304e579a3d47e4f15ba336e1 + 1;
                    I8c3d927ec93e73c5bca489a2f2b43f55  <=  1;
                end
             end
             if (I92354deea988f3beb25bfba90735c6ac) begin
                if (Ia4ae7c98720d43a604f28dfc5dd67d50 == I137e343ba2386bbe31813bbe37e87dd9 ) begin
                    I2d2c2997dcc5167fc6ddc1e90f0ebc49  <= Idd302bdc6ff8368a6b73d53bbc8f8425;
                    Ib41ff881898782965734bb0cc333be79  <=  0;
                end else begin
                    I2d2c2997dcc5167fc6ddc1e90f0ebc49  <=  ~Idd302bdc6ff8368a6b73d53bbc8f8425 + 1;
                    Ib41ff881898782965734bb0cc333be79  <=  1;
                end
             end
       end
   end


   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
            I748f85f6680918a2e992df339b4b6558                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic93835a022c46b7aa00a465c407d7da2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I92cb615e2c439914e72ce001256518e4  <= 1'b0;
            I2e30088bf29cedd7debc15b1e6ec4ada        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iad799775eb657f8973e6dfcf70a9875c  <= 1'b0;
            I38f512bfb84094d1e92a10a345d5505f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifb064c69c7110c014593149ae69c75fb  <= 1'b0;
            I1e878f00f056f637625cb013a93325a8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7f7b30f2acbb8e31f50b58096b738254  <= 1'b0;
            I25db27464b31fee41ccd7a3cfe4d403e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iefe4099ff7e457f6b9fefc83e176c1a0  <= 1'b0;
            I19417a224c5cdf1211e9790aa29c4c5c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icddb43f9b760a4597a0bb637fb405616  <= 1'b0;
            I16dcafa854ea9c67d8a080feb2ba9166        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic76e72b434b47c10ebac3fac4ea50bde  <= 1'b0;
            I7f63338eee2663fbe61fffd248433310        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9eb87e62d23bc87d7cd82c0f329f247f  <= 1'b0;
            Icb1e3c56c8729c32d43c69710e345db2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2eac5b39c6f485c9ae0bd341f894633d  <= 1'b0;
            I6ece8e3c1e89613879336936f77d732f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I76992221b1edff5684c482df7ac4693d  <= 1'b0;
            I72a646ae7e32a16af0f5930a6e95b36a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iada5bc4a51dc1bf57bb9cca11326bdff  <= 1'b0;
            I7e72d119dd93a6ab05a23fde0a865866        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I364ed3f83c49626bc3b939e53524d9c7  <= 1'b0;
            Ied4fdf5805039cd2fcd042fd13755fdc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic2b000c3b2ca3beff2d427caab04701a  <= 1'b0;
            Id44c2293b765cff450dd1d747c47c1f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8e873fb2321eea82bb590a92411e2e2c  <= 1'b0;
            I8f4ed02f7aeb823b745040f7f3f43ac7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If4cb744ee52b6ae793431cd038069b57  <= 1'b0;
            I6488b9b8f405d7d81a4874fab2678102        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7741e239c16828889d488cc87647c154  <= 1'b0;
            Ifff612d16828ec907a348479e19ddf31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7979161aa1e2262ebea862004c387697  <= 1'b0;
            I268262076f22bc6b1507bc8f91b98a0a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic62fc602da3d16fe13d03a49a21269d0  <= 1'b0;
            If1f732841adb7c0cad1ba37c0f5fd517        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I94009bb7239be96243902ab0f0abea7e  <= 1'b0;
            I0df8a24f31c027756d248c3bd1b9bf7b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iae7b72abf4d3c536330a229e3836b441  <= 1'b0;
            I8ef901e733b12e76412eb36684e2b575        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie5d9cc18b2dd300132470f206452ff17  <= 1'b0;
            Ia48916a02f68b1b8f5fc7fece04677bb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7c791c854d0bc28e8dd787545f8fbda0  <= 1'b0;
            Ib0f57837099e3fdf1b908d78bcda4a43                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia37409944d9fdd3b16e7007e13d82a79        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5b177dd5c14ad082516b47f550875682  <= 1'b0;
            Idd65f149afe9d5f63ddaf34b82b11e95        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I55e4ad2d71a29ad63b4999d64ac0dc4f  <= 1'b0;
            If2886d560854faed32ebd8e33d868973        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I59c5da6338f431a626c86a065a355c35  <= 1'b0;
            I77778118bb3ea900c080754ff4c49c26        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia098bbeda8b755ece6b88eac83d03e55  <= 1'b0;
            I7292ed752d8741594d757730950feea4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie7470dd75b54d14038de19e4d3043ba9  <= 1'b0;
            I68cfd7868e061793ee8a41e69e80219b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie95662d4faf6b5a4cd5ecfa41697b983  <= 1'b0;
            I667ead814b303fca64ef047bb8246b19        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia1b617e3d141263b51e58c5ef0bd7a89  <= 1'b0;
            I4f25c7edb12e868cb5532e42b4ba5133        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If9a5d830e3ade0fd96b98f5949f165f0  <= 1'b0;
            I5aed2d82717f359bb5ac5a0ab91b7beb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id3de87169c440f95d406693ef77cacd6  <= 1'b0;
            I92835fd54631deaefa7b214e2c4b9bff        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3751f191f5009322acb7c9be4f8d7129  <= 1'b0;
            I67e067da565635fcff166e3a7d0c446b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic1927bb3335f6a28c0816eba12d3975e  <= 1'b0;
            Ifdb0f307b1b9458c0487a1574ccc094b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia659126b51468cfef48c97a135a71500  <= 1'b0;
            I5c6b7d143e42fd3b8bcdb7d7ed4da2c2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3c3c22bf63e55a81ae91b1dd1ef615a0  <= 1'b0;
            Ie679a21d0136a08cc5e6526e9f8d1843        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia62832d325f86160285c4d1a790a32cb  <= 1'b0;
            I611942a72a5e12f6afaea6bde6699ef6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I83c7d177eec2dad0a924557cdc91ba77  <= 1'b0;
            Ica9883c97f823a4491cbee5b45c43590        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7050adb9d06f767549b7f35c4679e391  <= 1'b0;
            I8e6addfc61f5bfb7af74fc2993639565        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I04aacd95d9e44657f616e01c9053f0fb  <= 1'b0;
            I9d53619f10e2a426f7297bbf7c81158a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2ff317d57f59747c4524ef4278d51092  <= 1'b0;
            I8a055c27778913287ad951183fa0d4d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8bd2a9d90074500698b302cb8db7f03a  <= 1'b0;
            I8f6ae5c80bb2f50084b5f5ee5ab0ffc3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3b8cdfb1440732ce98cd1676e05a2af1  <= 1'b0;
            I3db8b3a342e8e2f13a448246aa001c2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I671de3d408b5b783541663c7f1e3a6fa  <= 1'b0;
            Ibbee0996ea0f5e16b1f711345be7f2ae        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I446857735e680cae93a24dccb59b1924  <= 1'b0;
            If75e99660e3997f53f7b903bc366f47f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Idb777f1eb4c3cbba103b9b43f948ccf9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I77b05a8aa92c66a235195a66dc13c0cc  <= 1'b0;
            Id5e46b1f8844c7587f99d22170581a24        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie92110d19f4886cdfcfacd0920c06a4e  <= 1'b0;
            I67aadabd3cf49456cace7392a1e7a35a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I36ba87b69b5b9dd919319230f697dfad  <= 1'b0;
            Id5635595d6b7b6dd7e6d510a27ad6702        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id20e72ac258d1d1b6cdca1e6c9e3596d  <= 1'b0;
            Ice783314a4868f0bba8bc3c5e3b65ae4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifc34f5d6b7a7d0533439794958959856  <= 1'b0;
            Ib2d9b7f58cf571b904be02e6073f9b94        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I849ee5d34760be03d4285185136aa52e  <= 1'b0;
            I61b6effae91ae4bdcce4550eb5cf0796        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia3559d98eb372b7307f30ad1f7c4c7cd  <= 1'b0;
            If5cf6e81b0e3b77f6a45f2555201acc2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7332e088bbff69db19c62685e033d26a  <= 1'b0;
            I62fae5bf51588f28c3521715b834909d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I44daa5992b00e7af19adbee70bf01f2b  <= 1'b0;
            If5cbdab78a4cf86b6285a400d0e0ac90        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie517386cb5832e406fefc5e85eb2e7d1  <= 1'b0;
            I6e481cc49441c08bcd9fdcabbe90a000        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b096ce09467c10f448496fda13987d2  <= 1'b0;
            I3aa663be3dd604564ef68b9a2b9d7319        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If1c0a3726041f70e508d68cbf6e40e04  <= 1'b0;
            I8031632ee8700c63c207e2d6a6bdb630        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaf36ce8598a29573979c683a5e2cf9fd  <= 1'b0;
            If9be2701858da0bdffbf2dff7bcfd7e1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice82cfe55a5f226746e59e5c8beb46be  <= 1'b0;
            Ief209532f4cbf1c6a41bea414577f825        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iea1297491d1dfe98f395d8c73808a893  <= 1'b0;
            I1c8953ad3f64f3c3cc506808aad29dab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If43dd31198c8a0da6fabd194cf13bb70  <= 1'b0;
            I1b519d88bbf86cfb080a50ea0480a128        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibeb8c72b90b50c6897224ca1a792fa56  <= 1'b0;
            I5b8258f35d889071109216b464abb2a4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8e87530a131b5a73cad6df68b9e4967f  <= 1'b0;
            Id9681d4e0e4d375f9279de115a4337a3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idf8d15c7bd7705b9aafbda09c3a5b46c  <= 1'b0;
            Ib42144ece00b82debd70011724a29c91        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2aea17846a53e2eb2968581ee2c48226  <= 1'b0;
            Ic5717058a1815f63f164de1b1defe8cb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I169d8f2bb5fde5b202b4239b7a7f1ed5  <= 1'b0;
            Iea41672f012f225d64d9c75b198c812f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I40a223380fb4414a3f26a08cb90025ec  <= 1'b0;
            I3253481bee7dbfc0f3eac94c3252ee4e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7a070bd014e1d2c5e55e5fcba88a5664        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie117f6ec475f5d6444998af151ce4e69  <= 1'b0;
            I4a0a8b28429b708363458c74230b0fc2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If7f3174da35dd39af7f4792aaa649bf1  <= 1'b0;
            If585e4075ac1740f3b141ae6a50200f7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I719a892ad54e63b217c7271741b29cc5  <= 1'b0;
            Ie1a68cf09bb21a1629369fde87f51bea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4acf6d84471cd237f65c9b2391b7a20c  <= 1'b0;
            I72b8547125d0ad6c1ad39a68b55c818c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7a387a1f887c32e9d0f8e89912a8618c  <= 1'b0;
            Ie14ba4a8657740f9a8d057258db2cb09        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib862ac63c230ccde7fae0e62f9d047fe  <= 1'b0;
            I27490a69fb2a1f6f298639254c37cf9e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8f1a8a22637d37c3692e808d5eb3d543  <= 1'b0;
            I49b9c212fbe74a5dd8b087e417296186        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6f420c64640dfb0c001f57df7e3b4504  <= 1'b0;
            I0a8e6f5cc8b6ea599b7605abe6479bec        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3600031716c2b4e21c9f577d34e033dc  <= 1'b0;
            Ib6d94b34d3886717e4016fec196f277f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I002820a37fa7c6c504c487df4368e2cf  <= 1'b0;
            Id7e53d36da7171e036ebfc984dbcea6e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8a4c1f23212ff846400651b100add502  <= 1'b0;
            I2ec254d80fd0683d782302cf3839559b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice1ce5b4c30841dd92268559ebadafcf  <= 1'b0;
            Ibbedaef61051d5df82cd6d55e05c80da        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3eeeb1949945032d6c1759875426b733  <= 1'b0;
            I501336bb7ba172c05dd5840036e6228c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I384d5377ee6b8f7eb2db23a2e444ddbc  <= 1'b0;
            I8e5c4c6c63e42054359cee697cc0d026        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I30d615203b697787ead37394953925cc  <= 1'b0;
            Id3daa6db921871b752bf92366446afcc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib16548d471f0a4f4625852ea04335dcc  <= 1'b0;
            Id8367ec60787bfad0da8aa76c6ed8ddb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0987c561670b7b2b6683303c1be39561  <= 1'b0;
            I533649312ec995f1f9e514c59a8675b1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2bdf4736022e5da7294a0e851006a124  <= 1'b0;
            I0621d0b2c83e70b4afd65eb9dca4b514        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic6fd9592d2ffcb8f4ca83c6f0bd19975  <= 1'b0;
            I2ae01892a3cd0432618d7280b31daddb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I14bf11ad80890227e47fda26ae1b9c24  <= 1'b0;
            I5ed8a2f30bd2ea269341c2267ae3fe83        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8ca17b6cf35e1b1f8f601604575d3f27  <= 1'b0;
            I2c819e7f62c0dc0aac650074b203163b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I275cd09649a750edb8ae8313e4e1e279  <= 1'b0;
            Ia80693da8182ee2c3708b6ec21d397d2                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I30e20b58913d6fbe5817e1956ba8e570        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7d6a6026eb3c4d06e682523424f9628f  <= 1'b0;
            I1b922bed7f3c4a6705f3ce7a885a68cd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia0c192e590d8c914555b434ce5a634a8  <= 1'b0;
            I2f65f0917713ecc8585392d3b557c1bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic98c8641d2022080297c54ff2539e75d  <= 1'b0;
            I3301533e7d9e527118a67c462f1b4357        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I87f34821cd0b58f8855b25c75f2dd32d  <= 1'b0;
            I52a88bdb1f03da82730f7579b7b5305d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I87211ac14d832ad3205d47fb83cf256a  <= 1'b0;
            I644c730662b3725d26cd46fb46106104        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib81431cfb3b281555fa7e5b4582a2524  <= 1'b0;
            I3da3e36c76c4123bec6879bccb39e933        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I835b902949c2c4c09b757d4d35574a76  <= 1'b0;
            Iebde55cddc8170f7dd8855ea55eff0ce        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8510240df7dc41f85ad58a39868a1fd7  <= 1'b0;
            Ie673e2d92a7090b2fa1c5e14a2e03be3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1b6abc8fbab3849b285e9f88a4fe867b  <= 1'b0;
            If90afe75714f8660ad0eb9f9ea06cd6b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied638fee34f8baed4154b0b72e43a21e  <= 1'b0;
            Ifd96e3a6e0050c30a4308328cfecb21f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I14fa7aebb608d4a3d67176ba27d34d9a  <= 1'b0;
            I68b92cc2d83e9a718edd2aea82314016        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iad90879acba3fc2101829549264960f3  <= 1'b0;
            I6bdbb92363f0e072ed04654e9aad17a5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ife0952b85f14a960007b67646b0cd969  <= 1'b0;
            I87a4267db59b97ef1b9bca8743cb0322        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If876ca6a14ffb4323503ed46666bc25f  <= 1'b0;
            I44eacb2bea725efab7c0dd560279f0f8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2dfcbf493b761fb5d7c622e739b23f3  <= 1'b0;
            I87a2736466c5ee62b7cc55f17e715ffa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2c8f4a147b363d9c5ef0e080d9a9ed40  <= 1'b0;
            I7a66c7713ba126fdc24940cd92f7e10b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I485f9d1104a965d5d035feef912a2ca8  <= 1'b0;
            I1f11c579f34c41aade41c53f53468057        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I10fca5f2cbf5e2bc3433c0dda579a051  <= 1'b0;
            I651a438f70583d476ae10f066e035435        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If8572800d5d80cc92dd917b60447b63b  <= 1'b0;
            Ibdf17fa73794c846e15fe0a915b071e5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I24645082ef16129eed1c574f5fc601ca  <= 1'b0;
            I76d3221fbcefc0ee08655f7ba4919f3c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I207a0f6184a0b3be71766a8b47ea5535  <= 1'b0;
            I3458f69c90ea8b20b3d1f67e9a13ec2e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5cac08dabbb6de3b01c821d4db93a8e3  <= 1'b0;
            Ia2d6e9e1e92a30c7028af50ddfbb9bf9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe6b8c57d7ff47b6fdad5fadf1f6b841  <= 1'b0;
            I7fa3f2648baacebf9e4b59c179601fa6                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I66c91b5133d9812a03daecc0b14211f8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I477326720157df2503149125a43ee987  <= 1'b0;
            Ifb5986949e88167526d9fcfe07b417ca        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2c741a5fed7d88e9bdd6b7459feac649  <= 1'b0;
            Iedada801ca6cd173ee523ef335e91ff6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17a6511072c7fb4846be5844decf17d6  <= 1'b0;
            I4e2722e547586da7565b2d91a7fc91e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5ebc3047985651f4b9a957d502a97e95  <= 1'b0;
            Ib321a8ceda62c64ab25dc1c718301bda        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifa09fc1b009d073d5a9973b430c63469  <= 1'b0;
            I58daeebec4873e6c1c07c090ff81235c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie6212a29c7c6b035cfff4c869f945b68  <= 1'b0;
            I3f103fbbe49c86c9db46129bd4632cab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If343015b4815b01dae88bbb6f2017b3d  <= 1'b0;
            Id6697ca17f1bd6ddd112951b9d89a8ea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia0116a3cebf94318ed5b287960957ad6  <= 1'b0;
            I445ede2983c7470b4418a2ec0cbbd5e1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id75c23e80cdf25d883806ed20d4ae783  <= 1'b0;
            I034e56cd77ee400ed81b78177b202930        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1b43f29e0ddb72467befd6f3a9c1c829  <= 1'b0;
            I08edadbd9366786f96b44268d096b4aa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3fd0fa3b774d30a267d61e9427d09f3f  <= 1'b0;
            I8f86a7af86eb04c5df18e09888cdce7b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2eb08ebaa07a1004638cdd61a7209b7d  <= 1'b0;
            Ic00d037a11f8a27ab34e4daab8c9c2e6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I258c45897919cec5c6acaddee7f3a41b  <= 1'b0;
            I4d95ceccc6c3ad37f13c98339c59e5c4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib42d37576e3aff3d205f1f8822cc58b5  <= 1'b0;
            I1ea967d377f462a0e06d7d0d4d95b342        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c2ee281cd47a8414851c5e1c758ea65  <= 1'b0;
            Ib0feec63123e66bd6ad6935e9b7fa6bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie644d131c4f2c603e8e64c5581fdf822  <= 1'b0;
            I7d120060ddae9ff8f7206b3ef63eda50        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b76f0121a3f7e887e7121db50024ab4  <= 1'b0;
            Ib47f8f72386e2e65a88fbadd3a705225        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9eaf4e9ebe07717503ff69b51f0e1905  <= 1'b0;
            I4e0efc35346e2934f5bb4c34a4bc5f90        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icb0841ecf142687c3aa23e68f01c927c  <= 1'b0;
            I3ca1014802f58087e3434a1e0df19c01        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie8c0fac00a9de74870e59cbf9e87a39b  <= 1'b0;
            I688a3879b7be1544e6f94b4221c03213        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iae5d6faac1f5685cb1d400ee2b1d85e0  <= 1'b0;
            Ic22988138610c8671ec342f65f34c7ae        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib62b02ddf0f57bee49838d19783ef6c3  <= 1'b0;
            I0b85fdd83569e5cbb7d71eed50cb32fd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibd59d0e5a062f149bd0e91ba76985a13  <= 1'b0;
            Id7699f8f89380c315303644fdebacb32                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Idf55390c11e5b41ebc2a28e0af109913        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I876fdba97e755b74532f7ab191fbac14  <= 1'b0;
            I6b48935ea25672ee9a42f49eae9e519f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8edf1a08ef943f06ee28771c6e140e28  <= 1'b0;
            I6a9e6c39c20e45773dab7823a7ff9486        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7e12ad8a8ef857e02f4563b2f3a7f0ca  <= 1'b0;
            I42907182010c5889ddb7a700ead16525        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17b3a9df6752da6cc987e902e6bbad48  <= 1'b0;
            Ib6c26f3e3358cc2ed6fbda83eabd4bd3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I487496233a32f657171b3789590d0522  <= 1'b0;
            Ia50d85808790790450f87a5246874b3f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie34534dfd435b3d1cf35e82ca71e83ba  <= 1'b0;
            Id4a1744702d7808a80bc40697c864765        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0e8679271ba733bb87c44b6b9f0b6ed2  <= 1'b0;
            I0cf3d2f3e6793a2dcf15949da16ad28d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic14760b65c6fe150c3c48e64389a41d8  <= 1'b0;
            I90bd9107f4c931fa1ccb92998ea8cdeb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied6c684cdd280b41ffab93a026d27282  <= 1'b0;
            Ida1c729e6bfcec2c31a92aa9002f2c68        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id0f4dbb72da33748d8baf723c5a32567  <= 1'b0;
            Ib848feeccd0ea78ebc8ba8368534c3d1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib0bb71b1f8829347b3a9a7543f9dd964  <= 1'b0;
            Icc11970bbae3adcfa33a0e5dba3e78f4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I47cbb92d2284aef7b9e56e88f0ba6f7e  <= 1'b0;
            I86bb4ef4bdd7af8861280ef30fbeeeea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic69094123b75ae36e3e54f179a9f2cb5  <= 1'b0;
            I7e0c259c6c7bacdff5edc44a22e005ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I07abbbd75d91018ac53f53e64cffafb9  <= 1'b0;
            I897ddba059b27f7ed009b0cb70cfb46f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib02268d5048c7c8e83118070e927453f  <= 1'b0;
            I4496243eb0542a514b551b4d09bffd7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc2a9c6dd8d2aa912548c918c8a488f4  <= 1'b0;
            Ic931fb08b2e8441321ebdeed84576a0d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5ad7eb9d3ce7c712515254f892d1670d  <= 1'b0;
            Ieb6af5390b98e893ee05a939c16d2ffd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ife25829fb3c5023b7d69bbaadf9cf77e  <= 1'b0;
            Ic2a54bad4c5a8885dd24b8687c6db0de        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8b2a79aa4ac88e6b4ca8188a7852022e  <= 1'b0;
            I6ecbad763d2b48b78a0584beaefc78ee        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I081e2595b18f306a74d070203447ecf6  <= 1'b0;
            I20556d23c873c71c7ebc8a961bf40251        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I68b152a599887c0039dd9d45c528c219  <= 1'b0;
            I79012e6351e6320c22437aa216ea4df1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id051f1d5454802e0eb37e22248efe8ca  <= 1'b0;
            Ibf74ab9af877d27c3a6f3881f00ddaf1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic4c6f707f461cebbc4c93f2ba664ae7b  <= 1'b0;
            Ibf3e1ead3776901898d4b154aeb61267                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I843d35db35d7b42a87ce78d3772cec2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia538dadbd6ae3711740595a18c89b65d  <= 1'b0;
            I2b1398b4bfd374d7221b0a68da28e979        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie7d9730b191781c78391141d95d4f8bd  <= 1'b0;
            I6f615d6e74b0c02f8e4265523ad16404        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I12f2f886517647044cc251861721bbb9  <= 1'b0;
            Iae8a98dd4a7cbfbc56c1404b6a2020af        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I615053b36a1851a06125e2ed5ec7f880  <= 1'b0;
            Iad53375a54d01c559c74981bf279dfb5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifbc6aa14cd448bbe416897a3671ba857  <= 1'b0;
            I5db1307f922e0c742d7d9f3a79a4a4f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie596289582a73e37f78f4ca4cab21e3c  <= 1'b0;
            I9f78172ed5bf73752196f9a8810005f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifad8c7bacf72583f91be27fbe5b7a1e1  <= 1'b0;
            If85a22d670d47f491dd7568d0453ba1d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie74c72742807ae4243748fd27d80d626  <= 1'b0;
            Ib9e529170b2896e930a839295796fd31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie7a68c2b368a295f95571bc4a109b9f1  <= 1'b0;
            Ib7af536846bac40c1f221d1f72c6c25c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id88a7edf897eea1b4a137141789a04f5  <= 1'b0;
            Ib0eb61a2cb831dd35ce9850994e7c2da        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib13436ad16a37d656d6b1ee95b9aee20  <= 1'b0;
            I89d338f59960af7a47595d6afa206abc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc07dc30c0a957e474546ac7a60df38f  <= 1'b0;
            Ib3c1176eb8991e3e85855a9fe845c303        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I595665d8128bb87ab62741d7ac520a4b  <= 1'b0;
            I93073d05d509b821a743998cf32c58ee        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I256050251d23250854ff337bef28e460  <= 1'b0;
            Iab6dac1909c1564c3890ffecc13418df        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I82f0e5a32d1bcd761a74f1f9ce8c88ba  <= 1'b0;
            I1b75eeb29167a171d89f6e67039436d5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I98febac90cccb5fc1f3d966b6e38c4d3  <= 1'b0;
            I3a31adc52a1405555017b2ddf219b407        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib534288c2cf976b6ec85db743bc2a823  <= 1'b0;
            Iaadba89c6a370240fc0758029f7d8db0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If988b82b86db1f4ff6d3695f7b0197e4  <= 1'b0;
            I4f4a64fb3ced7d9f7ee4513178e9655a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6ef260ef75e47b011a46ba2080ac3684  <= 1'b0;
            I0c76ca58f69c91758e755cd581241284        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifc1da524e7670772834d521a6fc4c96f  <= 1'b0;
            I2312bce18958346149c868846e04643b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I852d5295a32984af00c95f6d9389555e  <= 1'b0;
            I3e154098cb0a48f1c23234f46613f406        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3c0a621dbef864fd1f566bc2e47f32c6  <= 1'b0;
            I1645c1c588bcbf15dd62d47e08b8e139        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic04828ba2db8239b093043c27476d345  <= 1'b0;
            Ie486617fc1d6354c7f347692cdbd894d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4c25de66590e1745d37112e08d8c8e2c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I319012bc6fe93d78de57bcace0caaef5  <= 1'b0;
            Ia03092ac621b8dd1c206fea1e8b0215f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibb35bace971548c9fc98d773d1aff712  <= 1'b0;
            I5c9bdb033436dc9f6069baca31f24c2d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I90023493600924a76d2192080cf6194e  <= 1'b0;
            I8f07cf4865480f18ad6945974ec2231c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia9f5ce4603af279bbd9b486b67016482  <= 1'b0;
            I4a7119e8862fe4a6a4100dd9ac67dd24        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I05721e06a1acdcc0571907c7d853f18c  <= 1'b0;
            Id78fcfc6724a05f46d44d7c3e7d0c756        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibfcfd3151af0d82bfce293ada44059b3  <= 1'b0;
            I7cbd9d619623cbabf8ed6b1fece8f012        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9539fcc40d26b13015a864718b116d5b  <= 1'b0;
            I58951165d251e370b0f3b3fb537aed18        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5490039998187a1a2efc3549e3dee7d6  <= 1'b0;
            I21daac106f526d84cb8fa5239c19499d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2b97a79c90f6578c8b2f321f8d598cc8  <= 1'b0;
            I178029cec3a5d6141abdfa91b91fdbf4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0c616f736879c28a5222de3d6f49a587  <= 1'b0;
            I7ba403c6745e7d026282ad704e065702                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I96dfb2efbb55a644616e3474ed07c364        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5590d801fd7fb496019d4c31b7c6d898  <= 1'b0;
            I7a17d8f0e2d16c441044db68ee037731        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I27e1d2e0e980216b27b90ea48c061025  <= 1'b0;
            I2ced9bb3ae6bdc5b5ef2865fb46abf07        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I474f6bd977f4197742d0bddb3bece684  <= 1'b0;
            I89a93384020d93cf4d26b3902e06cd9e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaa1e981134f5a5c02983c49562683bc5  <= 1'b0;
            Ibbb47d29b9a45559c13ffa3b046c66f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib051eb1091a85f85a1e50007f1b27cab  <= 1'b0;
            I0034177eb1049577a3578b371527f34b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6b5645cdde4b35a16fe3e91d90caaa4e  <= 1'b0;
            I22d9ea7bb5a1a3405bcd04b9af40fa62        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8850ab26807dcd55fefadf6310729ca7  <= 1'b0;
            I8a632e7a911bf5726fee587189cb6f16        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic5cb81c821716a8aabf8cc2283ff73ba  <= 1'b0;
            I3765afc490b34e8a310998a4ebcff8cb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9a6923c6368526a53ef70e16471386ef  <= 1'b0;
            I7607e800ae46a96e016b303120da4247        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I620b8ecdcaccc1ec80ebcf9fa6af0017  <= 1'b0;
            I93cb3974b8594665b2e7ce5593fde69b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I29b2f1fddee5e32f217d25410bcfce4f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I141cda06bae0c5666e3bc61c6fe5ad66  <= 1'b0;
            Iba5f8a31a81f6aa06f5e38c03dc6db54        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia9c273b32d0701c7f185ab2de9e57829  <= 1'b0;
            Ifcb5c907ad503331317599e4e0ce7be8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic3fb524ab434e80b3289c9241b65d224  <= 1'b0;
            I62d6f2ab4ec8b6ecfa544ad4d90eb30b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I23c8b64e433af0bd00cef44e38df99f8  <= 1'b0;
            Ide65414c51b3cb182c0f2f238903d60a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If6a5dc79c0f6ce348956286737a369d8  <= 1'b0;
            I03a8dc2288eaeb619e746990e20cc868        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I34e6e9d2153e4a70ee36ab85e72d5318  <= 1'b0;
            Id81c1b44d16ddbcd466382c60fe84986        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifdabf743a8cb46b7053000ff48ea0c60  <= 1'b0;
            I503d72f4a2fd20dbf35aa27321d2ede7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I22f5bb821a2571d1764978fd76c8f1d0  <= 1'b0;
            Id6595a4cf33062d1f05cbcee2d0685f1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1b695aa715615662eff7065c742b0859  <= 1'b0;
            I83ebdd7331ca8fbcf5250851b346c0b0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iec91b3ca3b54010755d57f8b8ea4a544  <= 1'b0;
            Id6a9ab06d58c3a01e1fe04fcf61406fd                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7f6ea26cdfe5986065e7b5aa6842cc1c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I06ad520cb02e46d34c45f207d42a9243  <= 1'b0;
            Idab1ec32c20f93c4cc1acb38158f92d5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9d18ff3465afd8cae63abba68487542e  <= 1'b0;
            I0738add83419502e73674ded2f1ad6c7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I914dedc1d5e5e21c9b8d07ec0ecc01f9  <= 1'b0;
            I6c93e63a8e5a2dbd598f1565c7323b39        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3375fff5ee0d4b4b12c5a70fbdee59fe  <= 1'b0;
            I4aa57a9d46371f1680d5f95596f60b5d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia8e304ca12c82e41cb8e4de7be199394  <= 1'b0;
            I5369a7203b78951a3c006c2d3b22507c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3566f2779e860008b1a5d305366a07c9  <= 1'b0;
            Ie72a79a6966cf198687b7c8a8bcdeb13        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie68b31360c12a83c6095254b6f14603c  <= 1'b0;
            Ie917ae4c44ab0f9c2f1747ff0d2a754e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I42ae0c42360c977b35429ce290516a6f  <= 1'b0;
            I0b1a31ccb34a742552c11b1945e23dd8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe01835305315fab50269c72ef849b61  <= 1'b0;
            I9a65a845cf2eced39050e8481665f557        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id806a2df1c4519bbbe811791cb4072f9  <= 1'b0;
            I261bd53528b82128acabd405389c8d60                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3b402b35d38a9fde312c89b82297c1a5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifb70a30f8bade95f402e71f95fe6644b  <= 1'b0;
            I309fa33562370e339c19e2377e6a6a7a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I592a495aecc800236c3470ff8e6adbb5  <= 1'b0;
            I7d06aed81222a030837cad2074c68e19        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c8024aa9d81704d2dcf63e34853f8cf  <= 1'b0;
            I835cc6af0cd8189035f2441c2e0d3100        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ief03713f5cf37200373a20d42c7fc9eb  <= 1'b0;
            If6f768d12f04087246a0d65de1aef99b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic3cb34aae74c5f1a870b3635f8a40764  <= 1'b0;
            If7fa833bf1b1438e7a5bc783ee745252                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie4b180e1e2cadb865b0eaf6509f99dbb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifa3df8b249467cc1e827c69925ef415f  <= 1'b0;
            Ie329a11fc3f6f59f6f1790612fde3250        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icf3ad912aaeaa0c5cd1ab0edb898d6e8  <= 1'b0;
            Idb7ddbee4076f7bf49177e69f5e4d112        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib774f380e3d7cfd1f5f064e93d8134b4  <= 1'b0;
            I614d66a7dca2d08efdfdc157ca803d5c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic07c650e6e49892a41cfaf3a37471426  <= 1'b0;
            Iea16eb0ab70ebb1bc47ae55e11ced62d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib1073489d63ea33d7f3892f4ff875358  <= 1'b0;
            Ibb103853fc21f8f3d466ca16557ccd3e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ifa8db43284d5bbebaed4f72d65cf9f92        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I174b6c36f2af82f8047cc76543a3b4ee  <= 1'b0;
            I365d9f3e8b2a9890427f07386deeb093        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I953b975a89adcc88039284970e9b3404  <= 1'b0;
            I466aaa0b6cde2ade1901797b8c11e32c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2b40d249c531e10cc22d1335f350441  <= 1'b0;
            I7057e329a65ab240ed6cfa824307af65        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I44ccc3ae897109dd51f9afeef93daca4  <= 1'b0;
            I624e50e3457d33d12680eaf8e7c34aa3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie9236599cea94cfb603c6b977fdbb44a  <= 1'b0;
            I37446eb66ccfd268cb418655b8160fe1                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9f356fd6820c33fdb5baff05a781e192        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I25f1ee9cee4d04bd8fec1fe601d016d7  <= 1'b0;
            I39b9c7c664fe7017731877d145d55b44        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5ec1e530b9007a75a778af4d82ab427b  <= 1'b0;
            Ic62ffbb9e58e0d08b0dec24bba1dc6f2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8a9e516aa824260998d10db758642bb0  <= 1'b0;
            I8da2a532288fb817e7dc0cb7b4e3761c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I70dd1350d65155ee7b562f4c79024a3d  <= 1'b0;
            I6a6e559f5c98f846014e8107fea5a5d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic9146d8b3dd0c612073b70b8a8791e8c  <= 1'b0;
            Id17f6250f8c7f1d7f75fd27f92698da3                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ibef9219f577b1a62dfdd77296fbfb24d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I857d3155df0b6dd704514b039c66fa97  <= 1'b0;
            I52e6688b5bfff75529d18e20b22832ce        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc1b8aa2f81a7fbd87e4f5821d14bf01  <= 1'b0;
            Iff22c49354eefca0ea3c5959c14b782c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I68b585571699a57bc6ba5e8955467119  <= 1'b0;
            Ie5377bbdb4111ed00356d5b7737102f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib70e99c3acc76286a6811bcacc9284de  <= 1'b0;
            I55bf0f3379a8c44634b8f0a3d06c049e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iee17ece482d04964d3c21a092ec955a4  <= 1'b0;
            I9957b02e8d0d888e6950eb553d9084d7                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9bc9541607f4f6aedb686cdde297bcda        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5a247475beb737d470f03507e55f5b24  <= 1'b0;
            Ia4620554fbb1d81a71a15a846e4be2f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I13b0c9578f7b6b3b7e6704d7b44079c4  <= 1'b0;
            Ibb31b35388ba8ba2ecf98449308ee67d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I41eff06fe1dea8be4613945de596d3ca  <= 1'b0;
            Ia20410fb3d56587f89a54c00b943b305        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I08f22261d5713c0636d77c7938f592d6  <= 1'b0;
            I9d268f3da12e35b9a4229b7340c0f018        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c7e41b9cb1bdb6f649c88c0ed3f4100  <= 1'b0;
            Ic71258b745437bc8463fb4f847c55e27                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2fce29bd666082eedb2fb3ec8b5ae4dd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idd59a5357d4c835379ed180ac0924bf1  <= 1'b0;
            Ia1e8b61e2579a90f5c88ded11c7322c2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe7e5c2cb9c50eca34a3859d13e83a92  <= 1'b0;
            I8cf3718ba65b7fed72e3955f190e34d1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibf5c141c5cc0a6a20c05b52bf8282476  <= 1'b0;
            I7e802d300af54d394b4ee041798c0513        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0038305f94aaefe2cd1a243580d95932  <= 1'b0;
            Id4fd5a4b97cfa1e176a26f3a823c5516        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5364deb983adc2ae505ed2b8c57f876d  <= 1'b0;
            I24bb5c315eacf0f4e8c86f6582389e39                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icbf8d4e75fc66c05eb49c5075696fb07        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifdb5589982db805a0416e1c01276249a  <= 1'b0;
            I746a7e90adb2f213b75ae12a161aca0d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8bb5522183b65583fda83067990b3e94  <= 1'b0;
            Icb1029aaaaed8c698862ea9c5e22132c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1e77fe6aeaba852aba34ed37dd53add6  <= 1'b0;
            Ib93ea7028c172373b53cdafecae32a67        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9171019227f35760d02d0c8ce786f4d3  <= 1'b0;
            If9628275b000e418f3903daebfdace92        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6e92a48aaab94074a555efa9bd1e7243  <= 1'b0;
            I607f203694ff76930cfee4103cb73c30                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I830202fb6f08f98c7f71893a881bd555        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3bc094d67805664859fdcb66f1360e64  <= 1'b0;
            I6f38bc9359562f57c1603355e9ee312b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2518ccf385b3b677d95983bc550282e8  <= 1'b0;
            I4701b732d59c26e3790a63c1936f9a24        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7547c56b32513ad45d775b4502596d9d  <= 1'b0;
            Ib5d28d8f73d17ab6df6a1291e50c04ab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I013d84bfd582acc7accf07ec522961fa  <= 1'b0;
            I81259f391db792339824ad5dd1a0057b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0ec27b590ee6dcdd9c1086105e3b6c23  <= 1'b0;
            I6f09ac63effe67a86798b9b4e1690664        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4cdc955fa9afc75c2c977de4ec540e1e  <= 1'b0;
            I370b4b3a0048a93ba374a40e170c75a3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ieefbb5d6f4ac1e586832c5c0f513c5a2  <= 1'b0;
            I3f8476d0aa0ea2439b67ea1a4adf36c5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic828cdd5dfde844df4c150921af2a443  <= 1'b0;
            I35b52dba10a8a5b22b518388fecac82d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idf1ecab26889c4adcb835fda6b1cb368  <= 1'b0;
            Ic7db274ed18e6fdecf30381a31238777        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I00d3f14b20e1ea7d726533386e0eba27  <= 1'b0;
            I2c4e538a8db759e9799541d9178ec61e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7f720a18542528f0c9bfb14f699ff4da  <= 1'b0;
            Ief6d4c3f5ef8663e111ef99347b023f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia98a6f01e4eb5bc74d50d350e79be426  <= 1'b0;
            Id95e964e5faecb52c72669b0d28a4bf5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I182b43872d50de6f7afb700f178b160e  <= 1'b0;
            I0fcef4538102ac6d24aa7090d5405afa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic9b72b2a91d951cf08cf54ed215ecaa8  <= 1'b0;
            Ica8e4c56ebb37e189ca8e6b3daafdb80                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I055019e38eec6badd1739033d43d7d97        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I93084ccf5b5e4efaee968b497bb2a775  <= 1'b0;
            I35c20a6e823da77a870b421eef2e0a95        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id38852415486e6989b89a0d85ad6771b  <= 1'b0;
            I32cc12cdacef1a4ef64577e0fa977f46        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17cf58ef5326978c62c03c56090a299f  <= 1'b0;
            I26b3f2360ca4a8caee61b2f3a3a08267        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie41ca18c7d11a47e274f9c33f75393ec  <= 1'b0;
            I5ef9b7dc0c63e9ca6a5fb5f7ffa06041        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7b80b4902fe98c10dd72c9eb082346e5  <= 1'b0;
            If881473b05090f40a027d7eeee7f7ed9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I20ffba20af04b99954bf719589e90d1a  <= 1'b0;
            I23bd59ab5b038935301396aaf2acefc1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If8fe5af7e5c3c97b5a713f6bcf919f1f  <= 1'b0;
            I874386d94dacf84e699d159af1a49836        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc5fb0f3a04ab32948e249e088a11b11  <= 1'b0;
            I95bfe51a759bf4165168e5e3b99d6b34        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia9f1e580e8f441394d719d52a7bad688  <= 1'b0;
            I4ba5b2f9b7ec0937ecd2c9945cf6de87        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I02849282dd1bd663fd39baccf41762f9  <= 1'b0;
            I0b08fb8db0e8a1de3d416907c87fe700        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie4cda4648f6ceb76b8fb74f290ab6439  <= 1'b0;
            Ie030d12e5acf9ef4975a17c83b2481c1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I24135210c23b2422a42c90ee25594191  <= 1'b0;
            Ia7a0e852d3dfcef950804ea0ebb0c80a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib08897f9216599042f7b97b137e07fe1  <= 1'b0;
            Iaa4c38d030eab2b7899399aa0d7886d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I51e14ece9ab6607f83e6ba27f3f046a9  <= 1'b0;
            I7089386c94261e0febf3b4f7dc1aec30                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icce7ff1d652d4d9c2be5ecf679059bbe        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7a626ec321bf963a5401892a7e3891c7  <= 1'b0;
            If816bc5eacaea23443602e575ddf60b8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If76f04fe0baf171d7df2c0cd849aea2b  <= 1'b0;
            I3b224a4ded05446cc5300d430bdd1947        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia9c8cc5e3becf3d48feedec8fa2c93a4  <= 1'b0;
            Ia5fc5cfb0e52237b407b37a3858fccb5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If3b77c41fabcdb283f2c6fdacaa5e9a4  <= 1'b0;
            I92f8ba6e7f8e9b30fb5b6973eb8fd03e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie5373b01a92f2ff85be8077cfef2175a  <= 1'b0;
            Icdfa60d2a024dd934f7e6639c6cb2c28        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5109afc4dc91780e05704ea5e1399e3e  <= 1'b0;
            Ifff70b976513eaa42b6bd4b80c98611e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3e0b41bee4c76eb5f3340ad23bfa01ad  <= 1'b0;
            Ica12fa8b631b70a6bbe9f6e92bf73ea0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic0732810fd355d59a3168be896a0f9ac  <= 1'b0;
            Ie69c255335760f706c644b115887269b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I220e32641265b46527ca61111f7ebf1b  <= 1'b0;
            Idb06676b41de19bc86eae34c292183d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice59d2af73d0b0f2ae91a2ef0c2b7f04  <= 1'b0;
            Ib21d2306d5ded3406fac754e69a10d20        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic308610ea8bb62ecb6094192e02dbdba  <= 1'b0;
            Ib41d1aa2dcf81879976fb8964cbf6f79        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I33ee415d85e2bcd8f975d34b880f6ea7  <= 1'b0;
            I5f8f5e246f008b8d8c75f72828337bab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie61f299252b8fecfd3e8634b64df5a90  <= 1'b0;
            Id6625e78da0e14d2eeb19cc8ac6520e0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icc67656ad2dd3fffae4e5abe02f8fff9  <= 1'b0;
            Ia1e4f20f32f7371cb0078d6e80fe8b7e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6d9ddc6afa559ac35c042df1a9390ce9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0c47ccef4b55410286248884a7249703  <= 1'b0;
            I9334055c7833676469670372d3c5cc31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I94e4041b482064334fd0ed92b91bde89  <= 1'b0;
            I0c97d772c737c6ff85b584bf69ccaf93        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I39d3bce4060032a81e6b6a1c1805cfe8  <= 1'b0;
            Ic6ce97ae85d91dd8a79f3f9d0da375a2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifb422c30663eb4824caa72326b238df6  <= 1'b0;
            I83ff9a2750b298b0f7c9b6ce13f574af        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I41ab6fb6ec6ef7ffff70e50f25f217b6  <= 1'b0;
            I85699a2a05c343a6a9e828af6d445e9e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ce10718a2211184999663c3c2493cc1  <= 1'b0;
            I51f6e39b24b2554884e381be79f47ff2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I877e8d94236c3d8b0a31858a98fba5d6  <= 1'b0;
            I9f65fd05c6929300860c8cbbde5607f2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iff2f1716cbd73b406d8f07c22dc79fc8  <= 1'b0;
            If09761d8f06051d4287ee29ac9c9fa19        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibc48fabc172f27ebce18d0a9b5120dc5  <= 1'b0;
            I33bfbe0bcca6d32c86b9576577e3f265        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie562ebb336e476a81f20a652d4cb20f1  <= 1'b0;
            If2921210b1c05ecbf00af3a2bcb96ef4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib5ee5a6ffc45ed1fece0822dc4619b57  <= 1'b0;
            Ib074e38e280474a782da831a3e0028b4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I86ba73ee348f80e2f9891d2ebc8a02ed  <= 1'b0;
            I507449dde0bc0c8f53a10759436ec731        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1e96d5af3d0e3fdce39530dfd0131a7d  <= 1'b0;
            Id55a3e3f2d75baeba71a345fad695c69        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I38352b363fa37f6f822fbc1a39100968  <= 1'b0;
            I790cbca796af58b1726d0a4680cc164f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I20984f43d22671639a7a178ad15aec04        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4ba41864bb1d2130c6971e0b2903027a  <= 1'b0;
            I59f88336d6bdd50ded87d353fb5ce3e9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib68deeb7bec4ca3585d1a4dcbf8793f1  <= 1'b0;
            I488635e3f7ed77ea88199f5bffd4b1d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ida3d808d100e0bba290f96ed9e744e65  <= 1'b0;
            Ie6893017d21c050ba10d206854f4a9f4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4d4901ff372f6820ca9c8c29cefa664a  <= 1'b0;
            Id3f68b4dc0ab60673208b7d2081f3533        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib99e1b93fb7fbda260d93eea3d24c3e9  <= 1'b0;
            I433756b944e061a824a89bda241e879f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I019e399a1cef87745e025a7d74e94db0  <= 1'b0;
            I2eb60a922aa4f7482dd92b9351d53a2d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia8974083bfd064f2c27dcd421490fcfd  <= 1'b0;
            I0a93f095f9efb1542116a295c0db9c8b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0867979e1b159c8ceae548930376f482        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8fd5787ebf758919e7cb75d7419441e8  <= 1'b0;
            I4accfbeae8a5ee0dbeab23ef3a116145        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id14074d5230885c38b89b09b130ecf68  <= 1'b0;
            Ic7570b0b7c5bef5758f68562ae4c90f6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I86fefad34d3c864dd0e725133f303b4f  <= 1'b0;
            Iceadadc4456881fdeea85934a9bf4d6c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1ca188bcdebbf41d84f7a5220bd1d195  <= 1'b0;
            I7b2b617ae67424f54961eebce42de77e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifc640243288c9b37b7eb9e00351b23f0  <= 1'b0;
            I953f0f8af76f89b2d9ab4abf19fb411d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3d149293f106ae8680c7f4702daa0bd6  <= 1'b0;
            I915b4736dcb20f831d02e48f4e79f008        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie232799bd6c4ec99e24c78f3ad798265  <= 1'b0;
            I989ba39f188a44475a83e65a4960d2af                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ib7eec587348ae1ca1f00c0a3ad10ad27        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifebcf64858d5e2d07ad7894d6182eb11  <= 1'b0;
            I001a212686304248c8359e5fc01227c0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibab55499323660588ec82ebd07ab0572  <= 1'b0;
            Ibb7554e012c0fc1223c29b759c900666        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I89af7644c48a80d7d22f50b008d35841  <= 1'b0;
            I9aeb9c42b54a05be6bf9b7b88b6860ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0152dc6e6a7acd72a2144623e63998ef  <= 1'b0;
            I6a5a5966965b0790b906c6fda71aef80        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I951dedd7af44c3865a8f36888432d0c9  <= 1'b0;
            Ic943083ca65ace6c42d73f4234739a06        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8188dd7cb03854c6f709de06ff785d91  <= 1'b0;
            Id0b321686d4c39621024cf0dd99822dc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3b30b4ab00a49e10a75587aa324d6132  <= 1'b0;
            I9bcc1d9b3dd258fa7b6042f0185d48cb                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0839dd3787442f1b79b87e02436bfdce        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie50aca688b3433fad7565998cb900155  <= 1'b0;
            I89e6a9fd97d8aa4dd3b832c3be4697b2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3342fe0c5d3ee5021892d53eb45bde21  <= 1'b0;
            I93d4157f48b132642752220059861e98        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5134b762ac428bed07ce102d8927a418  <= 1'b0;
            I8fc4faa2891d7fd3479ac1f788f481dc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic14f948884da19a272a4760ffaab9ea9  <= 1'b0;
            I440f30e9cb4bc89233b46ea00b4cbeb4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I46e1047bca2b38e62b4de80d1d2249de  <= 1'b0;
            I6568bfd8780c11e0b1b049a01f92abd8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I866b30a63b3b5fb708934a1cbb0e1d9a  <= 1'b0;
            Ibf7dc4da07f9955d5d4c7e1f63f1ad68        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaddc1f2e822fd2fe9d9046d759a82cb4  <= 1'b0;
            I9ba14715d9f33ef45681ad52f5be9593                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7ec1a328587b72a39c462083efea0ee0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If9285bf7611bcc5ea6432215c349e021  <= 1'b0;
            Iaf028e7ab4dc77a7649f15d603834b5f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id277f5f05551eeb5dec1701056330da1  <= 1'b0;
            I58db79a8e9f0cd1ded379897ba2f27ae        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9963d0b24763ed8038b1f3922b8f9548  <= 1'b0;
            I6d3cb4ccb4e51c7e6603d0abd1a082c4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia98de3691917dfb63bebdc3f8655c8be  <= 1'b0;
            I79f75f49ea8a29d684af396014b2f3ab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0bce960fcc58938e6a1e01b912eabbf2  <= 1'b0;
            I9c5ecd86bedb189fada40fae9d751a68        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice5f7168aeb940d48093cc9df7cba36b  <= 1'b0;
            Iad5f06e1989ead7d306c70a3b02cb8f4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I859d795a7d141eb777c1f3c038203794  <= 1'b0;
            If6d1a410df5a4aea6a01337a6074fbd9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0dccb8eaad52ce4d780696a8485420f1  <= 1'b0;
            I3bc40a4db14566b5099b14cee5f61135        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6d4fc81ced37c159303c243af04d345e  <= 1'b0;
            I7e683fd8235d7cfbf4ff407a286f07de        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iefdb8bd28839af9413a3906cbfe715e6  <= 1'b0;
            I97afcedf05e588b7976d6005191dc916        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0615acb0f7cf79b5f6ae8e91cb525dc9  <= 1'b0;
            Ib8d8eec0aaa662adf2837c9b705fce7e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ieed4c810a5bb69de112522dcf00b16ed  <= 1'b0;
            Icbd765be950123705955e2c5d7ace84b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If533578cacb685a95afbb8e1c05d3c07  <= 1'b0;
            I396a897f79b519f4fa02af39d0274f64                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I706e8f5617cfae1e6fc83db18c8b5fe3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia858ff5551286beffd4cf82f876d30ac  <= 1'b0;
            I1dd8f8c7f1b673898096b1f3ae383197        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4c66570630a650fa7b9bec543f685487  <= 1'b0;
            I10ca8978cf4659265ed25a27d09acc1c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If10f33385e236eaba56cbab8c2883399  <= 1'b0;
            Iec4656b32460def4a608b6b0f6486af9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7cb58e4c486e683faa4acad4756815d5  <= 1'b0;
            I5f4475897d1d58965da1b35fe0ef8c01        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I452e51cca9acec44e36e4efd21b43034  <= 1'b0;
            Ife61469306df3cf220666b187f1496a9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ice0234f25de4ab1f03a3cb01a2d61dbf  <= 1'b0;
            Ib49319b9dfa4914f92f423ceaf840014        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I12a18a1f8d4416e9bc8abee6ac3dacfc  <= 1'b0;
            I93ff2f879233cac9b9f0dd2f4c082c09        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id17ada8dae3f9810d1892d34f2288859  <= 1'b0;
            I44597d694e9c5d29280e503d72a27c8d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia2c5fe53cb5b318fa63d09881609655f  <= 1'b0;
            I04a19448c5e75af8021ad02d1a708bb0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I579c7926e7b78f4ffc606adc10522f53  <= 1'b0;
            I71a3093121c2f19dcd1412b468652fa8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iffa06a336949f56f4e5a88a06d8b7e60  <= 1'b0;
            I3ae09c82029c617034fe6aacbe9e94e6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaf82668eb49248709540f2f529f1b3e4  <= 1'b0;
            Ie7af6b3b441f910b000a333afad6c76f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I90b3708abdf742370f06cc513ee307e1  <= 1'b0;
            I197c0cd576e16ee2197a28c86397f801                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4d71dfea8407aa5b5cbb991bc4fea963        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia17906696bd0e095d7a5297da2e049ea  <= 1'b0;
            I1a082caecc831a90e74674ba35da4183        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I180d4f3b23b518271d7cb8189fbeadc5  <= 1'b0;
            Iec1de44616a2354a56ab1f681059d4c5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id79636d195efff260c430978f0bcee9c  <= 1'b0;
            Ie3c2318e64d0e218c3db557404c4aac8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idbf4ad11ab2a27044193448c8739fec6  <= 1'b0;
            I9a251d50f41e51b1a5cc2475f267e8a0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3051f561a5e1131ebf167cb6ccb5adf4  <= 1'b0;
            I9b5767a49f7b9dcb8fdaea924835033c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9322a2a61900943075bbc23c72a3f65d  <= 1'b0;
            I6ca1e6700a19d03621a193c7240bff54        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iedc463e359dd3003d9f7e50f3e858e93  <= 1'b0;
            I931c597ff12bffce581f653346202f83        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie7cfdd25541414ff3f8d6e5d7677fbe5  <= 1'b0;
            Ia3a2c5d59f6340917ca3933c05ba4678        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1e93f0470d2818249f1c28ef2a399a0e  <= 1'b0;
            Ie83d0a8ee5ed214bc7577467748aaa04        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5d6e576b0fa7e3219aaf9ccc345085b8  <= 1'b0;
            Iaac29552e5fc65aaf4f0116f917b707c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id962beade26396738ba0e97f67d5e261  <= 1'b0;
            Ie2c8eac7204b98139c03b6fbfff9af36        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id0ab747d92288f23cef793567b2363d1  <= 1'b0;
            Ied7fcdaec662cb3c2f89f131986fa102        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie536879e6fa9be65376d7f00e0fc40d0  <= 1'b0;
            I094a178e55425f27ac1ff6195217396b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ib16a17d6430570b45a304d847ee2b11c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibf312ae4f51fbc44b43848f9df62a45f  <= 1'b0;
            I42169e454756fe4d1c5f17f2eeb2e091        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icfc03646b36b971b9fa57d04a26dbfc4  <= 1'b0;
            I6fde38a3a92e06fa77123e3279813c41        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4f134c0669b5a6a8c7e03be7eee30c6c  <= 1'b0;
            Id8ee16437e8d6d6da6d37440e04097b6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6c765e677f42fe600b848698c8a78349  <= 1'b0;
            Ibf249d8e5acced9b064132575f40e001        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I284b23051c85300c2a1e3afe8f25e99e  <= 1'b0;
            I580659084e3d17b48de6b1c66154fcf5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b560d9baf8a7422b0dd84720e924ced  <= 1'b0;
            I7a14e45d43ab77b265501902152c8616        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I457ae11ad90c8478751eb4b42764e158  <= 1'b0;
            I81ba868784103e0eb05a44d981d4d666        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2b7822d5d77aaed61eee87570564df76  <= 1'b0;
            Ic6b88783957cbaf253648a30b22f6b1c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibdad0ab78e4404c852e60a2b04c3a5f6  <= 1'b0;
            I4103c218a85a1d08db5c4f4b5686b2e5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic4efba3932e598784f5b9ad6ad04772d  <= 1'b0;
            I0e6c0958af503e4a120a49d02a432863        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia03836a4e93d2f36513227d1dfaea0fa  <= 1'b0;
            I8f76b31e8f15c0e5fe24dcb723418111        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I138fb0c48f2d27e3315e237d9e61d653  <= 1'b0;
            Id1457221b58344b60070aa026436df2c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id0b1c46fa4caa63a4c63a44ba3c5ef8a  <= 1'b0;
            I3177408f7d08b431be99297fb10586e6                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icc31966508e03d8869e81d8aeb243705        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3566033cf5c9a06977c9182925750707  <= 1'b0;
            I9dcccf542ba434b6e0fde6f012f98f92        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I02812a8a833bb69eb168a1004b6fafdf  <= 1'b0;
            I51ccbb824a5e1e340eefd173c4491728        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie886c5effc85f1fe0b6411db4a2cde77  <= 1'b0;
            Ib7ae1730dcd8bc708bbfcc6a9f97ac66        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibab1d13cd6a4f7b0c79c9f845339e53f  <= 1'b0;
            I4714f5c91203fcfa552f0fcf71b87442        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7b813d83b13bb7bc13940cf5714c06ba  <= 1'b0;
            I3b6d1e84fdd1019249886fa5fe65895b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I09031235f61238b0e32ff52641aab70e  <= 1'b0;
            Id4948c876d48bdbf317d32f135e645b4                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia8a7d4207dbabc7970bf36f3fe74f72d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5402fd208dc7ca81dfd2920a9cfa2715  <= 1'b0;
            I84047457b43ef33874f4550c3b773460        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia01c82761aeb124cd92fb15ee367ee8b  <= 1'b0;
            I5e51563c3e69beca0b463742e6e5f9ee        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib1a40247057324b0bd810c844bf11f51  <= 1'b0;
            I6c8d14e31c80811ccab1b6ab09d28089        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied8bd4b6fd0e4fbcced6d20eb7435f55  <= 1'b0;
            I50b3b7490c9b65b6e662cc86b163a2df        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4ee312036de8c08300c358edcff1e1e9  <= 1'b0;
            I8351a2110a3d73ad8803cf17e3317017        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I477a920e2326828bf026b0a6b6a18e2b  <= 1'b0;
            Ice5ff01d4fb4583898498651a0ac0171                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1e6c696951688d581f21ab2302593335        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic11a6b77b84c44180eb99220a0c4c9f6  <= 1'b0;
            Ie9840e28133eebdca0be313552195c7b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If0970d9f7b053fce3ced3521b4885588  <= 1'b0;
            I82812258a8032e273cab7139266be1b6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic7ebdc317c978eb275eca41d5b9106a5  <= 1'b0;
            I27ab6fd9927518e29ed36d7a7a241498        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe3d3e6bc58efc2e9d9eb1f96cdfe424  <= 1'b0;
            I05b0f33a3808ac53b29d8d8309447650        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1dd4671765f8826c2fe20c592c5e32c8  <= 1'b0;
            If150ebf242231f0d22c996a71552f6eb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6cde57127c5bd2732e71ecb7738fad6d  <= 1'b0;
            I0fb33a5ced3d15622c9aefa188052e24                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If2d0a2b58510715e74787cb60719cb5b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If6ce2fa9f0b8bc74442ed8262b5089cf  <= 1'b0;
            Ib6745a6d17034a29501e022bd846bf2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib0001d7298ad1f3b1c7603173a70d8b5  <= 1'b0;
            Iae09c127dfe86c9f7bdbeff447c777f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I05e739fc87e962848f265e2c73338cac  <= 1'b0;
            I742128de6b237ed48e3a7ccd3788f0d7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaaaf373f7e6f55214915b93da9bd71d3  <= 1'b0;
            Id5e8fda13ba8f6d95d694d0f30da75bb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I47b0847946b0e00961233ac0101fa2a7  <= 1'b0;
            I1aa5a04e40f9b1685c77e4d101c3ccf4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2f23d4cdb6f5f827513aa60266936e4f  <= 1'b0;
            I0074e1c3ca0ff903a9201ac5fe7ca841                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ife1adea26d13bc299bb2de241ad4a6ea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia67f9b902a21de0414eb8dda52171991  <= 1'b0;
            Ifcf6c761f0f253921710af87ab1d2247        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I87b10521099179c18652c86d5887c908  <= 1'b0;
            I1478e6a9113c124bdc4361908af6643f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I84057a3b319ab3d6a2ed8f2310f970fc  <= 1'b0;
            I0afd42151925883835844cf5deef6156        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I67d57e38df8cb35ca686ac2eb44e233e  <= 1'b0;
            I2b4ab0aadffb3a1bb86f45ebc8acf085        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I23955b54e486f0f0d21a2809a9472b86  <= 1'b0;
            Iffa867719ba9c31a8756cc5e6bf81147        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1e11f0088959aa40b4ad1a047b59caf4  <= 1'b0;
            Ibb62b6cb003f0d5549c864075f23d19b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I68c35d63dc95baff41b4dc27a86d2342  <= 1'b0;
            I3690d101ae99f258cc58b4482cc378c8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I837183265ee22d080e81fea468ab0887  <= 1'b0;
            If65f587e987a51c093e8dd4df532e26c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id597e95ce8a168ab67890085a26870d0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I413b1c1985a6c9c6f202e85ff901e3a8  <= 1'b0;
            I98df60eb8f65641f9cccce4023be905c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic32c6734132776c290155a80025fe366  <= 1'b0;
            Ibcb4fbdee372353b79c460cdeafdfe4e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I624958486d181501c7a8ec2642cb503c  <= 1'b0;
            I74dbf75966d047a4a9e91c1bc793666f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I04864c28351edb33b61a103add6fb875  <= 1'b0;
            I79b8d9f9447c4c1b551ec6c1e8903040        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ida3dd5e990ce3c237e9628a9a090901e  <= 1'b0;
            Ib34b66548621fabe0753223712b1369f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id182a776b03f48fb139c28194ae7ab6b  <= 1'b0;
            Ie5b3eb4c00bedfaecc3215d43ff28362        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0c5539373b3868d0664a92157b4b4226  <= 1'b0;
            Icf3a1b0b6dbcf959b44379024f3c4169        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic0191941cb968bbd7644c21767423d2e  <= 1'b0;
            I33d7e77d08590f0dfb1867e741dd8b6b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I918c2bbe7c71f8c6a07b0bad8811f4e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I163cf58b9a308e0439a8dc7c1526e6b5  <= 1'b0;
            Iedd960a21b1c08b4a5293cff200218b3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie08ad9bd71329858c1742c8f571a1c36  <= 1'b0;
            If9722c28747df3a59b0ecf8200907e98        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3c10d579f80bd0106506ad047d75f188  <= 1'b0;
            Ib83df72c8b73a333d0699a8bbbec16be        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ieca2767ac27170058499d83016447aa7  <= 1'b0;
            Ide3798a77f709a9f694523338b081f70        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib9c194ec16f435a9357cb344cf25bdcc  <= 1'b0;
            I0a9722a805604433562f85c62b168b96        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic920452d5997a8477724fa78c86c0fba  <= 1'b0;
            If9480ec13cd538ed03a43e56bd6264a6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6eea5fde8e2517554ad6ba25018572dc  <= 1'b0;
            I433ecf86b7704c5552e5fb5cafe0d529        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9ad2f6fd2d7f68011fc926ec9abd5c34  <= 1'b0;
            I678c22563e0273403b046df4261f21cf                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8326f0b2d25139609e2c5e466724f224        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied33f18cbb778d5ba744d249f91c950b  <= 1'b0;
            Ibbe211d9955cdf2810c9003d1fb78074        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibabf61085ca7af8dfc7927b3656a76f7  <= 1'b0;
            If15e950b569a92b590127d0ca6f20a16        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddc5b5b4501f9f13bcaf22081e5a70f4  <= 1'b0;
            I03e0532841ba39eb1d4ae823c4de2f7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I67f87fbb746dd937fffc534c596f36c4  <= 1'b0;
            I1be81a7b73987ee023e396cec87312d1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I45bdd0cfe107da0d57cad1333bf95e3b  <= 1'b0;
            I4ce1a767a78673590c4074f3f03bad8d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4d54dd2ee2f32909098d3cc2b6689220  <= 1'b0;
            I57806bb7da625881e68ae315543f70d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7bfb4c5d9e22d1bd8811844d9c74dff8  <= 1'b0;
            I8b0ab476b4790150575abb06bcdce2b3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib9d58222da98f29fa302b4896594fe26  <= 1'b0;
            Icca700c12ae2e8155ca6b41e692e8a8c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8846a8961b7d557df4fc62dada679c33        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iea3e35ece9fdb3aff3b9ff5369e9a7e0  <= 1'b0;
            I7909a0f96a92e93f95023cddc742a5eb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic44eab478be232721e7a43d14beca32f  <= 1'b0;
            I43ac4857544c0fb79d04e850435ef673        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifab075b1437495268b6a3be4cb022e71  <= 1'b0;
            Ia6dfa47c465325c1d9fb9b9c5ce08f01        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2919272e9ae3996a3e1d602ff72ba86d  <= 1'b0;
            I2e9eda5bea0cc3d88359ce8a7a82f21f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib6fbe376477afa58bfcc17a8564f78b2  <= 1'b0;
            I53ec2486418e41b2ccfa8fd82777eaf0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I659322a9fd0d5eac514437b02e0491b3  <= 1'b0;
            I18387c05cef21970ecbc39c20a87aafb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic68f500938d80460ffdb33a0adc48298  <= 1'b0;
            I2b23eae78cb925008ad59f45e80e165b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If5ae6fbf843fdeee17945bc5ce81aec8  <= 1'b0;
            Ic69eb7677638a90b7a54389d47be46de        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I94460b6ce7b776bcc5eca149eab80c26  <= 1'b0;
            I5ed74e81d2497681af5a0ca13fe23088                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8cb9a216f4da7c27f678386cb214c59d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3347717ba9556e69de30ce7533d4f5a4  <= 1'b0;
            I48cb720a6323697084ac3bbd8fcadfcb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2db290170ddae8dc52ce07edaf48b365  <= 1'b0;
            Ib8dc3c1885c92cdcce7fcb58d65d03e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idd775d9fe6fa8dbdbfb07d4071b9caa5  <= 1'b0;
            Ic3aa51a5c758405fa6e2dbed707555b2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6cbc06919b9c695d99621db6f8d768cb  <= 1'b0;
            I4d418179c859feb8bc7d750416bb1004        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5b8a1e1a6b904b0f6822c224ee0486e3  <= 1'b0;
            If207b2adc6f668f85cb76bf54673fe18        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3f5053e519a928640ae49cf4e5b39d1e  <= 1'b0;
            Ib08b8067ea75e210e83526ca4a37217e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7c965c047d862c973d09a81abe03a845  <= 1'b0;
            I95b30f641cbf7bec1886643c4468017d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b8023f4dced915cd52c91bc9d4ed78f  <= 1'b0;
            I1978531a6f8d1d25ee6d404025ec4753        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc6b6357741c9887a9db1037ccc2d922  <= 1'b0;
            Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6c9698ba88db16b8d22ccebd58cc541d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibe97860165dc5d9a076ebd935385ae51  <= 1'b0;
            I0d8ac5e09b200a55bf5ba6f834cc9174        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I777ee54ff20d0544af18ad8a870d6915  <= 1'b0;
            Ib58b7d3d77a54ff1a180c6fa5f1400e6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id18c5a1d4eaa73a94e699e5f9e3c3d35  <= 1'b0;
            Icf6b990098b7ab91800bfcf1e643153c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I72939e49bf2d9c6a84e404419fc644a1  <= 1'b0;
            Ie4308b9ac6fb6de9329ba02b1eeb0e8a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I57b7b48f13436b19a8d6a47e014eb41f  <= 1'b0;
            I01d4f02a356c51d7e4e1993de0d8eebd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia3ef2f70c5abaa852586a33c505aee0d  <= 1'b0;
            I36c351e3641b01cc43e1dd5de0a649e5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6d423a7d17e05a3c597ec6ef6c5a7cba  <= 1'b0;
            I4fc983e94c5b8f7bafca61fb0d351c08        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I48e3309c61918c3991852b45d9c72ea5  <= 1'b0;
            I1fcb82fdf96cda14a55fa6358cb62c1e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I472352e7027b9df2fa957d9fd68443ff  <= 1'b0;
            I26010e26e22d8a2ea831e86fae34a24e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I665e54ea6bdca483149d3b7f3ee42a2b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idbbf2ce4a30787c5f07c3b908a73da75  <= 1'b0;
            I925df2307b5af6d1b166e5435641d3bd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibc9a860879ccc58c815b9f6caa23320a  <= 1'b0;
            I9b14f48aa357d09e460a445da86cdf89        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia71cf07b645c58cffe33be1a9a960eb2  <= 1'b0;
            I78e94ecb6c92fa8ee24edaff33b6f82d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0ceb14ac0187d804f9692e0c55b8e941  <= 1'b0;
            I5ebeb9ce5adee72a7c9527ea6d3a3028        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ief18a19d451f05f6051e3cc8de16d73c  <= 1'b0;
            I90d7b28ec09142ca8086836fc0c5ea0d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I30be0b18e4415ca50f2d8149efaaafe6  <= 1'b0;
            I27d9985415e6d0b117e5a4c2863aa7f8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7ec15b73b2811b44e1e50c74a9f921e9  <= 1'b0;
            Idf9b563e5d10c2bdbcc07e81d74467eb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0fd2f706e374a4eb57ee26ab50201e15  <= 1'b0;
            Ie351922194483938302ff6cafc477e4a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I44f170d02bae7fe044456e125a98451d  <= 1'b0;
            I578efe5c2c504f12c8f2466a7f734215                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ifb2da5faf236ca8636677bc1dc35c4db        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I30c0fcd89e0cc7c5fa348df7b4fa2ccf  <= 1'b0;
            Ie15825d216685ae241b528fa9c158ff3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I13a98f98c54b2e412cd88c96f016c41b  <= 1'b0;
            Id92c2d8bc61245c0c8e40bec2424c3c8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9890f7fc708c7b8cf460849b4a30025b  <= 1'b0;
            Icd9fd8d7114b6e894dbee493b6797df6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5e69e930a318dcb0594a823b3129d650  <= 1'b0;
            I29ff688c085f2b18e7a3af969f18af76        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I403303228c0df825f67436f4a7e64061  <= 1'b0;
            I6d56db9fcfe69dfcd747521a1ff62297        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I946246be5b4745508b7d4b578f83aaa2  <= 1'b0;
            I2f17f7c79a0118b39a63894917c6affa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I95f0acd4f955058041c035789c3a4d99  <= 1'b0;
            I7350af5d5ee09ad28c459e3674a829ab        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4082b3564c1949a19ed35bd5a88e1ef4  <= 1'b0;
            I67b6415c5135e3d6a41d56d98d3f8315        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia7606050c683ecefc510ba92ac539a9c  <= 1'b0;
            I4a6fffd8bb7244599383f2aa3a1c8916        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5446c1c323774715371c73bd1be66697  <= 1'b0;
            I7dbcd21016231546b76aab175cac9f74        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3a8e9e7d2cd6751e8500a5567cef5acc  <= 1'b0;
            I9aeff3dc44ed0d0f32518590a900dcc9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I621b20d29d3a9a9f41065bc3c3bbd2d8  <= 1'b0;
            I988b7d5d56d22d2c77c5c8c125129a50        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I263aad78110a1136eb7012c6983b2a8d  <= 1'b0;
            Iff35cd97f2a6d37a7861b9cc1a655ef5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If4308ed204e33952c9931f8fe257aca4  <= 1'b0;
            Ifb3f2a1bedfe41c73d198046a2a3f177        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddcfab4a7022e0f12fd20cb34e9b9d02  <= 1'b0;
            I37ddc6ccbc188a3eb8c33a501de820be        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I759409e242eaeb144a53e630a8cfd514  <= 1'b0;
            Ida86d05f907d23ff9fed06927c2ec9d9                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ica608f1136da397e2ab61bd4a5d83201        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5f96a68d20e3ebc71dad4b43305baa20  <= 1'b0;
            I80636a3df4541bf29780bcb4d0ee48f9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5d92fdff96b9cd64f3af2b28b13e9956  <= 1'b0;
            I9ad99d544187db3cc7090b92c9933a31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iab2f643f81921ed8464e1bbd9fa8c68e  <= 1'b0;
            Iaa8a2b6fcd469869efcf0b75ca38e68f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17d7f36fdade16dbcf621fe302bd7e57  <= 1'b0;
            I9a171d2d8eee362a0073ab7b139d3037        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I23afd747ecece714e32fbb896b5c022a  <= 1'b0;
            I84cdcba86bc5991feb391003cd7be40b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I388528eaf83566cc56b23485a9c05962  <= 1'b0;
            If9e5c3a848acce5daf570458f78f6aad        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iea424dd9d8916c4951b8746408b8a521  <= 1'b0;
            I73247d4348333f67a491fc607b15af0e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I73bbf90b625d56f663ad10f9d21d8e76  <= 1'b0;
            I021c745eee4b85a2cd91d9d8d2b18b2c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I41796b587316c600bf583edc62649bd8  <= 1'b0;
            I1381c0a0bd28b1c5542992084635b355        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7009c18515dd43d8dd2e5d1ee6779641  <= 1'b0;
            Ie74eeddc21428254a8fc4c3e293b5eb7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I797c9cb725f88c07be28f017871d17f8  <= 1'b0;
            Ib1d0f94258b45de4bfe610086d8990c5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I06b48093d4c9b0327c3efc6fa4ca7daf  <= 1'b0;
            I138d6d5d60df37870cdbb1d9c51a94af        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I04c734eb876aa722e84d6b9edd297978  <= 1'b0;
            I706378735e63e15c8d5395446ea41db8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifb89e7ad8ef661959d82b7c22f187243  <= 1'b0;
            If8680a7fc4f5532a660006bf4ca6a66e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id1dce2b9eafc35fa71df33ada4aac539  <= 1'b0;
            Ic59d1ff3051a95166c3c2d5a2881221b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied19cb51636bfb029ba8a2c390f97105  <= 1'b0;
            I9d9f8c7a23d9750ec44e706bf763df76                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I54a551af28c505601cdfaf8faaa94afb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie46b71f55aef4d00168202431d47dce0  <= 1'b0;
            I6a3124c03eb83d41c16704133bd1cfde        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8c0c1a0a35f4f7a688f516c567242d39  <= 1'b0;
            Ie9ee27b9761af611ab96f0010abd47a3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I53222c82827cab7c770e057ae91bc10e  <= 1'b0;
            I305436919f84066a22ab1417ebabd737        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8015717cd36aabbf2cf4aa3a5c234690  <= 1'b0;
            I78e63717f436493b756efa32d66cdefd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic0c13c9a929c8c46e8702cef74de8955  <= 1'b0;
            Ic965ba971642db19ca773eb68dc0b9bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I71d7f72d83b7410de31e09ea96adb95c  <= 1'b0;
            I579480a66a5f6331fb46de13090ce888        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1db4ea6916125702e7fb09d0f742e60a  <= 1'b0;
            I38d78b447217271a63f30f78b424e2ae        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc445d3f5b3b62562b0ac83e5f17e92a  <= 1'b0;
            I4c8d7e5474b19a7c63444d0cb6143728        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iee6e52d75c093a24eb4e5e0b45feb256  <= 1'b0;
            Ia4bc4b7414bf31305ec8f63e7eda61e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id48fe0672aa98f987162931527e9f9bc  <= 1'b0;
            Ibbebe287d56c7d627f3ffcf706575e77        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idce46f6d03376bea1ba361e8c59f8bd1  <= 1'b0;
            I83867e6ee369fff7e39ef5c8d5398fef        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie79ce8adeef2c3c24a3386f054d0cf5b  <= 1'b0;
            I1d40df7dbf99674f987bd06db714a702        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0d41bef808860bde56d48792764612d5  <= 1'b0;
            I92f42789cb81760ff2973e3a5fe915c3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib6ae81df8db1dae269437861ee11ec0d  <= 1'b0;
            Idbd5f2a25ab05808721cf9c403017565        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I33ddee677715877c11a1df45cbfb01ac  <= 1'b0;
            I7ca5f07d6d3c2a045dfd55ae5214dd65        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I433dd5092cf1851cd196feade3cfa6d8  <= 1'b0;
            I0b41b002a32b8e9e2fe68e819f228fb7                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7f4e1445c68abbadce23944b99d206f9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I71d3a999d88e591e102398409b3adebf  <= 1'b0;
            Id9f28016678e5e2127d9f0aa93e0b534        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iebecd2d19f9174d87deedc1a273e7baa  <= 1'b0;
            I6b939c57a8b7c7c51ab43e1b1df12f6a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I168afc1863f909dbcb6a9230db9f3e00  <= 1'b0;
            Ic5d0df586d56bf4cb322d4c3ad677385        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c4b29e48d0effac4839037ae5688334  <= 1'b0;
            I2e287724873cf6761799eaf464ed6302        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I431fc2e9533012c8571d8158d4777dea  <= 1'b0;
            Ia7a10cffe31a53aafa1104b97543280b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ief72606c77113ae37845e4aa4a2ae5e7  <= 1'b0;
            Ieeb089c6a18791a2227c8571913d689a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I641539560711ff1824bd90baa0f21f96  <= 1'b0;
            Ib29b00328971c3cd67209a5ea5b63b0a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ac0799861144b599995318bdade2114  <= 1'b0;
            I517e0868f2bb9a22c287a1f3eeaad2f3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie83fa8157a7cce44c2e25f46ce897dbb  <= 1'b0;
            I2bc9f76469e2a3f9846560ad1975cf54        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8be4711146486fea913843e497065b50  <= 1'b0;
            I9f089315e435cd69d2929fdd936a8a77        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I65171c9ee8449407484e5c82d13c6751  <= 1'b0;
            I9b54c9fb4179423c731217286e329930        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7353ebf3a1cde89d2bb3fa667f7f5485  <= 1'b0;
            I82fb41ab743146badfd2e82258afb310        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I669d34b955d2991ebbb31c149ad1b6f8  <= 1'b0;
            I5619b91de99eead78befdcba1c62411e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iabb01dc9980b4879a7356712b51df0d6  <= 1'b0;
            I83dd2047dece99cd841b2e7955819d57        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I373841aa2bcbad8232d54ac9035a3ef9  <= 1'b0;
            I8c927e66ccbf4d19f07af5ef9fbfe3fb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib6124faff821158c6a2c9a9c454ab68c  <= 1'b0;
            I0e872d4c07169cac84549178fa144274                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0793fa8938acdf65486e5582d01b9e5a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6f7a45fe64ffeda9ed120be3a4519aea  <= 1'b0;
            Ied68d7ba0ee9974eb33767e737760b4d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id1dafb7e45b860d506e0c2c91b28142e  <= 1'b0;
            I95ba37056659b29fd4318a68d85445e8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5f1609647f1e71cef4ba2d605c6c8445  <= 1'b0;
            I08d7051a18f358d08728f1c401c15c47        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If17c0096ce34b88007247bf4c429d5c4  <= 1'b0;
            I768b6f55827ac49eb6ac2655e9397be1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifc2963762403a00c4f3662b2863c991e  <= 1'b0;
            Ic66f737fe60c55d4c10e5d72b307a061        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5fdd8e1550feaecd81b82069fe73ed7e  <= 1'b0;
            I5653779f15c6c9b0f3b26927c48d6234        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I85654bd3a07b4329aba17d8b27777f4e  <= 1'b0;
            Iac550729fc437fd67151fab57134ec88        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibf2a253afde05c905d0b2404c5a808a0  <= 1'b0;
            I853b03c5826eedc3c67a2fae7a640212        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ade5535a79ce83857481ac771cd8618  <= 1'b0;
            I6f4ef0f404ae046519b8436171d51e09                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If46a6b47c1c52243cc0bc92d1edb594f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I221524a69e18854f029cad30e8f94e8a  <= 1'b0;
            I75b36a9b429cd657afc8151b9613aca6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied764ee7730ad129b6f62837ef50774a  <= 1'b0;
            Ife682dd9f677da4d27294fb61b141948        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic98f33c6a4613534bcc9b6bc4b4f2d17  <= 1'b0;
            Ic2b6177a9c586b274b68b25584e6df2c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I92eb6f60c14ee9eecb01718b01ea980f  <= 1'b0;
            I0d23011c4381496a19cced7bf7960546        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I97e82e5f6775d1e31537b891597223bd  <= 1'b0;
            Ic5992d5eaeafd5dded641a7d9801e763        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iba1c0ebd9cefeb0dd7f690bdbbbfec58  <= 1'b0;
            Ic9e7fe68b9045c6c9eb86185b5f5872e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I235c3a9fd3e8ea1cee762c10bc8e2c53  <= 1'b0;
            I51ad746720b5e6e09ab50f0283552f1a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idd474d80b50992537d6f527faf279800  <= 1'b0;
            I0c8964888a1315507f5d71959dd24cf0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I88a89b2d938552458dab9bc34728959b  <= 1'b0;
            I4d04e66ad9103a685fbe088b74517452                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id4d4f814a0bb3418cbf70c306acf048f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib105151d91678f81978495ff94b1e651  <= 1'b0;
            Ic91bd7b4bd148e526ca21d4a5ba87be9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4edd64d1f1da865b1eb886e22726a033  <= 1'b0;
            I7959dddc32f0f181b3ba39149afe1016        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia7c9c24f8e993526e76c6915e56908c4  <= 1'b0;
            I087263600b5f38be072a4f1db787aea7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib0dadebad37d9ea9d01350054872863c  <= 1'b0;
            I78d17a56de5cbe08191ef23b9731c485        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I76fd9005abd511c3c5bf6c77de8bf2f3  <= 1'b0;
            I82f713a43596df3b935d6da6f8041dc2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic124975d36a292816146a2fe61ab3ab9  <= 1'b0;
            I422987396853a6a39dabb6e7ddbf91fb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I70a4926e9e6a05fa9ee51a26988862fe  <= 1'b0;
            Ibb6556671e104141dd33188ea5fc024d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc5e98f6958786ccf95d39b922b42ea9  <= 1'b0;
            Ie42ce76076a2a5e887e0112086012da6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8879df010bbdf6e5fc9370e2fb3289b4  <= 1'b0;
            I988e525020c1e43d238fad41dab4e6ea                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4aea430599b9c0702b3bebd5960b5c91        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I94a9de743d5bedbea3876de954f479bd  <= 1'b0;
            Icbe11a3970136e485eee1bc5053e7273        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17c9d8f658dd6b2916b645d103f4702a  <= 1'b0;
            I0a7f1ea1719c1f5ff104445a4130a5a8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I384e50fa8daa639124f083dda56fac00  <= 1'b0;
            I1802d759f26dd919bc315bfd4156238d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie165d0729542c81ca89f45d15e0afd3d  <= 1'b0;
            I2148493e253783fad70f4f2807b83008        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie8e29053f122a9247b0dec291c6ef4f3  <= 1'b0;
            I39e7f78d33aa7f50264908d2efe23634        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I453dd7d7c0a2f003f0b67e909630d641  <= 1'b0;
            I844be5874def16af98de935019f35fe8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5707d30ca29842b6a96cfaeb44ac6668  <= 1'b0;
            Iee5172ba70a6e368b4903f9ff1d93471        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3fbd40faa4c3b78b547b8348c466fd1f  <= 1'b0;
            I1f34b473283291e0970879465c005e2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9a403c511fe2d44472ab319a9477199c  <= 1'b0;
            I90d92887cb2526a2956d5e8c9fad760c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie1e0b5120737a7f4bf845618ccd22239        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9db50007841762c9a10f6b7e9d40f858  <= 1'b0;
            I8abec3020ee5358f8768e5595e9992b4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I89c5af1a6176cefa1f77ee69996473cb  <= 1'b0;
            I6fe683073211a484cb6e3c416b365d9f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5ede62333e0f7ddc5446b653ba9a2382  <= 1'b0;
            Id7d764da58ade36853e8a45b5ee19dc3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I69d82ab774d52c219509e993e7cc4deb  <= 1'b0;
            I3cee2fdf353643deac7d6bca20c8fb52        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0eaa22f5eca8f33dd254fe241017a098  <= 1'b0;
            Ie9b8f8f0434fe3783c3d8f68fef30e50        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I570c036d0237c53bb069c52d621e539e  <= 1'b0;
            I68cba8ad7742cbb34d0b1fb16be4a58a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9d7614d286377329eb3999213889b707  <= 1'b0;
            Idcea56657d40e0fdf9a1c2d920938fd6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3eab1582cc42db0ac7739386cce2a712  <= 1'b0;
            Ic549ffab8f0ce161a177faa2ffd1326d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie4827dc0983c1a63053c08de6e36d375  <= 1'b0;
            I4d463d500f93f74b2724972ec1d62439        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2eed3d32a27d51036e17c4a21382b4c1  <= 1'b0;
            Iba2f362e263953331649c726afa9c481        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie039ab562e9cf90289047b5425186123  <= 1'b0;
            I6a053d931fb030e03d4882856d3bda75        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iefbdf686d9452a62cb99cf023a4d9fe7  <= 1'b0;
            I00fe3792cde1eeab36e576fd6634c4fa                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I27ede93004e0c240efaa56cc8c570910        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idc5dd6caa4ed17a63746d30d381a944e  <= 1'b0;
            I61a11c1711ca10eefea3438722b40bff        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17086dc5193aa55e5c6f56ecd365cc00  <= 1'b0;
            Ia7924c88692cfddf24fb1eff66eacb7e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib2fe0f68044c11f879e512a200f8099e  <= 1'b0;
            Ibcfd01e622f7f5a5156dd9b335b4e5e0        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I768720af835b02a8dab376ef23d17a15  <= 1'b0;
            I7f6f418ea51b4298da8758bda3f6a21b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1d98943b01a6a2d8c4db18b98dd62f5c  <= 1'b0;
            I7185da8937449e23abdd0f39a4b3ed7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id3b089fb6edd5bcfdbca142fddd5ff89  <= 1'b0;
            Idc3e3ffa31d9b76c7cf9358a5b2e65d7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5196382b75d16892d550f17893de15ec  <= 1'b0;
            I31fe8c887c4aff7c69336676cd31aaa1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6387919f2426c283e2d70e471cda54a6  <= 1'b0;
            I59684d5fe6bbb4b54ac097bd25fceef5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3b84dad6d0dd8730312b3e20c6d5a2a8  <= 1'b0;
            I86a7cd69148f9590ce91d0aa270d6c54        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2a4bbedf880a9a7b4e1bf946f9f96c0e  <= 1'b0;
            Iabce1ccdd968980f622f0e137b159d11        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I49d35ec6369de10afb15be8e0cf135c3  <= 1'b0;
            Iff02977d7b4c733cca1794246f630931        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic3ba4531855366e9a060cec1c7694844  <= 1'b0;
            I6e586c5ac59a28b30c377e51287bf04d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9026c904e5ead7ff2994c4f781d61466        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4dbabfd592b74aef93b819163130ef5e  <= 1'b0;
            I99d7489ba87c629c6dd9702a9bbfd3c8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9ece87047aec25abc02a5eea72f0e647  <= 1'b0;
            Ifaf191e0d00ba6da7019c2efcf08e1d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ed6426fbdba8aaf1c948cca7442b3a6  <= 1'b0;
            I4c295991fb08c90862a2f3ba6489000a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I24075f37c6bbd90c83370de1a2e58af2  <= 1'b0;
            Iee61d179da125934298400256788cbb8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3175159add7b814df637c2db8feb43f6  <= 1'b0;
            If87c84440426fb24070372dc1d4bf315        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0a569f6536789efb7ad2377c11842830  <= 1'b0;
            Ib9259a807b31c1b7a528d336bfc403ee        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iae6ed7748692f2edf1aa9d73380075f0  <= 1'b0;
            I411c4d909b2a571e685cd703245516d7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib4ae1cedd09d72c235765a6cd7e91366  <= 1'b0;
            If8425453cca8fc8623cb85375c4b8a1d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie2d946edaddd3c87f328e861f3e72c0a  <= 1'b0;
            I654b497f62df75fa283127b5de29b1ad        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id6b508145cd21ba088ab8fda34577c35  <= 1'b0;
            I2768519342f7b8a1ee40c1d5ac502b66        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifa6e3541f5e12bf9677ffc51d0392749  <= 1'b0;
            I8e354c1c5ba44fe5430887248ce0c43b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I21e72a7e5870151c3247d15121e5fb4f  <= 1'b0;
            Ib5dc74106d8841d25a793010fdac599a                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8970d8a8aea29913e8696c14c153d16e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iba283e99a57d0a3b78ad2e309c316b65  <= 1'b0;
            I3555c6e2fd480a6be11549bf95a9b0b1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifba3e46933049cb093d2c1809f3a8a3e  <= 1'b0;
            I8d5600a352e8ba4756f917f912fda6dd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4af3e2bf2ebc913ac902b48da672c5b6  <= 1'b0;
            I7e99d73c95e7ae5c3fe07a3c60ef52eb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifbadefd3a7ab50719a703400ddd742c6  <= 1'b0;
            I831633aebe5c6a52b98d630205376f3a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2042aede3390bd208a281f0380c95a4  <= 1'b0;
            I82e35482de74223be0d2558334ac2dfb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I19b73c5c93a71e90f620572f23f0e6d2  <= 1'b0;
            Iae2a6f9649ef1bb193e4f0ab5ecbc3e3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4b99891bed4f5c149cd4a5b4f1dde0f0  <= 1'b0;
            Ie8eca65d791ad2f6e8f4ed244f22ae3d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3472ee8c06644490252e606b62bf9bd5  <= 1'b0;
            Ic24146b01094df9b9ccd455a791f239d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idb1efe99b5d7fd567a7f82cfd52f7eb8  <= 1'b0;
            I1c9031fd54ff9417d44c9fb17dc1fc63        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I24f82a3f2c0e8df486fe495dd95cf8bc  <= 1'b0;
            Idefa20487bc5ba6daff03e6b327d76c6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I83ecf12f3b38fc14c3b75e47b71ecc09  <= 1'b0;
            I6f984fd9ea27b40ab3afeac8afd29ade        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I74cbc0ec3bb682e0f927890eef8d7a58  <= 1'b0;
            I3eaf142d2734d2d0decef084dc037b50                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0be92debced4961df5f461fe81e80bf1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I989dda9add29306d7b3c0f376822763a  <= 1'b0;
            I2d171ad83e27a3745d204849a6f46954                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia7bdaba4c6601b7146498aea6c9a3e07        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibc929201e2eeb3e61cc8f0acbade497a  <= 1'b0;
            I977f1083f5e4f6f8ac38e2c5aecf1b79                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id450c0a1cabe087be051fbf4158e6016        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib0dfbbbca2d3d264065f73b4241caed5  <= 1'b0;
            I9bcd673a4293e14fd20b48fa20492df7                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I656d0d69f6e243746b87ad67764dbc3d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I339786aa60d4c71d12c65db27ac420fe  <= 1'b0;
            Icb7422ea46b22b9330c123b40fe343fe                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iab9d870dc1ad159bbaecb20a9b72f005        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3ade020bbdf8f954821f737439513043  <= 1'b0;
            Ic414cdba230d7ea73972b0eda1ec6b1b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id53b60854f19e095c38f2c255dc57f29        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia50526cd3a3174bebc5a7a0889fda661  <= 1'b0;
            Ie4e1e00503dba189b0f871c3c0810d76                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If9ba44a2e4a8f0b61692fc69ebeb82bd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie9f37dba0791359bc426a73639ce33ad  <= 1'b0;
            I721c43ab62b42a18c3f5228fc0a73262                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ief95e8620a1c8ddfd6df673a3a223bd8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9518532a8617fc8290eb6a5e981dea94  <= 1'b0;
            I1f7cb03cf806b247be1cace4d75de942                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I61519bc0aa02ed461dbb91851d0ae19e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If66524125bfde5aa48ac70c4e448b38f  <= 1'b0;
            I775cc766b069022bc00220050feee4e4                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie0c11d584811174a66ca221baf87c36b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic3ec6375998b05a3e48f6c5fe7b3910b  <= 1'b0;
            I08b78f774ed494fa7f119977bd92679e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If10f4f45ff0fd17541735934ad20f187        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0ac421af6e311b6005c3e02e93ff94ce  <= 1'b0;
            Ic7dc7f94af108ca7c8003a2d07e1e168                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I445919f07a6fa8654211301a9a6126bd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib9db80f43718305a8a8774d8d80c86c9  <= 1'b0;
            Ibe1327961152cc2d26b3f19476a6e2c9                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I64102b82893352549abd2e2132b19476        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3b775b06b5d78fcd7373c966a62f44ad  <= 1'b0;
            I5ba97de444af4e8c9744c3b707502edc                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1fc1933fe891ac26f35a42a1b242d919        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2372a5956f21f97eeb9c76281b6675e  <= 1'b0;
            I3e4f1314042010b5d7384693b580da7b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I84dfba8bcf8ad3b85f9472fd60d607b5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7b32c2b108e24750e2a24785668af3ea  <= 1'b0;
            I4a47ce6e21c1a274578397e480c184c9                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4302fccefe5ee13161f9ad49f9ddf43c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8ec99197a7d823f5745d382c10161430  <= 1'b0;
            Id184731beb200ad6a53ce273b963bb3e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I59d7153724d3b3805af799692fbe245a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib895fec0b3756932b85962c1d129a03e  <= 1'b0;
            I3317f2f6eef9a8ef1fe1ff68b47c5d03                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id1650d0e39be078027493f58e9bbcbdd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I76aab345d13c6678fe37a4a7133cfd7d  <= 1'b0;
            Ia6b9fa10c79e6f3847f89b35afb4cc59                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If40ad4aca8dbb3bf7dde8c2ff2e5b8f2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib4f368fa3d3ec11d9ffb2ae9a2ae6310  <= 1'b0;
            I91e98b804ef82eea53c5e8eccfec827f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie49f173549396caeab1d13da36e37c65        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idd0f3cfc5599481c954a2bfe69f044e5  <= 1'b0;
            I5f1e0d0c6b50f70a6f5584124e095501                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3002a0e0cdf8e79bc7186a876410d106        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie624c4dad5036a25ca314b94cf3c4b95  <= 1'b0;
            Id61fcc605b4b581f5d42024c2610c8b7                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2b50fa03f584d10e9af3be085a02a12c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibf4b3caa5655cfb6663f9b7e2383bbbf  <= 1'b0;
            Id64738b7668931553151dbadd5605b71                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If473d172a7bff5aeae99245bbb72978d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I049d1c09c15def12ba7bae95fc1c3d55  <= 1'b0;
            I3bdfb451eb96d256da542864d39024df                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ib89f7b5625995290a64bcfb143d978ca        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ide06ba186ddb179b489ba6e3e209e3e8  <= 1'b0;
            Ia740d8ccd8230b28d078b2ea3e58d6ba                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iebe0c9b4a87d58a1c55e2ee6b01603c4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1b78785ebe2e7f77a3125a6334c4dc54  <= 1'b0;
            I574050722f82569d34bc2cfae1eedaa9                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I104411bb641d2445c7e1385a809bb682        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie79c93f1703121713fb9401617f349a8  <= 1'b0;
            Ic8f7ec6ee09fb9ee2467e3cea30a44a3                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I47dd28b4ae4f7151aff5bb271e35b716        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icf25f076eec2bf81c899c66f6cfbebc0  <= 1'b0;
            I2b77d922a74fdcef0d57debc789bd539                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3a27d5573b748df459b90a5a347f9d09        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic5c837a0556d1cb66edbf0294d08283a  <= 1'b0;
            Ia1d8127af4944b23475bd7deac91d60e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2dbef85d2b2b95af39c3a98c4e143253        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I51ff4bda38746682e3cd4c68118c3216  <= 1'b0;
            I247abcede9914633c0a33fc402bf58ae                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I510d39830ae7b0a857ac11baa7c144d3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1c074a53e6c0f2467bcdd7c952f51670  <= 1'b0;
            I1f413d3e081c6aea012b122fc94f73d5                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2751a94a66ea4cb44c512df4c509937f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I37c49c5a2af240496f5a5706b0d42ea6  <= 1'b0;
            I1b812fb764d3b48511c0d15a7efaea29                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic9a003bfb70ac2da6c229fcad09246d4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia94c439131e1df5c95fc8ad3cfdba473  <= 1'b0;
            I88882bd8a9f8718411564221ad85b223                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I34ed986182a3311a8cb005b3dccc224b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I723a6fee3b2496f23c48b3584f8bf9ce  <= 1'b0;
            I232f24e2798488ee66003f3b8cc294c0                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic79281755397f6099ff30c5d07d7e6de        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I648b62fa0bc2185c1756ee531e8e34de  <= 1'b0;
            I856284e951773518eb6c4232ea7f3d40                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8d6559ccc33cbc663584923a55b928b5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ife631f9a3c4c64a3d92aa9586ae75f3c  <= 1'b0;
            I82cbeaf5b3e4796b2aaf33dcbd119f4f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4f0a4c241844e390318f11899a0f2c5a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaac1d82f0846fce1bd88ebf8e60300ac  <= 1'b0;
            Iaa7791bbc193412e5fe25000ceec23d6                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I45fffa266ce3838f82d755b59216a4d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I48cd09f035f668536cd288a23010b07b  <= 1'b0;
            I44bdc0baed3d51ef54ce2728618ad339                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8f0e65f5db47d5460d4ec2172807a3e1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I119b2e5c2fea5338244c4019884af26f  <= 1'b0;
            Ib6bc7e75ce750a26113cbb8895c2f024                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I34127c0d1af2438e13b6f4709ece80ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2bd34b2fd12f12bc301fd0d5d69c0fb6  <= 1'b0;
            Ib4188380f7e96d5afb99f5045674193d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3a67de0e76bbf29d8c77c21865abda2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib715b1e0061b84ce614a30d961a83e7e  <= 1'b0;
            I5bba219c5024301e420e9a5acbdc5845                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic64e64aeb754249b868e14311ea19759        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ief8c2838abac83370fd7ec25c06d509b  <= 1'b0;
            I1bb52988c9ba03e16b1b69335d3d7e7c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic4aa0dc9014c8445f8d9a7723d7263f5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I561d79eb079915c0b1732cbddb119c2d  <= 1'b0;
            I1b9990aaeae716f66b0f89fb02be0a74                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I47b988d017580bdfe8f443904b1f3aac        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8bb75bf828d5ef337fa6a965808e4638  <= 1'b0;
            Iceec2cf6aba9138648a3340390f39fe9                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ica9ff13e8c3850be6c70b0b06c1d9fbf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I11ba339c8250d07b497c88a39a6df1ac  <= 1'b0;
            Iad7842f3d4672f42c1064c28d4c8ec4e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If2efeb489911f295dd7722cb22ea521d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I173aa69cf52114e223ac1410d90b4bfe  <= 1'b0;
            Ie5a53cf9343fdcdb5788667c45fadc83                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iaa16dffcc01e41e6ff17e92bdefe3df5        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia4e89e99acb95f4183474b94798ca35d  <= 1'b0;
            I30e06d190906bc9eb6f1c3156c47f9f1                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie8857b9841fbd795a4192976ef7ecc25        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If4c36727ab1c29bf78f72e8acfc00d7c  <= 1'b0;
            Ieaaaced47e22029ad2945eac9cc45e6c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If12aef69eea28052aa3bdb6ac31af205        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6426943b4ab66f17c2b7b399ccc7a6a9  <= 1'b0;
            I08dc6f8e837b1f6b80bd3fc742290dab                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0b3c6162ae2b9221738a18a29489887f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddcffa815489773b3688fd68dba18bd8  <= 1'b0;
            I8eb6a9c907c5909dad6cda98022d70b8                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I08211bba29e87faf4079152bcc973e7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id00642563679fa9a6696f8e7bbdf6576  <= 1'b0;
            Ia5067b1b458af82c3c2cd50653099854                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ibff3da265f1c3f21548f5b019e1a9dc1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifda1c55899cd3506853cc82b450b3936  <= 1'b0;
            I198c6753cf12d423c709d1512e66fa9b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie9fa1762d7844b0d781afdfb0771cea9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib5d1a7cdbcba0b654c12063d4f1768e1  <= 1'b0;
            Ib600dd8a39fda48d28e1289d44d49a84                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia677d504b9f7fc2698c0345f236428ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5e8ed024e2f2548bb375a2ecf1918a5f  <= 1'b0;
            Iabf09191227584c76d7fbc634b706d12                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Idebce29121c0481df83d755b60ff632c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id25deba967318f049de8163e67262f4b  <= 1'b0;
            I4869ba08cab90a6dcbc454b0001a7a20                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iad2c780a6386674d50cca54d8c4ebd86        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I925f6b549a25cdc8f85152eb21ea3b58  <= 1'b0;
            If97974406672507f8c9a1c507c4b6951                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If1d7944e7c4828ddb91ffea28609cbc7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9b49e1acb81ef5b088b808d2e4ce9954  <= 1'b0;
            I4210341f99ac7cb08245137999739114                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I843a68ceb0adab829091f31d0de56eb6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6386a4dd26e7c36165dc265b3a2c93cf  <= 1'b0;
            Ic24f4dbd99c8f4d88c8450d4fef762b8                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I59701b9eb54dda2744a79cebe7d73f3b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia20709f08cfff3a51d4af1e81d640400  <= 1'b0;
            I68dffa1a13eb6ab54615347729c1d6af                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If63cf5e8f47e4e51176401f0d954ea23        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1ff042bdb52aac5d69791e96e2f9706c  <= 1'b0;
            I10153d5548b184b9ac2cecdba4ec4b1a                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id09454844b525697de3e3727d89551e4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaa2cbf59f6f61198b4fcf5a741cd5bc8  <= 1'b0;
            I104b7f0512440cffc0fcce25e477f537                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6d1b2ce4368945b56eee7814638471cc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I01c94743a11042e75638ba6618356203  <= 1'b0;
            I18b6758319272eebbe76e1eee5ae55b2                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6079945faa57335b1c902ccf7f960a70        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0a0340a0e52145f3597accfe4a4e8624  <= 1'b0;
            I780263b10b98f9bb0eaf66c045d8d37c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie7752906ac55cf51f3e96e8c0046f1aa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3bb4d24caaa0882a75125e466070f0b1  <= 1'b0;
            I37b772442e55cbcd44ba892a0608d662                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2d7d4135a94f5df949283c043228791f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I44ead0ab5ccc53226fccc03024643771  <= 1'b0;
            I0ac256a6659ff5c6673fd110a8bf578f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I99c75e3d26c5d01f6ae9abcd05407d8c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iaded125f7fd5c833e7206dd7071069be  <= 1'b0;
            If134e1d27e736005e5a390e7a2ea1f4b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I81e6f97621dbfb2fed6fc236005a2b19        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I373be7c3f9511a2906584e33e5048abf  <= 1'b0;
            I7b37b8f908cd82683832536e02faab0d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ieac60532dcfc916a65054e35cf31d6d2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie0b5f51835ebdb508a596eeebf0e4847  <= 1'b0;
            I08b4bf60c9c7e7229bd1952cc88bc7b3                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ib7eb83ba73e0dc17f69c357b6ca555bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddb75e0197b9a76b36a59ac2a7ccdf3a  <= 1'b0;
            I267d637eb63fef9f4723f7978fad88f0                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I5139d8a7a099e3c619c60647c15b7420        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I08c03198b9599b2f4590e3022e398f7c  <= 1'b0;
            I4fb56a70e5ffa71f58f715da36368e04                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6ccd2e11ebd5b2de80b120e20650a602        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia4f3cff223e24815ee1d86bf41756f06  <= 1'b0;
            I5e9e2acb258baf96ac4b525bba54a462                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie669cebe5fe39e1a841f8dd3c1f6bc57        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I56592e1452c4b559af19465b30230ec0  <= 1'b0;
            Ic40f61443a4d8f87769067fc39381cb3                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If32acb9fc212c4af34099acf6df2bc5a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I213ce488e5345fa405a9c5df297d6f74  <= 1'b0;
            Ieb36710c9a3726f33407436d62639c8d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I075ce236a181bf925c8ccce91d9bc8cd        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iefac1e428116a797c2c0803410ac5601  <= 1'b0;
            Ic804af393da2e4b9c8ef25d4a3b4e8d5                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I541d4e422b999a0dfca44d275178e1d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8b419d5827e5b1af9649d602401c189a  <= 1'b0;
            I52e4c446693c29a42bb3b665f72d382d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I3e02657f3d9f79338cd083ed024bf96c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ie989550c9101de382056dd60d5da0e01  <= 1'b0;
            Idbf02cf10add496d30fa44bbb18458c6                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia5e5537405ab8edcc7cd43c86837d43d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I259010e323e1e8dcd9dd719091131f6c  <= 1'b0;
            Ida095585ad26e215f1c1bf989912da89                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I07ff388e3b6c7288f0f6c35a345023fe        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I389ac86954fd70464c9550e3fed4ed33  <= 1'b0;
            I19f1ffa05c7c9a0df5e7014044024c7b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I56cb3b3e193ca5068734417fd0ec4e02        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I77371f0e55b4684d1af196ed52d3d997  <= 1'b0;
            I4d68a2fe778fa93faac38b138138291f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I5bbf1765d8f81581d0cf31c0bc755fb3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5a21996f5724a2a49fcf8e928c01b062  <= 1'b0;
            I54393ada6f76ac82c31f2668e228e29d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iaa1643095e518846cdede4d5a90dff84        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id46108963921efa50aff64d4dd7d1701  <= 1'b0;
            If5b9ef84f09680f3593250b13a852c1c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iee6e12f4717a3279dd31b874eabae69e        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8da50e5093acefb6f809aed64564a53e  <= 1'b0;
            Ibb759bc4179e5b7aa759d850c7cfa467                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic52a9edbbc5283844d2514ea142ca6e2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I03b0694777d0160a83cbc82ac1397736  <= 1'b0;
            I05e8b5f8b83f07b609b5ebf272bb2229                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ice3e978c8da2a7de5b28542a5589f0a2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I85c2bffb93569d9fe1b1bcb10b98bcac  <= 1'b0;
            If6ac15373ec1146d38e7aeb71c3ece64                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I336a425aed221c85ca80b9a97d21d6b1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id00274c88b93867a80606343add1cdab  <= 1'b0;
            I2ab3675e1eede757af80716ba980a4e6                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie477c0f3b77bb299ba8b1a410d211ef7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I61e829cbf7d6c0ef8ddc11677981e2cf  <= 1'b0;
            I388c271687ab31b57421ad57192273ed                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie62920d089ae762603cd33fbf97d92bb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9e8ae2aed048068b01b3bd46f30baae8  <= 1'b0;
            I6121679cec8caa51dc5ff0d1a61f9821                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2ca952e4e676537fd5a8fc71ecfa10e9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7dab71adbe62687846fc027d2789451d  <= 1'b0;
            Ia0649b990bf5716cfab230127cd5d47f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iefd31e7ff3c829c88f60bc89d70afcf7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If1295608bd218ed60922a0b95bf1d098  <= 1'b0;
            I867a0626ca22108b16267d95c0aadf4f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iafa987a413fd8fcacfe872bc0f5bc2d6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Idf04e08c120ed116af14a62659675b44  <= 1'b0;
            I1af54bcb73d7c6b93e55450871207976                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I305c1ea420d666f258e38c5a65847367        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ieb7614ad1b1bfed3e2b0089a72fe214a  <= 1'b0;
            I91883553543d0425e9c6dd726dce3d27                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9f040c4088bfab72d74e5332e9710d1a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I589062eca318b25dfe5735da455b6fe1  <= 1'b0;
            Ie95405659701278e3f87bf1f823a037b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia2f41f9778324a06daeb185c736516a4        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If3db87afb3ea184c9e4020c5e45cb161  <= 1'b0;
            Ia42392e2104b50c0908aad82738a5ee7                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id9778ba5fbdbed4d33a092da6b68c414        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ia14bc1fcd5bbdcb60b8e68298f7d716a  <= 1'b0;
            I68ad63230a51b9b9e3daffb307ea970d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I27c2c79d0d719c71c8e28218d1174a13        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I268b60cb371b3d46dc3f8b0009f541b1  <= 1'b0;
            I7a052d63944ccf42e598efe3a95b88f8                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2a9d6a774769b12ae20bc0cee0c36f5c        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If2cd93b57cd1c2b91ee7a73a97dd19f2  <= 1'b0;
            I2b3c6d69f79c8d51e4d1614c62c44fcc                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I2c567b75f1399c069b95284f4c36b6d1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id81305359a07db527e49fda05cd2784f  <= 1'b0;
            Ifcef0e92f50e3920bf1208af5d64c632                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If3d3eb609abfd6e315eec803d2e94490        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Id8292eca087c1a17dc8b5a572a76f21f  <= 1'b0;
            I111340a19625901a3c1b95fd0bd1570e                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9c58aea7ce986b1d28f5808b347c015d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddb19725b093506e5e521d8d68dcb8e1  <= 1'b0;
            I11aec4fa85c30f6fe1fd9fa72542ef6c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Id139c7a783196941100003b6cb0cd1e7        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0b573d3a86a3111451da661e46384876  <= 1'b0;
            I80cc333c181c16a96b7bd6501c27c2b3                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I524d7614b01460778da3ce98f6aaa3d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0ff479e61d1a0cede88ebffb073c60be  <= 1'b0;
            Idc6354325a6280ae9890da33c06c33ec                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8acda65f116d5c91cbe2662ac282aa31        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Icd6f8f5df6b4ca4c81855e974db76526  <= 1'b0;
            Ibb04cf82acc4ac16599ad3ddb0c2ada2                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If67dbe22f8d22b3430215fb0deae8204        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7ce064a756dad56d37684d5d7d168047  <= 1'b0;
            I3ed096dfd8a14f4acb4d53a70cf8aceb                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9a35cd7512787263abedd6d9913cf507        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ied2ea62cfb21602645babc36e27b8218  <= 1'b0;
            I0fa07f95e96326cb0599c0c3f76e2b48                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If9cca23469c5e6001650f1f8b1360ae8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I79b85da6e5ce0b02ebd1619115c98e24  <= 1'b0;
            I87d98fbc97d9a78c2e7d6a6280e7a49a                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icc2606ae8f9a3b425225ae7339112b9d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8e1ddd7e4185c28caa71d30bc28138f3  <= 1'b0;
            Ib7ddc4dca877f7cf5697a02c3d1915ba                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I34aa1802d24e074ae54563898929abfa        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iab0bff1633e2f3ea0bfbc291f3ab5d29  <= 1'b0;
            I3612ef280891f6017fad205d0484bde7                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Icb85b3464dc40e8504c53c377e889c45        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5f0751fceaa008feba5c6867ced453dc  <= 1'b0;
            I561547649aeb5b4c3f10d9506db1f3cf                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie595a7d10b5ac84c0301fb55bebd3680        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9f6751c15237c20b0cf2175575195ea7  <= 1'b0;
            I84cc76c0079b86da7b994844c3ccb875                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9c217a672cabc05efbdff218637123ba        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6ea50be10bc990a1206cdc9e28e0c4c2  <= 1'b0;
            Iec013c508d0c6401d7eb856e7eb60446                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If20f3780b4af857ffe8083056085517a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I43c2fab87f70ea883321ab82de85f133  <= 1'b0;
            Ifd8979aac6b6b24aa560b46b18240e92                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic2e275bfa8ab3d2002d2aa374ac9bfe2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1af02ed6cf00d4cb0704b5e44c83bfa3  <= 1'b0;
            If12394e78dc913b01890b56650856a44                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Iac5798fd9915b6778700da6a14f6a381        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib71611afdd0381cc1884f5ddbbae1acc  <= 1'b0;
            I94d18aa10695f3f22b23246884b72822                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ide3204bf317fdfb993410d338085b174        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I38fc49afce0298846ae8ed63ae715e81  <= 1'b0;
            Ic90b38835dd7e760dd54067b196f8470                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ic3a95140fc1029efa17a6557bc977719        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iddc3e44d83e8253e5129b6cbf5082df7  <= 1'b0;
            If3691ea51f6efe9b165a31964854d2fe                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I647d3a46bb2c7ed0f1ec08760b3858be        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I975a87bdda30c5b6be8d2f0e4b107450  <= 1'b0;
            Ic2ce582555add38a14f5006d3c87eb15                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4816747af9d9fc8dc85fd831336ec710        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I582bd96afa764ded148202f738b7a1df  <= 1'b0;
            I58cc950ee2cbe56b7c5a619be3792511                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1f66c026a5437320bd1f4df2ff71663d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I6fb88d97bc9ed37a06b729020a1df140  <= 1'b0;
            I0d8e329ec5873db96df1ec309445a096                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If347c58c328193f420286ea27a4afa20        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I1500943c4a550e78fc169437b0a663b7  <= 1'b0;
            I106325488e2ecfdba1cf9e5201e6bc8c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I7a126c8304be920f2a920315dc61ba7f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I0b83f4ef8ba9badb27e81b32765ec5b6  <= 1'b0;
            Iff73a0085541a511d3912b64686a82c5                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I237327d6a74df1fb05537dc3691ebf11        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2c420acf428e44cdd9ca9998e276f258  <= 1'b0;
            Icdab59de68f2870504598c9ea18f1d2c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I64a3e8bb4c87b066806d33a5306a2c53        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic7b6dae3017b55dd3cd27423d5f1b0ec  <= 1'b0;
            I75604d727e82c977741f90113719183a                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ibbca6ec39234473fb517447a8beacafc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4a91a7c9b2a0f3552b8f2ef4e2398be2  <= 1'b0;
            I6f50c4d0d2639857b2dcca300c2d7b04                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I78327356176a16fc996188b83b058cbc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I99ff29c7ba68b5d0819f1e1bead51287  <= 1'b0;
            I5cd013a2be2e761c10c6a957632517de                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ifec496c87a7a2474855067305ac8cba3        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If06b00be0356a2be5074d958ddcdb2f9  <= 1'b0;
            Iafeedddd02428bd2610c576e68d4ae25                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I41584165a62caaa37ddebbf79bb8b617        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I604283449f13c7b225ea03f99f2e296a  <= 1'b0;
            I912d6325e34180e0f668f0f024e63581                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Idf0916d6b025aad6eccb98ada5ba3aca        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2b600e5f5c146ee97c4044c08e1f5ad5  <= 1'b0;
            Id1e05294dfd02df499ad0c08bb5c191b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I00ef133d5a53f8f99f35b50327e5272b        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9fe16403fc21bb1159a5e0305fd1ef69  <= 1'b0;
            Id3bb9b100ee4302473b49ac14615e9b0                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I6f0e302d38d75982d0761e306ce9f146        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Iabdb9374e5caee281c25b003624b2c4e  <= 1'b0;
            Ief32db1cfc443119b6202b0cc7bf70a2                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I127eed5de00e10a020717e796de76c7d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ibd12036702fe60b57354b3aac921559d  <= 1'b0;
            Iad7dbe9909b5eed3261adf92d3813acc                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If9aad73aefb1b225f35e8c813b85fe87        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib1639811de6eb1c38257800c201fb704  <= 1'b0;
            Ie7daf0789c35caaadbba06cafabd2b70                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I00a89ac37676521a081a21b1ec1a0798        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If926d98f659e8fe4bbf36ad2c5c852c5  <= 1'b0;
            I2bd1f9b75d9ab94af9ddceb7528935e8                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I06f3a34f2b1770ef82ddc2a732b3d4fb        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I211f8d7f97ebb8eb3e50313513abfb1b  <= 1'b0;
            Ic3d9f5c6677758810e4865779ec303e3                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I4744d64a746f16004e3bedaaa41465f1        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I304ac9f96945546cdf1b6f1fa7136731  <= 1'b0;
            I00af04882a25e2832d913a67d4d86d7b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ifae0cc6cc1c65d24bbe84c4ba938e2ea        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I7a9800418bd5c195fc47a72370680b56  <= 1'b0;
            Ic9db631df0a1a9108c10c3e0eca7bf15                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1223c21129382d41e4f38ef4bbe60c2f        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I5f6a61c9f0c67510e148e596f553a4d6  <= 1'b0;
            I749f9ed1fb2dddd40ebc28f638e02935                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I14e36e16df00adcd7dc1973d3852d2d9        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I8e313ceb21359bcc44114ab217b1c394  <= 1'b0;
            Ia45b2a24df24bd5e3c95885c8928686c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0d05ae27b53fb6939e4c2f862a8d20b2        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4c9518755c33d725221ad79ee6badba9  <= 1'b0;
            I7427464fde340780aba7f9847b4ad564                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I97a6fcc08929c3b7d15e36d7706ed13d        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I3c3cffec9f47c9979cb9503f222f370c  <= 1'b0;
            I33fd1ae225e2b881b2b41e0358675e22                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I1f04e86bf27596718836d0a09adbe120        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I68d6769541fdc3df321e192f645c667f  <= 1'b0;
            I2e21a35d1cf560936fd19b944a208b6b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie40873cfd6d10a61a94a761becf588a8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ided55428cbb77f454c2607ac783d7548  <= 1'b0;
            I249522a3d42cc75d7a6b9ede1222ee76                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I61960ed74fee948cc12bd1fd8384559a        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifd3d4f3e2a388b3c70e7704d6351e0ba  <= 1'b0;
            I68b4c43d9f40ae4bfd70d2983594392c                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I8533a3ec4be4c49166184c94761eaebc        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I17d32f292758416fe02527dfd938fa0d  <= 1'b0;
            I63145e0fec15c7e7c0de105f348bfd31                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I00be319b5bdb85ffaf3bb0eca0b348b6        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I9ce3942aba354c1fd7d6b9a39c994d7b  <= 1'b0;
            I8af625de86c04016c3424d116fddab5b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ie889c916b5af185b52ff5e2e3cc23045        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I2c6c6041c9c69c84f4d64af6458955f5  <= 1'b0;
            I54c9c10527f83b4ee4e1e22f1e4044ed                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I89697be6dcb2e7f972db498c1b1dea71        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I830a4fffe1244e071eb82c28ddc4a308  <= 1'b0;
            I972559e47c7f83bd9000ca1cfc14d8e0                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If13dfbfff7cd8e197bb44006a3db73bf        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ifad8e46fc3844bbfaf434a14f6b5869d  <= 1'b0;
            Ib97a7f941eb7ce2a867503a04ff86a67                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I87ed6c3e172c7a06bf6aefe7bf718d70        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I10a6c6a8fdb0003de1f360c148777d0f  <= 1'b0;
            I5979b55f607c71017537f2b48b40cbea                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I0db87adc849839fab3a4c9884d5a4882        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I4cde586fc28f8d03fc9934d56f7ff7b8  <= 1'b0;
            I6a56760b621f238843b091279c69897f                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I535e01a6c35fd7b455e4b79b1d4bb414        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ib83a067fb08e118dcf794902beef9405  <= 1'b0;
            Icec45bf76c241d37c9a50a5cd092da9d                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            Ia2d1c752cc4b405adb97a815e90a7b96        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            I358cf9609272a4562423a85f9b2f56bf  <= 1'b0;
            I2f6d3f61f2890e584d3063a09587e99b                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            I9ac12eb3878f6fc7dc428fe5e7f35d97        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            Ic1e9d9113150ad57954c0e369259dc62  <= 1'b0;
            I7c396ea2e959d84fd9a6964617cb29c6                   <= {MAX_SUM_WDTH_L_P1    {1'b0}};
            If46fa11dfadb0691eaaa0a40836e08d8        <= {(MAX_SUM_WDTH_L  ){1'b0}};
            If7fe3f5ccbb5b279e41fd183c8ff3974  <= 1'b0;
       end else begin
           if (start_dec || I6d3acefe6d7dfb94a5d66dcaa1bbbb76) begin //d7 for Id0cab90d8d20d57e2f2b9be52f7dd25d I37302ccecb8ae11c64170bc6bfa44eaa I1d623b89683f9ce4e074de1676d12416
               I748f85f6680918a2e992df339b4b6558  <=
                      (Iea07d1adf9016a29cffd61d183e268d0) +
                      (If92db65b39a83e1c699e4cc6d7f9e57b) +
                      (I8f2986bc015fcc64ac5e5395ac6dd851) +
                      (I355725a804e0df68b4acf96ca98f2448) +
                      (I78212ae965ab2dcb2eed0b060d6b253f) +
                      (I0b56aa7a1b7549c91dddd3a06ecbaacf) +
                      (I71412803cc5229025487255aec62ec4f) +
                      (I32fcb28a27356bc6f403528836ea4c1f) +
                      (Iad354d876cb9fc72fc0143e6f7da9357) +
                      (If6e745bb85abba7282dae1f6f701225e) +
                      (I93bb43c1b89d4c70a57bdc019d64fd22) +
                      (I7a2e554d07bbea291f2cfc18694fca3a) +
                      (I3e59b2419c7dd1553b792d536208514e) +
                      (I46894c6526983bf1ce4b503159131b41) +
                      (I6404d0df952b5bf8292c753e4c6f35d8) +
                      (I8522c402e654d007abffcb0e904af5e6) +
                      (I5ed85845c39337c37791f16e718069b4) +
                      (I89013d61c1ea8da8b1c6071cc21c316f) +
                      (I4102100fa5f1dd299af0190862efcc42) +
                      (I4939f69abb1eac56d5021e06406a93b5) +
                      (Iadbd245bf842aebb456417579a3e6296) +
                      (Ifc8ece44a4e68c3117eda9e65f3084d2) +
                      (({q0_1[0],q0_0[0]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[0],q0_0[0]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib0f57837099e3fdf1b908d78bcda4a43  <=
                      (I91679dfab57a372eddc7f9b94a231edb) +
                      (I2213c1a2b831f421707a261f5a58b1b1) +
                      (Ic53b875b2ddcba11406eb2ca39354757) +
                      (I634484f00590216c0f74f975c9c83400) +
                      (Ib3b1db2d8b669988c887ed780e439b26) +
                      (I735db8b0ee0ec98e4cce0030b11508da) +
                      (If1607e907e626902ee26d15020a64c21) +
                      (I081b38dbb37d4c14a6a9fd3fefa13daa) +
                      (Ibac5e7b6d4bf5cd6926358318f0c418f) +
                      (Iadfc60386481092ae85cc148a2c40abb) +
                      (Ie0ee5445c56a5f9b41640b57422206de) +
                      (Ie5f8620371236cb11c9e88c16b509ee8) +
                      (I8d7c1fe2e33bbd45379b0325a3c5e989) +
                      (I4fbdc4ee57a3be42b62d9bd43078d6ef) +
                      (I5510b88bfd65811b3200adf4ef975b48) +
                      (Ib57ef2f577cca54713c16717cbbd1ce9) +
                      (I15943aa74e9fbbaebdc0d54eb6a3bffa) +
                      (I6ac24c46319a787daa5c545de8c6eeea) +
                      (I52403a0454e5fa002e79eaab7ea497bd) +
                      (I634f0ce28934600a1a31ab0d8e59b4a9) +
                      (I7103aa739616a39c03e675ea0efb0335) +
                      (I0296d01fd3f9a269a617efd4beea9b8b) +
                      (({q0_1[1],q0_0[1]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[1],q0_0[1]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If75e99660e3997f53f7b903bc366f47f  <=
                      (I065a81ba25962785215583e7ece27661) +
                      (I631a3300cb6685f47da7781940ec5d27) +
                      (I8bbe1a2ace8f51aa22cca5d9fc66f136) +
                      (I38c3e3e136acb79c8a0ff850bcc55f16) +
                      (I35b2c7e9cdc53a98913e1c16a3a47b37) +
                      (Ib1a2b31d49ae476e2f1fb9acba2d5af0) +
                      (Ic72f41f9bbf470aee3c9b9b8787b31c3) +
                      (I3ea4c33a9419820ed54460eb64134dff) +
                      (Ia0d940e16c8cbd4f7544f5a5cd7d83b2) +
                      (I4a8abfa0896ce414d9b98093ef84455f) +
                      (I680be647bf2a62e0ee9b5d379dc87b4f) +
                      (If4d75f83299a21802b6fbe136913489f) +
                      (Ibddfda6413e3dd2f483c3174ea836b6a) +
                      (I33bddb0adcc2af7b12a83bf843036385) +
                      (I529f92b82248efe2cf64f7da0ec8283c) +
                      (I2f34af0036985cd94ade9cc905bec065) +
                      (Ia1a0d8d7dfd6e877f15cce773f85f5b7) +
                      (I5dd29fd1a73df5662d2b636e7285bad9) +
                      (Ide530e6f4622c8a7b101b6dce9650e42) +
                      (Ibaf00a6780325882067a79f0c4d693d2) +
                      (I16e3559c63ebfed83d6698fc9a9cd93a) +
                      (I9747a02384abb1c2dd1f52b3a5a999cc) +
                      (({q0_1[2],q0_0[2]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[2],q0_0[2]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3253481bee7dbfc0f3eac94c3252ee4e  <=
                      (Iceb7a1d4c23806b8f5824016779ad129) +
                      (I40ef50004a60ae58aedc49eb5e6797c9) +
                      (I753f92da60980736440aba814a156f1e) +
                      (I4ac79b67a8904b95f7912d24af420585) +
                      (Iad44c932cfa5c249c5e59f8c706173a8) +
                      (I10f14b6433498e3b9e9bf021b60115e8) +
                      (I96008f47b9f134c9c4274cfcfb28e550) +
                      (Id0344146d1a53d418add6d2b185377dd) +
                      (I1eede74f12d37331b399eb7136bc621f) +
                      (I3e4754acc31d99bc71525789bdee0c1a) +
                      (I11c1fc94a3bd6dffa17e1571cc6ae97c) +
                      (I5395ee57418c31e11cf847f0f514ec19) +
                      (Iff125392fa39afebae1637a19c4e23ec) +
                      (Ia6308e16fae5428f4ab6560f5b21479a) +
                      (I5ea02b5349cd4d99ccbcb6b26f0cfdd7) +
                      (I21de4f6194dec9e3c401934db92c25e7) +
                      (I57d0920119f8901bd4dea2d5f8fb5d90) +
                      (I89537301987d6da0dbe6cff3caab3ff4) +
                      (Iaf0bbbe791bb71d0f557dc71caa5fb87) +
                      (Ic7ff9cde71054c1ee9eef81eabdd7061) +
                      (I88c10c47ae424fbdcb852fbf1e94127c) +
                      (Icd2e75e47cab1d539ba9ff1b6e1d7155) +
                      (({q0_1[3],q0_0[3]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[3],q0_0[3]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia80693da8182ee2c3708b6ec21d397d2  <=
                      (I37e6bc7aff363ed0ed1f84b23c5f3e34) +
                      (I733605337bf6972630c089d32fd7f98f) +
                      (Idcb1d8bbdeaed6768c2a418c3048e6ee) +
                      (Ia89da2f1890524ad3519ab403dd0686c) +
                      (Ie33a780b0221084898c9fc5b237b244a) +
                      (Iabbd1668e0014df518ede5216232834c) +
                      (Ibd89458312687610aa166a9538968851) +
                      (Icbaf92a8e9875bcb19a1d074779a9ea5) +
                      (I80f3c8559da8e97bc5397bb8b621a0bd) +
                      (I7a0eada108891aba06cecab5071232c9) +
                      (Ie21a2c9b22e7bf8425fb5c0f33e5f4f7) +
                      (Iaa5b2807e5cc2403c5787eeb3d10ca6b) +
                      (I6da2b3a481ee71b85f3087b36b399288) +
                      (I11094e852295755925c3c61f1df81643) +
                      (I9c633aa620cca127b0ff8cf882178e76) +
                      (I694d471fd353eb54aae08a2afa7b645a) +
                      (I816704585ad393f685731104ad3ec64f) +
                      (I85d95015a9ce27a18ccbf73bbbcdbd70) +
                      (I992e7c551b4aa818606c3465d33eb798) +
                      (I2ead0e9941e2280309ab53535b1e1ac1) +
                      (I56873feb8418005b5661c7382f2dbeec) +
                      (Ib6ea4a822da2ea32e0abf6cf8a33d295) +
                      (Id1659ccdeaea3e59eb2d3f65a65ebd05) +
                      (({q0_1[4],q0_0[4]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[4],q0_0[4]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7fa3f2648baacebf9e4b59c179601fa6  <=
                      (Ic2171967791a0329f3e39fc19d0a6bc8) +
                      (I7d5041a6796c00188f74936d283defe6) +
                      (Iba7608ee0a01af103e022bcaf564bf6b) +
                      (Iedbe9d0e48bd36064f59faea51afddb9) +
                      (Ic3871325d57b310c95ca02fcaca529eb) +
                      (I42f9b1f8ef24ad56c10086852678b456) +
                      (I3ed5d0fca86f35b3d4b4a89c6147d0cd) +
                      (Ib0126fb335e32793c400a97c5a4a337c) +
                      (I20590d8fb97ec0b2164ffe17826136a7) +
                      (I3c128efc9f80c9b8334bf7b61de71b43) +
                      (Ic7147944f8835e26b9838fdbdc18ca41) +
                      (I698b1dbc9d8664d1c86c7a763d97b3b7) +
                      (I508bbade361787127e1a2e8687ec884c) +
                      (I2afeb2a7b199c0c6738938f156ae4274) +
                      (I86255756ddd1f88b74e070b19f8c3bfa) +
                      (I7d4924388dc5373ad7936dca76797473) +
                      (Ie317e5ea2ca4ba2060d0f491290af96f) +
                      (I56ea52c50a188ec47e48740839a031c9) +
                      (Id9b9a8fe43992ec0793845715dd2226c) +
                      (I93b69bfb228db4b569a6772179d603be) +
                      (I71afab29cdb962e1f1ca21b61dfb50c6) +
                      (I9905e2686b350e8a6e7f790563a91294) +
                      (I524e78ae6a4204e17ba4532dba047d4b) +
                      (({q0_1[5],q0_0[5]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[5],q0_0[5]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id7699f8f89380c315303644fdebacb32  <=
                      (I71228fe4188ab1d9796081184a422094) +
                      (Ie19b39200436b0bfca13502ad36c21b9) +
                      (If6657f90c84ca5e2ba08ec705f34be03) +
                      (I60ec7459bbe99fce295406bee1f2af46) +
                      (I29ab844f80c105d247c5c15faa35863c) +
                      (I856fa68463aa5ef1ae53442699d38b33) +
                      (Ic3d00a27f15f8983a120395082854d6b) +
                      (I6b1d01c3cb8fb51e43cdb788b89816be) +
                      (Ib74a56900c1f8b159ad381f61acee801) +
                      (Ia5eba52d169755c507b9e0094e467fab) +
                      (I0899e8fec1a7209cd94757c0b2f87c9a) +
                      (I08ece7cd684e593e02321612b7a88cee) +
                      (I691c84d81c60a462e28e2b2bae3ea845) +
                      (I58dc9cce6384160c0a85c6efb3319cdb) +
                      (I56bf74b5890ec67090f499afdc0a9c88) +
                      (Ibaf2f1f8bda2f6b932dc30f8369c0e1f) +
                      (Id9364a29fd79b52d0442e18dc0227854) +
                      (Ica3a41ace27f7d94377981079952f4f7) +
                      (Ib57795a63d642a73456324bab41384b6) +
                      (Iabf572c97b48c6a7dcc19e56676e3a82) +
                      (Iefd370d0df1a93639af482f78a1e8706) +
                      (I995d2809ffaf0ecda6a004d01cb9c8c4) +
                      (I4e8ebc46bc068c3f9889d970db131112) +
                      (({q0_1[6],q0_0[6]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[6],q0_0[6]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibf3e1ead3776901898d4b154aeb61267  <=
                      (I7b561638da1b4a45ff59be81243e4471) +
                      (If0a3b88a66a816b25f17ced5d0e8f775) +
                      (I0374ada4fe50717f2158468b7ad205d4) +
                      (I357137b41bb91e0659b1ac6ead9b5c12) +
                      (I5d70bc64cf7b3d3ef4180e082e533237) +
                      (I7d9ad929660cd212387d893266b681da) +
                      (I34be4b353cf75603301372840c2f91c2) +
                      (I14834fc8e6489775359bcecf5a37ff4d) +
                      (I633a74e4dfa841c9fd13dbb6564c8493) +
                      (I157bd468200e63385583b9045758d81e) +
                      (I918c46173eebc5b2a95e041cfd91d958) +
                      (I4f8792c18bd07b23e82bbc44b4ca947f) +
                      (I8d0a1ae4c47edf1f2b99d1175aaa7197) +
                      (I734e601f5f9d568a44a48834559e04db) +
                      (Ie421da1dc5aaea57c50d0c7d9c5a2717) +
                      (Ief5cbddfbfb98fce4812a676849b9a98) +
                      (Id113cab2dd1949d32e3c1c15273185c8) +
                      (Icfe1a689e33b2b9aa9dba692d6d610b9) +
                      (Ia4b671f3360f3ce55db0dc0e4d78ddbe) +
                      (I60cbd4369e7ba9b6532f279e5c59084c) +
                      (Ifb6c65a00d9a2c31d8b1119b949828d8) +
                      (I4a777f0dd62b19dd340ad31517c4e789) +
                      (Ib75747cb32130d44b338ed8c8af8ca11) +
                      (({q0_1[7],q0_0[7]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[7],q0_0[7]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie486617fc1d6354c7f347692cdbd894d  <=
                      (Ic7e35cf8d5cd230b94c40714f16e2418) +
                      (Ic51bb9184dfd103703cd0c6ad6edff4b) +
                      (I103f1449c78c47396d6a54dc1c810934) +
                      (I56b3a97dc3037f0bb2eed93a9482c813) +
                      (I51e98035b35a35fdc52f5bab8f19c152) +
                      (Ia6a7f9beaceb08d81012f0e72171252f) +
                      (I21b062856ced09cb9131c01b5e166f32) +
                      (I4f1221ce7880729fe584b42ef3afe6b2) +
                      (Ie7f3f1d6cee7f02ae1b17740ed54c049) +
                      (Ib196f5bcf9152703dc32c5101076600a) +
                      (({q0_1[8],q0_0[8]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[8],q0_0[8]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7ba403c6745e7d026282ad704e065702  <=
                      (Ide9ef5a16d8fe32353c2c2a30e8ee3b0) +
                      (Iee6f2484a381bd42e441ff072ec582e4) +
                      (I53121a39de0bcba91a4d0438be2ae958) +
                      (Iff7950f24f0a6b0073942c37fff49d37) +
                      (Ide86f019e9573706c25bd8b4552396a8) +
                      (I2370042234b0e93bb66e44b97fca3e43) +
                      (If9efe7a1c359ec03014a52870ac13aec) +
                      (I6a6eb62960b616043415406ebfc21346) +
                      (I06c7728ef64be8311f48d10d766d0c44) +
                      (I9fe11f6c8147391aa4a5afd1a4e4f731) +
                      (({q0_1[9],q0_0[9]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[9],q0_0[9]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I93cb3974b8594665b2e7ce5593fde69b  <=
                      (Id50edc56fce48130247fdbc42eeff9ea) +
                      (If3e5161254eb9056914c46263b865c10) +
                      (I58703e8b6d04f8c69ac38f5fcfdc4efc) +
                      (Ie1f41720e296ced1b74cb325b666d88f) +
                      (I5d5701435c96f1078e741921b56e3c65) +
                      (Id96e744d9b10dcddd1ae0115ea57a76a) +
                      (I0c0060fe260afa3cdc72f35ffb6938ff) +
                      (Iaec1f186cb4a65da21d41e637fc628f7) +
                      (I9c15a6a5c0db11ede80ff6d04c9a56d8) +
                      (I8922487573e02d684a3d71448c3828f5) +
                      (({q0_1[10],q0_0[10]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[10],q0_0[10]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id6a9ab06d58c3a01e1fe04fcf61406fd  <=
                      (I47f17afcd5871fc3ac378316fd3d7ae9) +
                      (Ia9642d79bb50567348083b4435c7d66d) +
                      (I2b2bd845428c49346ef8e94e95b618f8) +
                      (Ib730fdb59198f23d1e590f6d6039e96a) +
                      (I644e83f0a7d432fba38ffb2d99088eca) +
                      (I97f2b15ce0a74e68d5a4438111adcb0a) +
                      (I84c88b631bed5311cb6e99e58941149e) +
                      (I45c5e6710240685bf54b73b0d7a64271) +
                      (I5827bc87b5db1801b7db16e1e61515db) +
                      (I1c85c8f73ef80a6808c6aec0c8eca8ab) +
                      (({q0_1[11],q0_0[11]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[11],q0_0[11]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I261bd53528b82128acabd405389c8d60  <=
                      (Id13c99b7f7500c8195b54627efbc4232) +
                      (I4636821315d702a677dc93113872e647) +
                      (I9c981b0614a29386ca5e8ebc06a17f15) +
                      (I4df3d4dac24877b14e6d361bafc1a800) +
                      (I913d818403024510c55b65b56a38dd89) +
                      (({q0_1[12],q0_0[12]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[12],q0_0[12]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If7fa833bf1b1438e7a5bc783ee745252  <=
                      (I57015930f5b09a6c6b030ed01dad2177) +
                      (Ib54d55a70605119e37e9898b940ff636) +
                      (If7e146da4f3bd255b8457fd6902005f6) +
                      (Ied00d87af99ae55144fdde41ebfc1357) +
                      (I7774313f1ae5a2de98855aad572b3676) +
                      (({q0_1[13],q0_0[13]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[13],q0_0[13]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibb103853fc21f8f3d466ca16557ccd3e  <=
                      (I679baea452c3c6d04c53baa88edd8eb3) +
                      (If4132b39ddb92aa02d8d0346fb0e6691) +
                      (Iba70e737d52e6812a67c159520e5192f) +
                      (Ib9ceb8315f0cd848f861bab677c2c694) +
                      (I7846bc2cc11e08d05f7c853c4920d555) +
                      (({q0_1[14],q0_0[14]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[14],q0_0[14]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I37446eb66ccfd268cb418655b8160fe1  <=
                      (I0865623d3350645e63fa6e6c9b78ac57) +
                      (I0262b30a4efa9f1cfb11d1c3940de9e7) +
                      (I7a2e79d42779ad235bca6ce3757cf588) +
                      (I09e9a3cd4c12d204f760758e873a177b) +
                      (I30b0b1d54912c1a41a02a25ab238bb54) +
                      (({q0_1[15],q0_0[15]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[15],q0_0[15]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id17f6250f8c7f1d7f75fd27f92698da3  <=
                      (I49fb0909ddf66fc0073e6400f1a07844) +
                      (I9938397dc94002481984f5b560fadc58) +
                      (I4378d139db4b710e3587aa72df22b70d) +
                      (Ifa43d74fa91b7b9884969f575ef9ca8e) +
                      (I7c19a79f441ecbb73685db5a505e7479) +
                      (({q0_1[16],q0_0[16]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[16],q0_0[16]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9957b02e8d0d888e6950eb553d9084d7  <=
                      (If2af8106efc1f7dd02c074af68278b3d) +
                      (I89a3f8d5f760d1a650f85814cbfdc017) +
                      (Ifae345c79662c3df3dff0fe68ad68746) +
                      (I88a61cf72347d695489909d0819332ab) +
                      (I9aaa036a6158d11c235bdc8406d79f4c) +
                      (({q0_1[17],q0_0[17]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[17],q0_0[17]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic71258b745437bc8463fb4f847c55e27  <=
                      (Ie8df350430970b5f1229cda772440f85) +
                      (I7d77ac9b64b2e8cae21c6e36947e3ca2) +
                      (Ic1faed76fca5a9ceb7db26c2f43623d9) +
                      (I3ca2b9b77ed8d78a10aff42a07a53b07) +
                      (I1f00849ea055a7893df386aed162a7b6) +
                      (({q0_1[18],q0_0[18]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[18],q0_0[18]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I24bb5c315eacf0f4e8c86f6582389e39  <=
                      (Iaf8a19fde3de660c3fa925593bebbe0c) +
                      (Icd1da43a4d95230e79dbd35a7ae41066) +
                      (Ice9079fb6e08d629f8c0c9ce332c8f11) +
                      (I15fafe2baba4d2f28037023a81ce0a81) +
                      (If4d5b48882e9e628cf51ad2ac2f38c22) +
                      (({q0_1[19],q0_0[19]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[19],q0_0[19]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I607f203694ff76930cfee4103cb73c30  <=
                      (Id0eef1adba01447c14a6f005782dd9a2) +
                      (I1d1a7c5928982c278d068ebd262254da) +
                      (I6354a0e638340378124e4df7f3d145b8) +
                      (I0236c912c6d684bf4862b725be9d5951) +
                      (I6f3be51d69b2b64a04e55b8946d5dd56) +
                      (Icde3e6dbcf985682041f30903ad95572) +
                      (I46ee30b46020d91707689f3468f00e26) +
                      (I2605f078c1a9006c93855a9a2b0cf6b9) +
                      (I4d226dd2f0bfcdbea6a2e6a6613c1b64) +
                      (I5c942076b173cf527e1be2ddb8560e84) +
                      (Ic95191bccb18e26c10e56be395ca6b1a) +
                      (Ia284f974dd8a526f31eb81ed71a06e94) +
                      (Icc93450a007cee4c0a42717ed7600528) +
                      (I9ec9f389d0489908d497487e44c6edcd) +
                      (({q0_1[20],q0_0[20]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[20],q0_0[20]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ica8e4c56ebb37e189ca8e6b3daafdb80  <=
                      (If8a527cc7f06a9963a80a880d225d34c) +
                      (I39ff4663007dbc89b403f3b08a69bb6c) +
                      (I9590eb28a81c730b83b92ef7653e71a1) +
                      (I2ba1acca919bddcc22a41a28d43a4e3e) +
                      (I62d8efd4227cb3dc88aa08b6585fafc8) +
                      (I749e987266a20840bb8a4b1a2a2fc5b0) +
                      (I7607af5d98e8070e3d15cee23cdf877e) +
                      (I2e11a697d7f17ac30302eadb500de72d) +
                      (Ia0886ce792e062e22d0c224158cdfb7d) +
                      (I6b3cd79aa87235ff174c0299b855dd3d) +
                      (Ie4ae993ddb776bdffec843db0def2f5c) +
                      (I3ed2da9b53daac0852a06ad1acfad21b) +
                      (Idefa29d4d4e2a6e9147f84893520096f) +
                      (Id1fbbe0594dae272856566522633bb3d) +
                      (({q0_1[21],q0_0[21]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[21],q0_0[21]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7089386c94261e0febf3b4f7dc1aec30  <=
                      (I8070a3b7d8b1a7ae90c1a2d27aed09aa) +
                      (Ie88285ce2b9c71de02ebd62e8f44ca72) +
                      (Ica1997c6c569c1d1f45224fbaa4e6b59) +
                      (Iaf08bcaaeb15bb0c971432f7f8b16d0a) +
                      (Idcb37cfc357cc088c775409fb9225b51) +
                      (Ic419255414995e7168afb97b051fa64f) +
                      (Iee6da3120d73373627b25ab7c0dedd28) +
                      (I56fc99a22960232b305d6e683c66fcc7) +
                      (I0a9a09b0ab43d2a0f1d1d01e13f0333c) +
                      (Ibc73d07e0c97a6fcae791e04106cb082) +
                      (I224bbdf94ac86c5c376d1db4f4d4e060) +
                      (I43f2b69c6b427de3095c44d4166b77cd) +
                      (I1e50c90010a3df1a8ce1cff811cc7a0c) +
                      (Ie1817cbf3a80dae435a5571dfbd2f5ad) +
                      (({q0_1[22],q0_0[22]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[22],q0_0[22]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia1e4f20f32f7371cb0078d6e80fe8b7e  <=
                      (I0052d562fb3182890c8828e52d437b11) +
                      (I1eedecb1d8ff505c75be7787199afada) +
                      (I7ef544597a185b1de63b4ffc4a1d44c2) +
                      (Iadeedf3870f0b1eae98d0f7dbbeff04a) +
                      (I70ae07db9b44d530be220f06401d3d3d) +
                      (I7992ea31927b4f0e268462a3b0f18c5d) +
                      (Iadf927d18644a232ad1f1eba7db82934) +
                      (I2a9c673cdd7ded79e09ada38c0f47e6f) +
                      (Ia86740e870d8063f0266b68ad6d7481d) +
                      (I6627bcdbaa8afb115123777abd45435b) +
                      (I96fe3eb633eff6958ac575b997460bb9) +
                      (Iefdcb71f2903b11f5cb0b8857f7a1727) +
                      (I2eb90278aaa54b9c8212b3b4af7c3617) +
                      (I43493f70f0336453d77caf7f27503daa) +
                      (({q0_1[23],q0_0[23]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[23],q0_0[23]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I790cbca796af58b1726d0a4680cc164f  <=
                      (I26a7fe395eb583258c1ac58aaaa3234a) +
                      (I21668ff77cf75570cae97f575cbcf644) +
                      (Ie48be9e6b6fd63baa104d0a6a4561a1a) +
                      (I05370777439b01811fe7f750d2f724f4) +
                      (Icdcd83341f6b5c404f91ec7e97d0550c) +
                      (Ibba4e82d1510ddc16eb4ef64893cec02) +
                      (Ifb00ae47340bc99669c71da34cccc59e) +
                      (({q0_1[24],q0_0[24]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[24],q0_0[24]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0a93f095f9efb1542116a295c0db9c8b  <=
                      (I75a4cf2948bebc58e12bb039ed273ff2) +
                      (I5a9fdec7d7ff99fe33ad6cd8afd9e059) +
                      (I47b1695a74e4d27389b97543415dcc67) +
                      (Ieb38fa62119a5a77c060d6634e051298) +
                      (I3459d98131faef5a5040a03847890b55) +
                      (Ie9b9221b2122087cd5f309570b6d31ca) +
                      (Id4451722e8e2393d627dcd0175dc9903) +
                      (({q0_1[25],q0_0[25]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[25],q0_0[25]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I989ba39f188a44475a83e65a4960d2af  <=
                      (Ic10356f9069e3651b9c045c906e63512) +
                      (Ic3a431f39c678b7175ed30fde1fa6424) +
                      (Ib01cfd833a63500e03333f263805db3d) +
                      (I0b7b4c0a8503c751229edfe0237cc903) +
                      (Iace01234164c8a9f7c98eeb83268745b) +
                      (Iace8b3b3a4c16763132b5aaa6b24212d) +
                      (I80a89644e278e96b1cd1c4b7f764dc34) +
                      (({q0_1[26],q0_0[26]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[26],q0_0[26]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9bcc1d9b3dd258fa7b6042f0185d48cb  <=
                      (Ia92d2276a8a23521ad1b88df7c27bc2e) +
                      (I39bbec42c442d1e8c818f46ad9c096a8) +
                      (I88f1b5c12759a5efb2d2ded8483c9ed2) +
                      (Iaf4ae293c576af16f5f43a8b86c1aa3d) +
                      (I68b575fcbc5321d4d26a22bcdbb506f6) +
                      (Idf600b93ee1018ecf969ed7944b6bc7b) +
                      (I1cd93172cf5996bc870063aa642188a2) +
                      (({q0_1[27],q0_0[27]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[27],q0_0[27]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9ba14715d9f33ef45681ad52f5be9593  <=
                      (I4af080cb4e5cc525db95e5f401019e8c) +
                      (I6fc8044eb226a14ff1a786ddc96d2414) +
                      (I27fd0073dbcdee599fbe85cf48806efc) +
                      (Iaee6d725a8b2653eeac6d5acb91f8f36) +
                      (I4afdeba4fc2a12a6cbe3567a519367fc) +
                      (Ib42816335dd8475dcc78662c4c0786c1) +
                      (I343c9efe71164c01e9c7d599e032864a) +
                      (I108c269ceec4adcff9afeda01101b838) +
                      (I761983331fb6e3c6c437b3f1660f0b6b) +
                      (I70d32affde22f9dcb2d77430fca39069) +
                      (Ic08e85346f61da036a15345a13ac12f0) +
                      (If5dfdadb3868ed5a495007362f7db648) +
                      (Ia1ee5579358b564de06c08ca418a9bf4) +
                      (({q0_1[28],q0_0[28]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[28],q0_0[28]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I396a897f79b519f4fa02af39d0274f64  <=
                      (I9bb81dda8102b829441be46460eb8900) +
                      (I8eef6ca0a61a21882ea28b3d63735228) +
                      (I438522d92cce6f7010246424746ca255) +
                      (I92496f68b44a94565af28a2c28d6fbae) +
                      (I66528f43f614f0edb715564eba3c77c1) +
                      (I8cab9fba615b94fd4bb6934325be8ab8) +
                      (I92d9fec22d36b1baac8bd78abfc1bbd5) +
                      (I4eadce87f47df6d8f0e4acd057de5a09) +
                      (I73203143fe37933c16fff873c1abf512) +
                      (Ibed2a63af723a7abf96dacf1951e5266) +
                      (Id667c80003b5541de9f84d3b8709c828) +
                      (I02cbb4255db2b21ea32140f9e9ddb36b) +
                      (I65354f2069de0c25bbe7cd50fbe892aa) +
                      (({q0_1[29],q0_0[29]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[29],q0_0[29]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I197c0cd576e16ee2197a28c86397f801  <=
                      (Ic279867ebf3055980f3d813d5dc8dec6) +
                      (I5c05da8a222ad5effb9815cbf3ec25f3) +
                      (Ib8bf21f32c0e8b9cfa42a53807bfe3a3) +
                      (I7208256bb198bfce1be71390b01bc028) +
                      (I49f2a06ceb3a59773c65b19f54ff362b) +
                      (I86e495dc894d2aace15c1aff89798bf7) +
                      (I0d53bb5344cabe5fa5ce3ecf7122a260) +
                      (Ib2f5f5fc77ea8b529f2471c54388f2d1) +
                      (Idcada1bfb3c0d1f2a09aab58a2071a57) +
                      (I814b62120953991f9da055f118967e05) +
                      (I123a212546a8ac394051425db4924812) +
                      (Ie95f1a7e0effcec0aa423dc803056a13) +
                      (I106deaff50b8480eac31ddbae2ec7c61) +
                      (({q0_1[30],q0_0[30]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[30],q0_0[30]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I094a178e55425f27ac1ff6195217396b  <=
                      (I68528be9951f5b8805411711cd11ea59) +
                      (I0f034a8f077b0ab231727b6298e366d8) +
                      (If9c12f8662333fb54a45cfa1bc5da487) +
                      (Ie1681d905517daafcc7584725cd6014c) +
                      (I2ff3edcdb6158f1e3c9a555aeefc0850) +
                      (I43b380be6df7df0d354223d0a0d6d6b6) +
                      (I23eb1dc4d1c992f804dd04a2d823c778) +
                      (I7f90f96c0260560ad5e6dc7448b2670a) +
                      (I07b417cdcc99eaea3413f563e26ddc73) +
                      (I2f3ab9654e515a54e22e73d6c130ccc3) +
                      (Iebdc41368d57498a04fa73e30b10a966) +
                      (I5b4305bef5b4350c1d7ae143667afddd) +
                      (I2795d21d343b83a69146314a2407cfa2) +
                      (({q0_1[31],q0_0[31]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[31],q0_0[31]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3177408f7d08b431be99297fb10586e6  <=
                      (Ic6386d7d8813731d612e24b715740275) +
                      (I4c366a57920ff090a98a2cb8b9caa00b) +
                      (I14cf5d43fc9864820a8a25efcc5c6d86) +
                      (I33b99994abbb5ecf8eed4de39033e4f8) +
                      (I7c3291f0250d13ca94802b0b071a95c6) +
                      (I2c926fd9d306e9ae13364e07c4b0395b) +
                      (({q0_1[32],q0_0[32]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[32],q0_0[32]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id4948c876d48bdbf317d32f135e645b4  <=
                      (Ib23edc35fa5bbfe0415fcf0861a22d9b) +
                      (I3e0e682047f7cc36142e668828cbff1e) +
                      (I99fb9030e8361e57818c07511479a9b8) +
                      (Ic87c3d7762a18772972552162e1d1a8c) +
                      (I7e393e6c1d1bc44daaab120d55f5dd59) +
                      (I448f126fd3932d5065abbe7bb2d92c56) +
                      (({q0_1[33],q0_0[33]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[33],q0_0[33]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ice5ff01d4fb4583898498651a0ac0171  <=
                      (Ifc8c6df8904b97674f2970ebc95b523c) +
                      (Icd0622a90782b9c451950e7ab0399567) +
                      (I6493b3c087d4685a6b3f98c73dc2ff49) +
                      (I20c2057240417146df144b518b43d052) +
                      (Ied029d0bdea3bf134744c99426fa72dc) +
                      (Icb82c9ff4cb58159a1c3115c6fdd5f8c) +
                      (({q0_1[34],q0_0[34]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[34],q0_0[34]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0fb33a5ced3d15622c9aefa188052e24  <=
                      (Ia3450e134e4086c35acbdee1e6042396) +
                      (I5a0f27df5158309f32f0df31e8ae3ae3) +
                      (I17d9e19854cef197fd3267618617efc3) +
                      (I2993acb61f1abe529f8a60c94a438550) +
                      (Ic8be2c94235fb40f78da33179ce4873a) +
                      (Ib3367565e4456da15e7c2315dccdb5e4) +
                      (({q0_1[35],q0_0[35]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[35],q0_0[35]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0074e1c3ca0ff903a9201ac5fe7ca841  <=
                      (I15a1671def323cd294591564ae6ef8b1) +
                      (Ic512effb493a06ece58a2af155135004) +
                      (I2c72248cbe49ec0a0febac2437b8a6dc) +
                      (I964e17c41a134c080e9c43412a514f3f) +
                      (I94f1724740defe5bb7e40041d0e266a0) +
                      (Ic19486b6ab0373b9c0ad8f7597782d8f) +
                      (I31243de90dc2a1656ca9d5e03bdd78da) +
                      (I242a30bdc8699d8ff550b25dd53d6c59) +
                      (({q0_1[36],q0_0[36]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[36],q0_0[36]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If65f587e987a51c093e8dd4df532e26c  <=
                      (I9d15f76bb68b214057566cba4b511214) +
                      (I9cc16a00912e7dfc05fb505a9db23cd8) +
                      (Iacf9640cbf486411d6ceb8fe1a2fd5c9) +
                      (I9015033ab0caf3fa41dae4de43f24a82) +
                      (Ia630e59cbce82a570ae3890a6c0221e5) +
                      (I4904ab14b19fa1b6befc218bc7be3842) +
                      (I282d2eb4e74e034694e33273b9cb19d5) +
                      (I3f33901c407a87e10d86c13c83dd52eb) +
                      (({q0_1[37],q0_0[37]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[37],q0_0[37]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I33d7e77d08590f0dfb1867e741dd8b6b  <=
                      (I43f41bf07836cee48069e9890c1de2a0) +
                      (Id88480a0a350bb5fcf01ed5fff0bbd4c) +
                      (I1d9b9ff357667a362f0442f19986f451) +
                      (Ice73589836da9028def6efb24a04dbbd) +
                      (Idb72c046c5996fbbd80b706666ffbd92) +
                      (Ie5757e7b1647ab7d43cdbcf98cbb77fc) +
                      (I6072331f838d82329a07a4ffa340c7b6) +
                      (Idf6875955525d80dc660ce956f4a84e7) +
                      (({q0_1[38],q0_0[38]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[38],q0_0[38]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I678c22563e0273403b046df4261f21cf  <=
                      (Ia96955d9c0a8a587e0afab37c8415d8c) +
                      (Ifec374bce7f5507438f550df22d61a01) +
                      (Ief67e897e57b96e2ec200e82bbc7caeb) +
                      (Ide604e9bbe35cb55892a4602e18b2527) +
                      (I262f2390e77ec486ccd3a6ed05816e2d) +
                      (I280e20c20c0b4f26278b3de9b2ff84e4) +
                      (Ib3a0307176d424a4733720416d71069d) +
                      (I76060709de3ea188748849f043c59ac0) +
                      (({q0_1[39],q0_0[39]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[39],q0_0[39]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Icca700c12ae2e8155ca6b41e692e8a8c  <=
                      (I8be20605d26d218911e80a883a90d085) +
                      (Ieafa9d74d4a61d28ac4a913db460bf33) +
                      (I6fd1b4395af175eff85b3bfeef4c329b) +
                      (I39e6d3fb468aa40ea73535e81556ea65) +
                      (Iae449b74e50e0907feae9e60f2329426) +
                      (Iebf769a6bdaf214c1006c55c608d4eda) +
                      (Ia030c08757123aae947f86ab8bfb6d94) +
                      (I8c35c5b343b552c22000e194c517ca12) +
                      (Ibf80bb564263ea85bd886a8617f09bb2) +
                      (({q0_1[40],q0_0[40]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[40],q0_0[40]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5ed74e81d2497681af5a0ca13fe23088  <=
                      (Ib8dfd9b8badef282ca00a4f793c3c868) +
                      (I596ad7e132f272cb196b74faa8c75aa4) +
                      (Idc629414f6d0236ce0714cfaae23f065) +
                      (I157fdf8775206858c08682db3039b084) +
                      (Iacbb4daf5ce5c7eb1a2afe30d0cb5382) +
                      (I4e08021c0235fafb60200aab97827a8f) +
                      (I730634ea15ac94d241f3ad2d6393a227) +
                      (Iee367c535d9c39f872d2ec043e7e7b33) +
                      (I68bb1f26f878862f288c1f57049cf58b) +
                      (({q0_1[41],q0_0[41]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[41],q0_0[41]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f  <=
                      (Ia9b5d9ede006c56a6d83905529c77b7b) +
                      (I1487170cb1f3370ad45efc801cefc8ab) +
                      (Id88568dd34fbee42c9cb8cc15ac5c31d) +
                      (Ia30539545e66c4cfc16828140149180a) +
                      (Icbfbb37bad6344005dd233b3605a784f) +
                      (I91a6408a11fab36a8ba3dbd3f895a803) +
                      (I47b878f27c30f79a37e97e022307e9e9) +
                      (Ie76b0739aec66f8860870e66e87a6445) +
                      (I50383e3d7c172eedfa00aa50a9faac4c) +
                      (({q0_1[42],q0_0[42]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[42],q0_0[42]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I26010e26e22d8a2ea831e86fae34a24e  <=
                      (Ifeaa99e03bda8ded058f98387de3d49d) +
                      (I4255ac1af4367c321567c4e46b06ab25) +
                      (Ia445bdc7def7d8c1eec31ab892c25c41) +
                      (Ic3b4752136ac08e343933ccc3a4ec47c) +
                      (Ica6707efd6d44ba6bbb87c0593a3d828) +
                      (I739267bcc50c54b8a685cb3c6afc5cc1) +
                      (I9160d11439c5140c0109b5190eb82e6b) +
                      (I6ff7b86cd7f63f9243646f1be10b2577) +
                      (I165653ab165cfafe2b74cd441331f9e1) +
                      (({q0_1[43],q0_0[43]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[43],q0_0[43]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I578efe5c2c504f12c8f2466a7f734215  <=
                      (I08a8cd6965c23af6650568b654831b20) +
                      (I9b6a674dbcbfcf65f1ae0deb8fc3566d) +
                      (Ie3a336de822ac7baf8486b1618ef1126) +
                      (I5fc3c26d6c5aa893dfd5caa0f677233a) +
                      (Ie22b94121b58f17af14c75bfb27f96dd) +
                      (I0d9f8c99194d9d6e187b4ad02fcce8b4) +
                      (I71e101962e766a4d1484b3235359a4b5) +
                      (If2539da6722562bbf31786fd0036666a) +
                      (I22c8ccd4a9018ad1c129aa058bf579d8) +
                      (I83330fef69470d2f5def8e6d7d9c50d2) +
                      (I0539d598bbe3d50940329a282c801328) +
                      (I202f88fdc946494d55fc8831c2e8a34c) +
                      (I3ee10f6a7785a236db317515fdd23a2d) +
                      (I453fdf4fbb5af5bd28a20d7643da9eb2) +
                      (Ic4a6c02880a9aead7353332708e3f388) +
                      (I7fb3b66cb48521f8715f66bf5642cdb2) +
                      (({q0_1[44],q0_0[44]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[44],q0_0[44]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ida86d05f907d23ff9fed06927c2ec9d9  <=
                      (I2fd872df07f50688486c0d602cfc5549) +
                      (Iccefa45795486757515d95e5908b306a) +
                      (Ib1357cb20f471f1670ac2448f964f8eb) +
                      (Iab953a8974a1eb619dc0f074c003b5f9) +
                      (I6e37582849c2c98fd15ad92d22c222da) +
                      (If004de0cac6e5f7701a1fce48c6936d5) +
                      (Ic1efa395cc1fd2c5a1d1559fb169a5a0) +
                      (I8e96c69e7d872be23229353808c34953) +
                      (Ib6aded6c73a8cc3cb964b0ae895b859e) +
                      (I939368b76d98b43826c68c7f468a5632) +
                      (I544f6263f16cd5e0b7cf28c511a8f6e3) +
                      (I484545c4d2c869d79eb17f51e11070a3) +
                      (I39289e6385a9bc378a9b8dd440249a7f) +
                      (Ie9cce5746a83479a567bbaeac6dbf497) +
                      (Ic044d7419cc43736d278c2df33b4a3cc) +
                      (I6714551e8885ef5e4490673fe1b2dad1) +
                      (({q0_1[45],q0_0[45]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[45],q0_0[45]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9d9f8c7a23d9750ec44e706bf763df76  <=
                      (Ie9ab3c88ac62369e3d92d110165a94a8) +
                      (If38feb4f76f761dce6145731ad235d7f) +
                      (I6359856a1843d8c8b65dc478bccb3acd) +
                      (If6f3d91c3c7a43622b9a522492cd83d3) +
                      (Id023a6298e65da1f4da3831f5136afc2) +
                      (I6b24690f394792edb0d82b3b9e110851) +
                      (I5b55c285f7e3e78447fee68532ab9f7f) +
                      (I32701d9e4b96853c53f0ab651a6a4ba2) +
                      (I82f266e5792cdb6e7ebd264e246161f5) +
                      (Ibfacfe5b83819afe7fbd4bffa2d6d4e2) +
                      (Ib8e68a77ad8b9e7cf415bee17645c3f9) +
                      (I644ee0055a55f54ab3544bb532e39c61) +
                      (Ic5467e42aa377c6ffd8f70673808774f) +
                      (Ic57eb4a034247a4c952d8224ea9f2bac) +
                      (Ia642db613c0ec1ca4e69afde7a14a839) +
                      (I432aa7cb844286c442356954f8814260) +
                      (({q0_1[46],q0_0[46]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[46],q0_0[46]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0b41b002a32b8e9e2fe68e819f228fb7  <=
                      (If520c1cd27f9d4bc52d0d029f693b660) +
                      (Ie87075ac979410cc11099a356966b8a2) +
                      (I6fab46b1766878b26b53f352fee98223) +
                      (Ieaf14683f40374c4531326d228cb43c3) +
                      (I5149125aaaad943d891df6a3c2be93a0) +
                      (I770dff588ee1f52f58bea1921cb23383) +
                      (I8f0a90e761111a613d2488285534a500) +
                      (I765a8825e42180a6c63f7b33703bb483) +
                      (I512cc8f6519aa08aee18225b56d47c9f) +
                      (If08370fd0e8af818c6db20f43e74034d) +
                      (I0ff382edfc8051459657ffa3899f5f73) +
                      (I9d2864024148337277523ef7fa2e1600) +
                      (I1c85a2d1df6749a194072eb731506bfe) +
                      (I3e3ce8b4ead150a6eae2e5c701c7b598) +
                      (I45bc13ae0e0554a79c62cd9c6aa8f2a5) +
                      (I92678f5b52c9c55556ff7f17f0f607b7) +
                      (({q0_1[47],q0_0[47]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[47],q0_0[47]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0e872d4c07169cac84549178fa144274  <=
                      (Ib4bdc9069d0c08655f5e87f705943eda) +
                      (Idbf9094c94c931f16fba468b9dd59a25) +
                      (I1c3c4ce44610e04c5eef2fcbc2ea5114) +
                      (Ie84be0ae8311d906eff08f7f5b214943) +
                      (Ic90b98708faa8c8b75d4bd9a52c292f7) +
                      (I8eba6f14f42701d22859fbea94bd1871) +
                      (I6d83efa9f988328f487e9232bf2633a2) +
                      (Ic23e01562c8a753fd70c343297be288a) +
                      (I5669856f88f5e2c98f64df696db76414) +
                      (({q0_1[48],q0_0[48]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[48],q0_0[48]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6f4ef0f404ae046519b8436171d51e09  <=
                      (Ic3a608b850709286ea0ad2f67425d9ac) +
                      (I5267fa34449e6eebe891017fc32d0749) +
                      (I599d01cfe6e54d8e45d64446c446818d) +
                      (I8f94dbafaac589ac9f14b56d4556ff96) +
                      (I754563caea429d3d0e22df5d193b84eb) +
                      (If7f373506cac70f8ba1222db135c27e8) +
                      (I69f563e7b7ad483893ac9c4684349769) +
                      (Ia0a02781c674fe5d769206448d475245) +
                      (I1b7a401bc11741e6f011fb9895b5c797) +
                      (({q0_1[49],q0_0[49]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[49],q0_0[49]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4d04e66ad9103a685fbe088b74517452  <=
                      (Ieb528d666fdb708279184bb59eac25d9) +
                      (Ic3ff7ce12c836bf0693252b9a7a7cfe8) +
                      (I19bba6a58ad3ef959b33701f82761984) +
                      (I8acc93b34974c1e708b0e1591f7b2d3d) +
                      (Ib60d4ac0fcadcdfce5a14fb92f58423f) +
                      (I039f05d5be891a37e04556f1eae674d2) +
                      (Id0f75e19b94541ed5c5c352d13390d2d) +
                      (Ife1190f76c2e251704c2960c23330a48) +
                      (Id3e0c98bff2636e216b4d3a0ffd51054) +
                      (({q0_1[50],q0_0[50]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[50],q0_0[50]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I988e525020c1e43d238fad41dab4e6ea  <=
                      (If4d3b31b87c0f723241d35ce7e854eba) +
                      (I72369dedfe36cb22269033cc305b730c) +
                      (Iec71fe7fcebccf1ae0d10a5d187fcc44) +
                      (Ie11da10808c4ca84f399535df6261307) +
                      (I280fa9d114e227cd649bf0e55e845651) +
                      (I94c4e11670b4233fa072517a8f19c901) +
                      (I4dca2dd40a7127ce44f83b430a34c738) +
                      (I1a24e98165afa62bd14986911a36fb6e) +
                      (Ife1164cad7cda4aa9a08d94dfe86add6) +
                      (({q0_1[51],q0_0[51]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[51],q0_0[51]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I90d92887cb2526a2956d5e8c9fad760c  <=
                      (I8d8d95ff26f33f69a182b32ccde23905) +
                      (I2508854bcbab37bd09c9465c377c06aa) +
                      (I140078292f7209eccacd53a8bab18016) +
                      (I141fb1cbe09f9abe282cffd4de815d25) +
                      (If79d1d378f7c6fd29fc3335ec5f5c51d) +
                      (I4a41999cea9357a85c73a0af509eeac9) +
                      (I8e517c401d62dbb10dcc96ab536f6afb) +
                      (I8ad3627f171eadcc960a688ac0afcbc0) +
                      (I85c4d3d6c8408c6f38741257ed177ca6) +
                      (Id66c47fd69c175a4393e975a269cf053) +
                      (I37dca40506d61bdeab1255ed4892ca20) +
                      (I340c98b886123c541a1b8d9fc8a6d48c) +
                      (({q0_1[52],q0_0[52]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[52],q0_0[52]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I00fe3792cde1eeab36e576fd6634c4fa  <=
                      (I2dc64c3b06588542b027f997437bee63) +
                      (Id92a37c091100e9df08e24498ecb4022) +
                      (I74a4b9365391fd20c34588002ad40547) +
                      (I461195b7ae78743e09ee50486ad6ebe5) +
                      (I356d747600182675699a2d2634d4c5ce) +
                      (I87d6a5d30c3e4202cf51f33c7a770c51) +
                      (I960768a84aec9d5b8bc7c1c523024a25) +
                      (I09b5273bb15d48a7fd78559930fa6d1c) +
                      (I5814a85c45fd0f7be21ed325235fe4b7) +
                      (Ib06b60cf9933dd8952206c5f3ccced8e) +
                      (I67347c413b5efd8ff9e0d5bc7ab2a047) +
                      (I72b1bb104bf2843f161448baf7aab44b) +
                      (({q0_1[53],q0_0[53]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[53],q0_0[53]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6e586c5ac59a28b30c377e51287bf04d  <=
                      (Ib23d889edb5a6d9f27de977d3b1a2616) +
                      (Ifaff9dd032cf96487be819c59b03000a) +
                      (I028ce03be0618b816e0ecdf43d4cd6e6) +
                      (I6ae2523095237282533e0b5f1c26b488) +
                      (I5aba6218461e8d571be03a3ef041ebaa) +
                      (I6ca8a1fa2c72b1c61d11dc7d1ba5f37b) +
                      (I3ec5819176ad4b0895a9118d90ab22b5) +
                      (I49b64469d298012dbb131d879bff38d6) +
                      (I95361d5f524ccb9feb42811af5c482e2) +
                      (I9c4b34b5fb1d59c132bcaeb6258675df) +
                      (I613d4b1e3b9e812b785c9cf14fefdfe6) +
                      (I848ed394bd4f0b199d11c0ff458394a7) +
                      (({q0_1[54],q0_0[54]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[54],q0_0[54]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib5dc74106d8841d25a793010fdac599a  <=
                      (Ie65a0634454381e24bb3223a333e3ad0) +
                      (Iad166146f7df5e8068fc6efe4d3e4141) +
                      (I63e45abd4d27219bddcef06108b72021) +
                      (Id1bacd13718f7c29c26b63c239d04dd8) +
                      (Ia3104c69fb4f7abfb5efa3874169a7ad) +
                      (Ie1b7257c99831ec5864f65958ecf14fb) +
                      (I4accbad1b451ed2b622e15ef9ae16d13) +
                      (I5ce8b2f633011e89356243a1a71edeb6) +
                      (I3e5139f24e3d082eb31b0e61ea9fa1aa) +
                      (I61cc8a0f49e393721a62a776e4793deb) +
                      (Ie631e40caade823a196370fc3358f042) +
                      (I4c971e714427664c59c6371e14781bae) +
                      (({q0_1[55],q0_0[55]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[55],q0_0[55]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3eaf142d2734d2d0decef084dc037b50  <=
                      (I36ca732e811d67cd742d24fd4cae887b) +
                      (({q0_1[56],q0_0[56]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[56],q0_0[56]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2d171ad83e27a3745d204849a6f46954  <=
                      (I354fdd241d5d07f0d8380fe8924e0a8c) +
                      (({q0_1[57],q0_0[57]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[57],q0_0[57]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I977f1083f5e4f6f8ac38e2c5aecf1b79  <=
                      (Id38b705f5d2863a020a475ffffc8afd6) +
                      (({q0_1[58],q0_0[58]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[58],q0_0[58]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I9bcd673a4293e14fd20b48fa20492df7  <=
                      (Id6e5d67e7bb7c4b999459374ea80459a) +
                      (({q0_1[59],q0_0[59]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[59],q0_0[59]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Icb7422ea46b22b9330c123b40fe343fe  <=
                      (I05341013abd4206eb66fcddfd63bfe26) +
                      (({q0_1[60],q0_0[60]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[60],q0_0[60]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic414cdba230d7ea73972b0eda1ec6b1b  <=
                      (I15da71a21f5842cb65b543d9bc3e267b) +
                      (({q0_1[61],q0_0[61]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[61],q0_0[61]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie4e1e00503dba189b0f871c3c0810d76  <=
                      (Iccf255fb3422c558465e45226068a16d) +
                      (({q0_1[62],q0_0[62]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[62],q0_0[62]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I721c43ab62b42a18c3f5228fc0a73262  <=
                      (I1c2674b2e6b269ed539827412c5199a5) +
                      (({q0_1[63],q0_0[63]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[63],q0_0[63]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1f7cb03cf806b247be1cace4d75de942  <=
                      (I6a3f405bb4a0c4448d9b9d3dd95d036c) +
                      (({q0_1[64],q0_0[64]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[64],q0_0[64]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I775cc766b069022bc00220050feee4e4  <=
                      (Ib528bb7a64cce4f694081d151fa6fa86) +
                      (({q0_1[65],q0_0[65]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[65],q0_0[65]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I08b78f774ed494fa7f119977bd92679e  <=
                      (Iaa40bd3abf668a21e0f87c7bda7b3f69) +
                      (({q0_1[66],q0_0[66]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[66],q0_0[66]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic7dc7f94af108ca7c8003a2d07e1e168  <=
                      (I919d36a7f6ad42c4bbc23222beb73106) +
                      (({q0_1[67],q0_0[67]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[67],q0_0[67]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibe1327961152cc2d26b3f19476a6e2c9  <=
                      (I648d2a279dd1f587b1e45eeb35f2fa90) +
                      (({q0_1[68],q0_0[68]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[68],q0_0[68]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5ba97de444af4e8c9744c3b707502edc  <=
                      (I194a64bef92ecf6714141eaa5d41c9d4) +
                      (({q0_1[69],q0_0[69]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[69],q0_0[69]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3e4f1314042010b5d7384693b580da7b  <=
                      (Id332e7f482524adeac7f7cdafcf5ca46) +
                      (({q0_1[70],q0_0[70]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[70],q0_0[70]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4a47ce6e21c1a274578397e480c184c9  <=
                      (I226383d68f89db716cfd8d08b837865a) +
                      (({q0_1[71],q0_0[71]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[71],q0_0[71]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id184731beb200ad6a53ce273b963bb3e  <=
                      (I2bdf5d319ba9089a4da34b108f5c5ae5) +
                      (({q0_1[72],q0_0[72]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[72],q0_0[72]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3317f2f6eef9a8ef1fe1ff68b47c5d03  <=
                      (Ia91800792941ec7cc60415c3f844e4ed) +
                      (({q0_1[73],q0_0[73]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[73],q0_0[73]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia6b9fa10c79e6f3847f89b35afb4cc59  <=
                      (Id7c507d96098ee7a955af8a48ee5d72a) +
                      (({q0_1[74],q0_0[74]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[74],q0_0[74]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I91e98b804ef82eea53c5e8eccfec827f  <=
                      (Ie15e4c1bcdb0e18085d4b320ac6a925c) +
                      (({q0_1[75],q0_0[75]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[75],q0_0[75]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5f1e0d0c6b50f70a6f5584124e095501  <=
                      (I5485d9edcafc6202f6e5f0969979802f) +
                      (({q0_1[76],q0_0[76]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[76],q0_0[76]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id61fcc605b4b581f5d42024c2610c8b7  <=
                      (I7fe364f9f537cbef782e7007848a1c10) +
                      (({q0_1[77],q0_0[77]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[77],q0_0[77]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id64738b7668931553151dbadd5605b71  <=
                      (I52dcf5bace9cadcf8a895aaa6a8c1da8) +
                      (({q0_1[78],q0_0[78]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[78],q0_0[78]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3bdfb451eb96d256da542864d39024df  <=
                      (I13a9eec6175e695ab8bc4516cf57d6ec) +
                      (({q0_1[79],q0_0[79]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[79],q0_0[79]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia740d8ccd8230b28d078b2ea3e58d6ba  <=
                      (Iee73a7c685a4cee03f33d3ef379b1c8a) +
                      (({q0_1[80],q0_0[80]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[80],q0_0[80]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I574050722f82569d34bc2cfae1eedaa9  <=
                      (I740dc91716e3906ad078e2c7cc3c925a) +
                      (({q0_1[81],q0_0[81]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[81],q0_0[81]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic8f7ec6ee09fb9ee2467e3cea30a44a3  <=
                      (I514d2dc697e9b39ba027c418a6df6cb9) +
                      (({q0_1[82],q0_0[82]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[82],q0_0[82]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2b77d922a74fdcef0d57debc789bd539  <=
                      (I782726e317a2aada9e755bcbc4b0d3fa) +
                      (({q0_1[83],q0_0[83]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[83],q0_0[83]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia1d8127af4944b23475bd7deac91d60e  <=
                      (I11eb26cf0f0b3a334e8f7317bf8d9eb0) +
                      (({q0_1[84],q0_0[84]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[84],q0_0[84]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I247abcede9914633c0a33fc402bf58ae  <=
                      (I26cb63ba20245b2c332b09e25c4409aa) +
                      (({q0_1[85],q0_0[85]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[85],q0_0[85]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1f413d3e081c6aea012b122fc94f73d5  <=
                      (Idd7691d31f8d0c09ee988116d574ec59) +
                      (({q0_1[86],q0_0[86]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[86],q0_0[86]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1b812fb764d3b48511c0d15a7efaea29  <=
                      (Iecc02842a2d2b9b9e8187f2d39e62e05) +
                      (({q0_1[87],q0_0[87]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[87],q0_0[87]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I88882bd8a9f8718411564221ad85b223  <=
                      (I5551342f1751fc64f32744a46b9649be) +
                      (({q0_1[88],q0_0[88]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[88],q0_0[88]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I232f24e2798488ee66003f3b8cc294c0  <=
                      (Iff7c29299f005c1cd5a16b64601e727e) +
                      (({q0_1[89],q0_0[89]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[89],q0_0[89]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I856284e951773518eb6c4232ea7f3d40  <=
                      (I17a5446e942bcc1dc2c96930e0a87a70) +
                      (({q0_1[90],q0_0[90]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[90],q0_0[90]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I82cbeaf5b3e4796b2aaf33dcbd119f4f  <=
                      (I719b67f84e07e90dfd29a8cd5d94cf39) +
                      (({q0_1[91],q0_0[91]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[91],q0_0[91]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iaa7791bbc193412e5fe25000ceec23d6  <=
                      (I2c835dfb3596b8bf057a7cc21122c81f) +
                      (({q0_1[92],q0_0[92]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[92],q0_0[92]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I44bdc0baed3d51ef54ce2728618ad339  <=
                      (Ib71b3d357c98dcdfae5c777ca3082275) +
                      (({q0_1[93],q0_0[93]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[93],q0_0[93]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib6bc7e75ce750a26113cbb8895c2f024  <=
                      (I086bf19f620c8a8f6888e775cb1ed7f4) +
                      (({q0_1[94],q0_0[94]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[94],q0_0[94]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib4188380f7e96d5afb99f5045674193d  <=
                      (I802c554d5b04af6b949677819a4966ed) +
                      (({q0_1[95],q0_0[95]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[95],q0_0[95]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5bba219c5024301e420e9a5acbdc5845  <=
                      (Iceefb06cb3715e1b41e6f7d89420e5ba) +
                      (({q0_1[96],q0_0[96]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[96],q0_0[96]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1bb52988c9ba03e16b1b69335d3d7e7c  <=
                      (I56948bc48c0220893d68004615a6ebaa) +
                      (({q0_1[97],q0_0[97]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[97],q0_0[97]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1b9990aaeae716f66b0f89fb02be0a74  <=
                      (Iec1368f034655d61354ab5b5e94d7d89) +
                      (({q0_1[98],q0_0[98]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[98],q0_0[98]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iceec2cf6aba9138648a3340390f39fe9  <=
                      (I1e43c0aeeb8a2461d208eba24967af30) +
                      (({q0_1[99],q0_0[99]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[99],q0_0[99]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iad7842f3d4672f42c1064c28d4c8ec4e  <=
                      (Ia6eb85b127cf9c1a437611556296b967) +
                      (({q0_1[100],q0_0[100]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[100],q0_0[100]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie5a53cf9343fdcdb5788667c45fadc83  <=
                      (Ieba89aa901e61218074af53a2484a74b) +
                      (({q0_1[101],q0_0[101]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[101],q0_0[101]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I30e06d190906bc9eb6f1c3156c47f9f1  <=
                      (I8b3b875c6c07bd97ba598a5139156fa4) +
                      (({q0_1[102],q0_0[102]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[102],q0_0[102]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ieaaaced47e22029ad2945eac9cc45e6c  <=
                      (I7b33ddad346077928620344542b9481e) +
                      (({q0_1[103],q0_0[103]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[103],q0_0[103]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I08dc6f8e837b1f6b80bd3fc742290dab  <=
                      (I11d967a5c5d14c88b5587d4cfed1d05f) +
                      (({q0_1[104],q0_0[104]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[104],q0_0[104]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I8eb6a9c907c5909dad6cda98022d70b8  <=
                      (I27458d76b3ac6520fb379405c6b2956f) +
                      (({q0_1[105],q0_0[105]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[105],q0_0[105]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia5067b1b458af82c3c2cd50653099854  <=
                      (I2525111a2fb5f10d64bbd16e148653b8) +
                      (({q0_1[106],q0_0[106]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[106],q0_0[106]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I198c6753cf12d423c709d1512e66fa9b  <=
                      (I7b7cbcd1c6d2a2eeaaff474536a69eed) +
                      (({q0_1[107],q0_0[107]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[107],q0_0[107]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib600dd8a39fda48d28e1289d44d49a84  <=
                      (Id2a7f0781d18dccc7c4e0b383b7cddfa) +
                      (({q0_1[108],q0_0[108]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[108],q0_0[108]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iabf09191227584c76d7fbc634b706d12  <=
                      (If8bc141d98ebe1be7fa81cde5c65868e) +
                      (({q0_1[109],q0_0[109]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[109],q0_0[109]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4869ba08cab90a6dcbc454b0001a7a20  <=
                      (I8645e1326c66f5efef4b9c923599d1a3) +
                      (({q0_1[110],q0_0[110]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[110],q0_0[110]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If97974406672507f8c9a1c507c4b6951  <=
                      (I0426ef66185128dd1ef4dbb68dcda585) +
                      (({q0_1[111],q0_0[111]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[111],q0_0[111]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4210341f99ac7cb08245137999739114  <=
                      (Iddd954df5bae9b4240e0512f746669a9) +
                      (({q0_1[112],q0_0[112]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[112],q0_0[112]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic24f4dbd99c8f4d88c8450d4fef762b8  <=
                      (I29e940970d87e8e09b26ab1b0b8f2286) +
                      (({q0_1[113],q0_0[113]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[113],q0_0[113]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I68dffa1a13eb6ab54615347729c1d6af  <=
                      (I488f6d9676aa85a55d030bf12e8997a7) +
                      (({q0_1[114],q0_0[114]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[114],q0_0[114]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I10153d5548b184b9ac2cecdba4ec4b1a  <=
                      (I99d761b75ade1fb2e8afbb1a77752609) +
                      (({q0_1[115],q0_0[115]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[115],q0_0[115]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I104b7f0512440cffc0fcce25e477f537  <=
                      (Iac4e3d20178049f9c59abf374752dccc) +
                      (({q0_1[116],q0_0[116]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[116],q0_0[116]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I18b6758319272eebbe76e1eee5ae55b2  <=
                      (I618d33f26badabfa578908903a613bce) +
                      (({q0_1[117],q0_0[117]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[117],q0_0[117]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I780263b10b98f9bb0eaf66c045d8d37c  <=
                      (I822d7973afe090b2764335f1b72dfd0e) +
                      (({q0_1[118],q0_0[118]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[118],q0_0[118]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I37b772442e55cbcd44ba892a0608d662  <=
                      (I12c1035353e553b3b6a13bb174ce6020) +
                      (({q0_1[119],q0_0[119]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[119],q0_0[119]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0ac256a6659ff5c6673fd110a8bf578f  <=
                      (Ia6d61947d36fc128c689808c82db80f6) +
                      (({q0_1[120],q0_0[120]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[120],q0_0[120]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If134e1d27e736005e5a390e7a2ea1f4b  <=
                      (Ie9b042f686381739b9ff219041f1e0ce) +
                      (({q0_1[121],q0_0[121]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[121],q0_0[121]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7b37b8f908cd82683832536e02faab0d  <=
                      (I0c4268c01aed70ce4fc71531bf4bb862) +
                      (({q0_1[122],q0_0[122]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[122],q0_0[122]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I08b4bf60c9c7e7229bd1952cc88bc7b3  <=
                      (Ia34e42f8de91fa4861b0c6cac5dcfc29) +
                      (({q0_1[123],q0_0[123]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[123],q0_0[123]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I267d637eb63fef9f4723f7978fad88f0  <=
                      (Ib7c5850b4f7cc77be2048d114a2128d9) +
                      (({q0_1[124],q0_0[124]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[124],q0_0[124]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4fb56a70e5ffa71f58f715da36368e04  <=
                      (I32bb50faa2b246b2d3b462a79be597c5) +
                      (({q0_1[125],q0_0[125]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[125],q0_0[125]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5e9e2acb258baf96ac4b525bba54a462  <=
                      (Idc6d40a49f05c5422758cee50f787eb1) +
                      (({q0_1[126],q0_0[126]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[126],q0_0[126]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic40f61443a4d8f87769067fc39381cb3  <=
                      (Ide1d7dc22a4b271ef764df14ac22366a) +
                      (({q0_1[127],q0_0[127]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[127],q0_0[127]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ieb36710c9a3726f33407436d62639c8d  <=
                      (I7ace6778ac86b3e05939a3fcc716136f) +
                      (({q0_1[128],q0_0[128]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[128],q0_0[128]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic804af393da2e4b9c8ef25d4a3b4e8d5  <=
                      (I044e01e8d2df46e03f00a0af2beb0bf5) +
                      (({q0_1[129],q0_0[129]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[129],q0_0[129]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I52e4c446693c29a42bb3b665f72d382d  <=
                      (I45a7ddcda2662e36b7617dfe64514346) +
                      (({q0_1[130],q0_0[130]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[130],q0_0[130]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Idbf02cf10add496d30fa44bbb18458c6  <=
                      (Idada779a1ac7b844867571d77054b657) +
                      (({q0_1[131],q0_0[131]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[131],q0_0[131]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ida095585ad26e215f1c1bf989912da89  <=
                      (Ieeba01b18a244ab8c0ac263c138fabcc) +
                      (({q0_1[132],q0_0[132]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[132],q0_0[132]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I19f1ffa05c7c9a0df5e7014044024c7b  <=
                      (Ie4c9797a955778694dd8615219cb51e7) +
                      (({q0_1[133],q0_0[133]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[133],q0_0[133]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I4d68a2fe778fa93faac38b138138291f  <=
                      (I28a5ed4c239e64c76bb6e566b50cfd23) +
                      (({q0_1[134],q0_0[134]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[134],q0_0[134]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I54393ada6f76ac82c31f2668e228e29d  <=
                      (I79a705ee1e414fe4a5fb14e9b3ce9597) +
                      (({q0_1[135],q0_0[135]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[135],q0_0[135]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If5b9ef84f09680f3593250b13a852c1c  <=
                      (I04f90a907f10a7fa1ae3591b48094d5c) +
                      (({q0_1[136],q0_0[136]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[136],q0_0[136]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibb759bc4179e5b7aa759d850c7cfa467  <=
                      (I31d25b1b49e65216e90b39aa27acd6be) +
                      (({q0_1[137],q0_0[137]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[137],q0_0[137]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I05e8b5f8b83f07b609b5ebf272bb2229  <=
                      (I1f6540c5f037d861dee2c0091cba01ec) +
                      (({q0_1[138],q0_0[138]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[138],q0_0[138]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If6ac15373ec1146d38e7aeb71c3ece64  <=
                      (I9632bb500b7faaaaeb649d74c21cbe8c) +
                      (({q0_1[139],q0_0[139]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[139],q0_0[139]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2ab3675e1eede757af80716ba980a4e6  <=
                      (Idd0217a35c3adc8abc7bb581a5df7a2d) +
                      (({q0_1[140],q0_0[140]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[140],q0_0[140]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I388c271687ab31b57421ad57192273ed  <=
                      (Ic05b46168884322644db4e331d37d759) +
                      (({q0_1[141],q0_0[141]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[141],q0_0[141]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6121679cec8caa51dc5ff0d1a61f9821  <=
                      (I53c88dc237bb2cd02d50fd7f0a168a48) +
                      (({q0_1[142],q0_0[142]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[142],q0_0[142]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia0649b990bf5716cfab230127cd5d47f  <=
                      (I7450d4ab3ef0227e93a02bfd620d047b) +
                      (({q0_1[143],q0_0[143]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[143],q0_0[143]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I867a0626ca22108b16267d95c0aadf4f  <=
                      (I2b16e5b4e279bb29c3c675b72083e5fe) +
                      (({q0_1[144],q0_0[144]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[144],q0_0[144]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I1af54bcb73d7c6b93e55450871207976  <=
                      (I70c92e8ada46476d15ef4b3c620d2601) +
                      (({q0_1[145],q0_0[145]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[145],q0_0[145]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I91883553543d0425e9c6dd726dce3d27  <=
                      (Ib193b07804d6d5f111b06bda487bfa5f) +
                      (({q0_1[146],q0_0[146]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[146],q0_0[146]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie95405659701278e3f87bf1f823a037b  <=
                      (I885433b0ab16c6d87abe45af13c9e529) +
                      (({q0_1[147],q0_0[147]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[147],q0_0[147]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia42392e2104b50c0908aad82738a5ee7  <=
                      (I198c055930cb89d0390c336eda8fed4f) +
                      (({q0_1[148],q0_0[148]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[148],q0_0[148]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I68ad63230a51b9b9e3daffb307ea970d  <=
                      (I688a2c72e69b217d2673e8da75146a83) +
                      (({q0_1[149],q0_0[149]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[149],q0_0[149]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7a052d63944ccf42e598efe3a95b88f8  <=
                      (I3b6fde4ed14cd68af1468ae1d4cc1a22) +
                      (({q0_1[150],q0_0[150]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[150],q0_0[150]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2b3c6d69f79c8d51e4d1614c62c44fcc  <=
                      (I5d3df1e7563630311f56143ee6d97a8e) +
                      (({q0_1[151],q0_0[151]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[151],q0_0[151]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ifcef0e92f50e3920bf1208af5d64c632  <=
                      (I90a7ea789d3bf7f9126c786474a56da0) +
                      (({q0_1[152],q0_0[152]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[152],q0_0[152]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I111340a19625901a3c1b95fd0bd1570e  <=
                      (I5029424c9d9fe923eeb858b1e62cd758) +
                      (({q0_1[153],q0_0[153]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[153],q0_0[153]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I11aec4fa85c30f6fe1fd9fa72542ef6c  <=
                      (I1e805c70d50c2765b4a03ad2982dc421) +
                      (({q0_1[154],q0_0[154]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[154],q0_0[154]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I80cc333c181c16a96b7bd6501c27c2b3  <=
                      (Iba58175a7fd5c5da650222193caff0b3) +
                      (({q0_1[155],q0_0[155]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[155],q0_0[155]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Idc6354325a6280ae9890da33c06c33ec  <=
                      (I7401a0501ba69c5559fbf00c77e58dc5) +
                      (({q0_1[156],q0_0[156]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[156],q0_0[156]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ibb04cf82acc4ac16599ad3ddb0c2ada2  <=
                      (Idd9f7ea657ea9cdcb45a7e4b573b9d50) +
                      (({q0_1[157],q0_0[157]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[157],q0_0[157]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3ed096dfd8a14f4acb4d53a70cf8aceb  <=
                      (I53f275395dd6be17961a5edc3e8da7f2) +
                      (({q0_1[158],q0_0[158]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[158],q0_0[158]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0fa07f95e96326cb0599c0c3f76e2b48  <=
                      (Icab010d78cd66b02e089c74f04bf4e75) +
                      (({q0_1[159],q0_0[159]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[159],q0_0[159]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I87d98fbc97d9a78c2e7d6a6280e7a49a  <=
                      (I376a48b7e0195a5aacc76a0ad8bd14b2) +
                      (({q0_1[160],q0_0[160]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[160],q0_0[160]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib7ddc4dca877f7cf5697a02c3d1915ba  <=
                      (I241622b0367dde514f96ece55c8c3964) +
                      (({q0_1[161],q0_0[161]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[161],q0_0[161]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I3612ef280891f6017fad205d0484bde7  <=
                      (If94a1abfb972f63629d07e64dc23863c) +
                      (({q0_1[162],q0_0[162]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[162],q0_0[162]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I561547649aeb5b4c3f10d9506db1f3cf  <=
                      (I07b9b1f4fa01b16cc69356057d3b6154) +
                      (({q0_1[163],q0_0[163]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[163],q0_0[163]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I84cc76c0079b86da7b994844c3ccb875  <=
                      (I2288a6ad3b748b716249f4adc42d52c4) +
                      (({q0_1[164],q0_0[164]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[164],q0_0[164]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iec013c508d0c6401d7eb856e7eb60446  <=
                      (I022df337bcc05ac5648b8ae2e42f3a76) +
                      (({q0_1[165],q0_0[165]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[165],q0_0[165]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ifd8979aac6b6b24aa560b46b18240e92  <=
                      (I60d9a7f95fb8623753002ecaf9a4efcc) +
                      (({q0_1[166],q0_0[166]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[166],q0_0[166]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If12394e78dc913b01890b56650856a44  <=
                      (I23a74ea5e7174d95e6d16a5e85ac236b) +
                      (({q0_1[167],q0_0[167]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[167],q0_0[167]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I94d18aa10695f3f22b23246884b72822  <=
                      (Ie697d28d757df82b3901564bda43251c) +
                      (({q0_1[168],q0_0[168]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[168],q0_0[168]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic90b38835dd7e760dd54067b196f8470  <=
                      (I8572aedc94f7243ce5eacb332c81eae2) +
                      (({q0_1[169],q0_0[169]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[169],q0_0[169]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               If3691ea51f6efe9b165a31964854d2fe  <=
                      (I6734123aaf6320da75638b212812732f) +
                      (({q0_1[170],q0_0[170]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[170],q0_0[170]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic2ce582555add38a14f5006d3c87eb15  <=
                      (I7f6dc6f0f403c58f9aaaa70c2383a666) +
                      (({q0_1[171],q0_0[171]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[171],q0_0[171]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I58cc950ee2cbe56b7c5a619be3792511  <=
                      (I66391978843c39b6acbdb4847a01050a) +
                      (({q0_1[172],q0_0[172]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[172],q0_0[172]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I0d8e329ec5873db96df1ec309445a096  <=
                      (I4f756e4125c8af5c412944b273e01cb0) +
                      (({q0_1[173],q0_0[173]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[173],q0_0[173]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I106325488e2ecfdba1cf9e5201e6bc8c  <=
                      (Id2c9f7ac95de07148c54803f69347f56) +
                      (({q0_1[174],q0_0[174]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[174],q0_0[174]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iff73a0085541a511d3912b64686a82c5  <=
                      (I5061e13a179d27e1ba5f89ce8ee0fd4a) +
                      (({q0_1[175],q0_0[175]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[175],q0_0[175]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Icdab59de68f2870504598c9ea18f1d2c  <=
                      (I0f7c32fc1548fb49b8041f55c157498a) +
                      (({q0_1[176],q0_0[176]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[176],q0_0[176]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I75604d727e82c977741f90113719183a  <=
                      (I89ffab735ee30423c82e079ed98216c5) +
                      (({q0_1[177],q0_0[177]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[177],q0_0[177]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6f50c4d0d2639857b2dcca300c2d7b04  <=
                      (I9494921d8487ee0b314f75cf0380fd2f) +
                      (({q0_1[178],q0_0[178]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[178],q0_0[178]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5cd013a2be2e761c10c6a957632517de  <=
                      (If2b3e7d1541cbd8ffc2b4cfc3ad13a57) +
                      (({q0_1[179],q0_0[179]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[179],q0_0[179]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iafeedddd02428bd2610c576e68d4ae25  <=
                      (Idf3d79da44f2d686f5bd43c3c1427430) +
                      (({q0_1[180],q0_0[180]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[180],q0_0[180]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I912d6325e34180e0f668f0f024e63581  <=
                      (If8125ad3c9e7f0a2b84106064d320996) +
                      (({q0_1[181],q0_0[181]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[181],q0_0[181]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id1e05294dfd02df499ad0c08bb5c191b  <=
                      (Ic9018b88fa91fb638bbab0613795ae13) +
                      (({q0_1[182],q0_0[182]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[182],q0_0[182]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Id3bb9b100ee4302473b49ac14615e9b0  <=
                      (Iad4ea0196eb32f9a152c9e6fe5059e46) +
                      (({q0_1[183],q0_0[183]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[183],q0_0[183]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ief32db1cfc443119b6202b0cc7bf70a2  <=
                      (Ia8ff29ed728e7f2ae4213f00328b495d) +
                      (({q0_1[184],q0_0[184]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[184],q0_0[184]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Iad7dbe9909b5eed3261adf92d3813acc  <=
                      (I70717726200ec02929f679ef05496455) +
                      (({q0_1[185],q0_0[185]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[185],q0_0[185]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ie7daf0789c35caaadbba06cafabd2b70  <=
                      (Iaf1e4c7dae6ad89567836877c08f57d2) +
                      (({q0_1[186],q0_0[186]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[186],q0_0[186]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2bd1f9b75d9ab94af9ddceb7528935e8  <=
                      (Icd09aa81e9b43528af73e23b2f0f80cb) +
                      (({q0_1[187],q0_0[187]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[187],q0_0[187]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic3d9f5c6677758810e4865779ec303e3  <=
                      (I6ebb2b94f0f80425f8401ae823d92a1d) +
                      (({q0_1[188],q0_0[188]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[188],q0_0[188]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I00af04882a25e2832d913a67d4d86d7b  <=
                      (I4a2c3204a6a9936d4a215b46c0ffd045) +
                      (({q0_1[189],q0_0[189]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[189],q0_0[189]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ic9db631df0a1a9108c10c3e0eca7bf15  <=
                      (Ib02c0694762c4815448b2c8d3df767c2) +
                      (({q0_1[190],q0_0[190]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[190],q0_0[190]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I749f9ed1fb2dddd40ebc28f638e02935  <=
                      (I98cee6efbbe565d3a4de16703189782f) +
                      (({q0_1[191],q0_0[191]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[191],q0_0[191]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ia45b2a24df24bd5e3c95885c8928686c  <=
                      (Ibf981c01a9d44cbea3c6d8ead92bc2ab) +
                      (({q0_1[192],q0_0[192]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[192],q0_0[192]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7427464fde340780aba7f9847b4ad564  <=
                      (I864c33e8ea204d20a9baef4584f22d4e) +
                      (({q0_1[193],q0_0[193]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[193],q0_0[193]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I33fd1ae225e2b881b2b41e0358675e22  <=
                      (I6ad3228e0e2e1f19648d73e83ba5a229) +
                      (({q0_1[194],q0_0[194]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[194],q0_0[194]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2e21a35d1cf560936fd19b944a208b6b  <=
                      (Ie099210a99a4899c53baf39559592690) +
                      (({q0_1[195],q0_0[195]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[195],q0_0[195]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I249522a3d42cc75d7a6b9ede1222ee76  <=
                      (Ieeec71d9df4613555fade2ced7b3baf1) +
                      (({q0_1[196],q0_0[196]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[196],q0_0[196]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I68b4c43d9f40ae4bfd70d2983594392c  <=
                      (I4931884e3544af182bcda9061091a42d) +
                      (({q0_1[197],q0_0[197]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[197],q0_0[197]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I63145e0fec15c7e7c0de105f348bfd31  <=
                      (Ib3fb10da528d450251764a9b9ede0dba) +
                      (({q0_1[198],q0_0[198]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[198],q0_0[198]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I8af625de86c04016c3424d116fddab5b  <=
                      (Icdc9e676957b2223d60c413331fa982f) +
                      (({q0_1[199],q0_0[199]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[199],q0_0[199]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I54c9c10527f83b4ee4e1e22f1e4044ed  <=
                      (I381f6051282c062ccf53866830344cd4) +
                      (({q0_1[200],q0_0[200]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[200],q0_0[200]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I972559e47c7f83bd9000ca1cfc14d8e0  <=
                      (Icfc21935c007fbbceb2a67ebe1a68a0b) +
                      (({q0_1[201],q0_0[201]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[201],q0_0[201]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Ib97a7f941eb7ce2a867503a04ff86a67  <=
                      (I120d597a80158374726e064fb0f099fb) +
                      (({q0_1[202],q0_0[202]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[202],q0_0[202]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I5979b55f607c71017537f2b48b40cbea  <=
                      (I2520aa556aadf851f58f0b1820498730) +
                      (({q0_1[203],q0_0[203]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[203],q0_0[203]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I6a56760b621f238843b091279c69897f  <=
                      (I6203f49a08107f7185ebadeecf2c16b0) +
                      (({q0_1[204],q0_0[204]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[204],q0_0[204]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               Icec45bf76c241d37c9a50a5cd092da9d  <=
                      (Ia706fb593b63cebbee0321c154cb859b) +
                      (({q0_1[205],q0_0[205]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[205],q0_0[205]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I2f6d3f61f2890e584d3063a09587e99b  <=
                      (Ia4b5f2b07556629673fc6576bc49a5dc) +
                      (({q0_1[206],q0_0[206]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[206],q0_0[206]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"
               I7c396ea2e959d84fd9a6964617cb29c6  <=
                      (Ic532c6b85b156f821e0742f47239a65c) +
                      (({q0_1[207],q0_0[207]} ==2'b11) ? ~percent_probability_int + 1 :
                      (({q0_1[207],q0_0[207]} ==2'b01) ? percent_probability_int :
                      32'h0));
                    // 2'b11 === -1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b1
                    // 2'b01 ===  1 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for 1'b0
                    // 2'b00 ===  I4a548addbfb239bbd12f5afe11a4b6dc I8bf8854bebe108183caeb845c7676ae4 -1:1 and 1:0 Icfd8f331d281b0da79e7c6ed6988243c I8b7af514f25f1f9456dcd10d2337f753 Ia2a551a6458a8de22446cc76d639a9e9 bit I2063c1608d6e0baf80249c42e2be5804 for "Iad921d60486366258809553a3db49a4a"

                 if ({q0_1[0],q0_0[0]} != 1 ) begin
                 end
                 if ({q0_1[1],q0_0[1]} != 1 ) begin
                 end
                 if ({q0_1[2],q0_0[2]} != 0 ) begin
                 end
                 if ({q0_1[3],q0_0[3]} != 1 ) begin
                 end
                 if ({q0_1[4],q0_0[4]} != 0 ) begin
                 end
                 if ({q0_1[5],q0_0[5]} != 0 ) begin
                 end
                 if ({q0_1[6],q0_0[6]} != 0 ) begin
                 end
                 if ({q0_1[7],q0_0[7]} != 0 ) begin
                 end
                 if ({q0_1[8],q0_0[8]} != 0 ) begin
                 end
                 if ({q0_1[9],q0_0[9]} != 1 ) begin
                 end
                 if ({q0_1[10],q0_0[10]} != 1 ) begin
                 end
                 if ({q0_1[11],q0_0[11]} != 1 ) begin
                 end
                 if ({q0_1[12],q0_0[12]} != 1 ) begin
                 end
                 if ({q0_1[13],q0_0[13]} != 1 ) begin
                 end
                 if ({q0_1[14],q0_0[14]} != 0 ) begin
                 end
                 if ({q0_1[15],q0_0[15]} != 1 ) begin
                 end
                 if ({q0_1[16],q0_0[16]} != 0 ) begin
                 end
                 if ({q0_1[17],q0_0[17]} != 0 ) begin
                 end
                 if ({q0_1[18],q0_0[18]} != 1 ) begin
                 end
                 if ({q0_1[19],q0_0[19]} != 0 ) begin
                 end
                 if ({q0_1[20],q0_0[20]} != 1 ) begin
                 end
                 if ({q0_1[21],q0_0[21]} != 1 ) begin
                 end
                 if ({q0_1[22],q0_0[22]} != 0 ) begin
                 end
                 if ({q0_1[23],q0_0[23]} != 0 ) begin
                 end
                 if ({q0_1[24],q0_0[24]} != 0 ) begin
                 end
                 if ({q0_1[25],q0_0[25]} != 1 ) begin
                 end
                 if ({q0_1[26],q0_0[26]} != 1 ) begin
                 end
                 if ({q0_1[27],q0_0[27]} != 0 ) begin
                 end
                 if ({q0_1[28],q0_0[28]} != 0 ) begin
                 end
                 if ({q0_1[29],q0_0[29]} != 1 ) begin
                 end
                 if ({q0_1[30],q0_0[30]} != 1 ) begin
                 end
                 if ({q0_1[31],q0_0[31]} != 1 ) begin
                 end
                 if ({q0_1[32],q0_0[32]} != 0 ) begin
                 end
                 if ({q0_1[33],q0_0[33]} != 0 ) begin
                 end
                 if ({q0_1[34],q0_0[34]} != 1 ) begin
                 end
                 if ({q0_1[35],q0_0[35]} != 0 ) begin
                 end
                 if ({q0_1[36],q0_0[36]} != 0 ) begin
                 end
                 if ({q0_1[37],q0_0[37]} != 0 ) begin
                 end
                 if ({q0_1[38],q0_0[38]} != 0 ) begin
                 end
                 if ({q0_1[39],q0_0[39]} != 0 ) begin
                 end
                 if ({q0_1[40],q0_0[40]} != 1 ) begin
                 end
                 if ({q0_1[41],q0_0[41]} != 0 ) begin
                 end
                 if ({q0_1[42],q0_0[42]} != 0 ) begin
                 end
                 if ({q0_1[43],q0_0[43]} != 1 ) begin
                 end
                 if ({q0_1[44],q0_0[44]} != 1 ) begin
                 end
                 if ({q0_1[45],q0_0[45]} != 1 ) begin
                 end
                 if ({q0_1[46],q0_0[46]} != 1 ) begin
                 end
                 if ({q0_1[47],q0_0[47]} != 0 ) begin
                 end
                 if ({q0_1[48],q0_0[48]} != 0 ) begin
                 end
                 if ({q0_1[49],q0_0[49]} != 1 ) begin
                 end
                 if ({q0_1[50],q0_0[50]} != 1 ) begin
                 end
                 if ({q0_1[51],q0_0[51]} != 0 ) begin
                 end
                 if ({q0_1[52],q0_0[52]} != 1 ) begin
                 end
                 if ({q0_1[53],q0_0[53]} != 1 ) begin
                 end
                 if ({q0_1[54],q0_0[54]} != 0 ) begin
                 end
                 if ({q0_1[55],q0_0[55]} != 1 ) begin
                 end
                 if ({q0_1[56],q0_0[56]} != 1 ) begin
                 end
                 if ({q0_1[57],q0_0[57]} != 0 ) begin
                 end
                 if ({q0_1[58],q0_0[58]} != 0 ) begin
                 end
                 if ({q0_1[59],q0_0[59]} != 1 ) begin
                 end
                 if ({q0_1[60],q0_0[60]} != 0 ) begin
                 end
                 if ({q0_1[61],q0_0[61]} != 0 ) begin
                 end
                 if ({q0_1[62],q0_0[62]} != 0 ) begin
                 end
                 if ({q0_1[63],q0_0[63]} != 1 ) begin
                 end
                 if ({q0_1[64],q0_0[64]} != 0 ) begin
                 end
                 if ({q0_1[65],q0_0[65]} != 1 ) begin
                 end
                 if ({q0_1[66],q0_0[66]} != 1 ) begin
                 end
                 if ({q0_1[67],q0_0[67]} != 1 ) begin
                 end
                 if ({q0_1[68],q0_0[68]} != 1 ) begin
                 end
                 if ({q0_1[69],q0_0[69]} != 1 ) begin
                 end
                 if ({q0_1[70],q0_0[70]} != 1 ) begin
                 end
                 if ({q0_1[71],q0_0[71]} != 1 ) begin
                 end
                 if ({q0_1[72],q0_0[72]} != 0 ) begin
                 end
                 if ({q0_1[73],q0_0[73]} != 0 ) begin
                 end
                 if ({q0_1[74],q0_0[74]} != 1 ) begin
                 end
                 if ({q0_1[75],q0_0[75]} != 0 ) begin
                 end
                 if ({q0_1[76],q0_0[76]} != 0 ) begin
                 end
                 if ({q0_1[77],q0_0[77]} != 0 ) begin
                 end
                 if ({q0_1[78],q0_0[78]} != 0 ) begin
                 end
                 if ({q0_1[79],q0_0[79]} != 0 ) begin
                 end
                 if ({q0_1[80],q0_0[80]} != 0 ) begin
                 end
                 if ({q0_1[81],q0_0[81]} != 1 ) begin
                 end
                 if ({q0_1[82],q0_0[82]} != 1 ) begin
                 end
                 if ({q0_1[83],q0_0[83]} != 0 ) begin
                 end
                 if ({q0_1[84],q0_0[84]} != 0 ) begin
                 end
                 if ({q0_1[85],q0_0[85]} != 0 ) begin
                 end
                 if ({q0_1[86],q0_0[86]} != 0 ) begin
                 end
                 if ({q0_1[87],q0_0[87]} != 0 ) begin
                 end
                 if ({q0_1[88],q0_0[88]} != 0 ) begin
                 end
                 if ({q0_1[89],q0_0[89]} != 1 ) begin
                 end
                 if ({q0_1[90],q0_0[90]} != 0 ) begin
                 end
                 if ({q0_1[91],q0_0[91]} != 1 ) begin
                 end
                 if ({q0_1[92],q0_0[92]} != 0 ) begin
                 end
                 if ({q0_1[93],q0_0[93]} != 0 ) begin
                 end
                 if ({q0_1[94],q0_0[94]} != 0 ) begin
                 end
                 if ({q0_1[95],q0_0[95]} != 0 ) begin
                 end
                 if ({q0_1[96],q0_0[96]} != 0 ) begin
                 end
                 if ({q0_1[97],q0_0[97]} != 0 ) begin
                 end
                 if ({q0_1[98],q0_0[98]} != 0 ) begin
                 end
                 if ({q0_1[99],q0_0[99]} != 0 ) begin
                 end
                 if ({q0_1[100],q0_0[100]} != 1 ) begin
                 end
                 if ({q0_1[101],q0_0[101]} != 1 ) begin
                 end
                 if ({q0_1[102],q0_0[102]} != 1 ) begin
                 end
                 if ({q0_1[103],q0_0[103]} != 1 ) begin
                 end
                 if ({q0_1[104],q0_0[104]} != 0 ) begin
                 end
                 if ({q0_1[105],q0_0[105]} != 1 ) begin
                 end
                 if ({q0_1[106],q0_0[106]} != 1 ) begin
                 end
                 if ({q0_1[107],q0_0[107]} != 1 ) begin
                 end
                 if ({q0_1[108],q0_0[108]} != 0 ) begin
                 end
                 if ({q0_1[109],q0_0[109]} != 0 ) begin
                 end
                 if ({q0_1[110],q0_0[110]} != 0 ) begin
                 end
                 if ({q0_1[111],q0_0[111]} != 1 ) begin
                 end
                 if ({q0_1[112],q0_0[112]} != 1 ) begin
                 end
                 if ({q0_1[113],q0_0[113]} != 0 ) begin
                 end
                 if ({q0_1[114],q0_0[114]} != 0 ) begin
                 end
                 if ({q0_1[115],q0_0[115]} != 1 ) begin
                 end
                 if ({q0_1[116],q0_0[116]} != 1 ) begin
                 end
                 if ({q0_1[117],q0_0[117]} != 1 ) begin
                 end
                 if ({q0_1[118],q0_0[118]} != 1 ) begin
                 end
                 if ({q0_1[119],q0_0[119]} != 0 ) begin
                 end
                 if ({q0_1[120],q0_0[120]} != 1 ) begin
                 end
                 if ({q0_1[121],q0_0[121]} != 0 ) begin
                 end
                 if ({q0_1[122],q0_0[122]} != 0 ) begin
                 end
                 if ({q0_1[123],q0_0[123]} != 1 ) begin
                 end
                 if ({q0_1[124],q0_0[124]} != 0 ) begin
                 end
                 if ({q0_1[125],q0_0[125]} != 0 ) begin
                 end
                 if ({q0_1[126],q0_0[126]} != 1 ) begin
                 end
                 if ({q0_1[127],q0_0[127]} != 1 ) begin
                 end
                 if ({q0_1[128],q0_0[128]} != 1 ) begin
                 end
                 if ({q0_1[129],q0_0[129]} != 0 ) begin
                 end
                 if ({q0_1[130],q0_0[130]} != 1 ) begin
                 end
                 if ({q0_1[131],q0_0[131]} != 0 ) begin
                 end
                 if ({q0_1[132],q0_0[132]} != 0 ) begin
                 end
                 if ({q0_1[133],q0_0[133]} != 0 ) begin
                 end
                 if ({q0_1[134],q0_0[134]} != 1 ) begin
                 end
                 if ({q0_1[135],q0_0[135]} != 1 ) begin
                 end
                 if ({q0_1[136],q0_0[136]} != 1 ) begin
                 end
                 if ({q0_1[137],q0_0[137]} != 0 ) begin
                 end
                 if ({q0_1[138],q0_0[138]} != 1 ) begin
                 end
                 if ({q0_1[139],q0_0[139]} != 1 ) begin
                 end
                 if ({q0_1[140],q0_0[140]} != 1 ) begin
                 end
                 if ({q0_1[141],q0_0[141]} != 0 ) begin
                 end
                 if ({q0_1[142],q0_0[142]} != 0 ) begin
                 end
                 if ({q0_1[143],q0_0[143]} != 1 ) begin
                 end
                 if ({q0_1[144],q0_0[144]} != 0 ) begin
                 end
                 if ({q0_1[145],q0_0[145]} != 1 ) begin
                 end
                 if ({q0_1[146],q0_0[146]} != 0 ) begin
                 end
                 if ({q0_1[147],q0_0[147]} != 1 ) begin
                 end
                 if ({q0_1[148],q0_0[148]} != 1 ) begin
                 end
                 if ({q0_1[149],q0_0[149]} != 1 ) begin
                 end
                 if ({q0_1[150],q0_0[150]} != 1 ) begin
                 end
                 if ({q0_1[151],q0_0[151]} != 0 ) begin
                 end
                 if ({q0_1[152],q0_0[152]} != 1 ) begin
                 end
                 if ({q0_1[153],q0_0[153]} != 0 ) begin
                 end
                 if ({q0_1[154],q0_0[154]} != 0 ) begin
                 end
                 if ({q0_1[155],q0_0[155]} != 0 ) begin
                 end
                 if ({q0_1[156],q0_0[156]} != 0 ) begin
                 end
                 if ({q0_1[157],q0_0[157]} != 1 ) begin
                 end
                 if ({q0_1[158],q0_0[158]} != 0 ) begin
                 end
                 if ({q0_1[159],q0_0[159]} != 1 ) begin
                 end
                 if ({q0_1[160],q0_0[160]} != 1 ) begin
                 end
                 if ({q0_1[161],q0_0[161]} != 0 ) begin
                 end
                 if ({q0_1[162],q0_0[162]} != 0 ) begin
                 end
                 if ({q0_1[163],q0_0[163]} != 1 ) begin
                 end
                 if ({q0_1[164],q0_0[164]} != 0 ) begin
                 end
                 if ({q0_1[165],q0_0[165]} != 0 ) begin
                 end
                 if ({q0_1[166],q0_0[166]} != 1 ) begin
                 end
                 if ({q0_1[167],q0_0[167]} != 1 ) begin
                 end
                 if ({q0_1[168],q0_0[168]} != 0 ) begin
                 end
                 if ({q0_1[169],q0_0[169]} != 0 ) begin
                 end
                 if ({q0_1[170],q0_0[170]} != 1 ) begin
                 end
                 if ({q0_1[171],q0_0[171]} != 0 ) begin
                 end
                 if ({q0_1[172],q0_0[172]} != 1 ) begin
                 end
                 if ({q0_1[173],q0_0[173]} != 1 ) begin
                 end
                 if ({q0_1[174],q0_0[174]} != 0 ) begin
                 end
                 if ({q0_1[175],q0_0[175]} != 0 ) begin
                 end
                 if ({q0_1[176],q0_0[176]} != 1 ) begin
                 end
                 if ({q0_1[177],q0_0[177]} != 0 ) begin
                 end
                 if ({q0_1[178],q0_0[178]} != 1 ) begin
                 end
                 if ({q0_1[179],q0_0[179]} != 1 ) begin
                 end
                 if ({q0_1[180],q0_0[180]} != 1 ) begin
                 end
                 if ({q0_1[181],q0_0[181]} != 0 ) begin
                 end
                 if ({q0_1[182],q0_0[182]} != 1 ) begin
                 end
                 if ({q0_1[183],q0_0[183]} != 1 ) begin
                 end
                 if ({q0_1[184],q0_0[184]} != 1 ) begin
                 end
                 if ({q0_1[185],q0_0[185]} != 1 ) begin
                 end
                 if ({q0_1[186],q0_0[186]} != 0 ) begin
                 end
                 if ({q0_1[187],q0_0[187]} != 1 ) begin
                 end
                 if ({q0_1[188],q0_0[188]} != 0 ) begin
                 end
                 if ({q0_1[189],q0_0[189]} != 0 ) begin
                 end
                 if ({q0_1[190],q0_0[190]} != 0 ) begin
                 end
                 if ({q0_1[191],q0_0[191]} != 0 ) begin
                 end
                 if ({q0_1[192],q0_0[192]} != 1 ) begin
                 end
                 if ({q0_1[193],q0_0[193]} != 0 ) begin
                 end
                 if ({q0_1[194],q0_0[194]} != 0 ) begin
                 end
                 if ({q0_1[195],q0_0[195]} != 0 ) begin
                 end
                 if ({q0_1[196],q0_0[196]} != 0 ) begin
                 end
                 if ({q0_1[197],q0_0[197]} != 0 ) begin
                 end
                 if ({q0_1[198],q0_0[198]} != 0 ) begin
                 end
                 if ({q0_1[199],q0_0[199]} != 0 ) begin
                 end
                 if ({q0_1[200],q0_0[200]} != 0 ) begin
                 end
                 if ({q0_1[201],q0_0[201]} != 0 ) begin
                 end
                 if ({q0_1[202],q0_0[202]} != 1 ) begin
                 end
                 if ({q0_1[203],q0_0[203]} != 0 ) begin
                 end
                 if ({q0_1[204],q0_0[204]} != 0 ) begin
                 end
                 if ({q0_1[205],q0_0[205]} != 0 ) begin
                 end
                 if ({q0_1[206],q0_0[206]} != 1 ) begin
                 end
                 if ({q0_1[207],q0_0[207]} != 0 ) begin
                 end


           end

           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic93835a022c46b7aa00a465c407d7da2     <=
                                             Ic05b492587d8d5083e8570900995293a[SGN_MAX_SUM_WDTH] ?
                                             ~Ic05b492587d8d5083e8570900995293a + 1 :
                                             Ic05b492587d8d5083e8570900995293a
                                             ;

            I92cb615e2c439914e72ce001256518e4  <=  Ic05b492587d8d5083e8570900995293a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2e30088bf29cedd7debc15b1e6ec4ada     <=
                                             Ibee9ba58404f1adb9e4e8e6f822a38c1[SGN_MAX_SUM_WDTH] ?
                                             ~Ibee9ba58404f1adb9e4e8e6f822a38c1 + 1 :
                                             Ibee9ba58404f1adb9e4e8e6f822a38c1
                                             ;

            Iad799775eb657f8973e6dfcf70a9875c  <=  Ibee9ba58404f1adb9e4e8e6f822a38c1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I38f512bfb84094d1e92a10a345d5505f     <=
                                             Ifab38317b76e52f9d9d64bed976e2cc5[SGN_MAX_SUM_WDTH] ?
                                             ~Ifab38317b76e52f9d9d64bed976e2cc5 + 1 :
                                             Ifab38317b76e52f9d9d64bed976e2cc5
                                             ;

            Ifb064c69c7110c014593149ae69c75fb  <=  Ifab38317b76e52f9d9d64bed976e2cc5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1e878f00f056f637625cb013a93325a8     <=
                                             I86195d9a1da88ffc163298c54401039e[SGN_MAX_SUM_WDTH] ?
                                             ~I86195d9a1da88ffc163298c54401039e + 1 :
                                             I86195d9a1da88ffc163298c54401039e
                                             ;

            I7f7b30f2acbb8e31f50b58096b738254  <=  I86195d9a1da88ffc163298c54401039e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I25db27464b31fee41ccd7a3cfe4d403e     <=
                                             I27c02895bfd59c762d5c7a725aa5cefd[SGN_MAX_SUM_WDTH] ?
                                             ~I27c02895bfd59c762d5c7a725aa5cefd + 1 :
                                             I27c02895bfd59c762d5c7a725aa5cefd
                                             ;

            Iefe4099ff7e457f6b9fefc83e176c1a0  <=  I27c02895bfd59c762d5c7a725aa5cefd[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I19417a224c5cdf1211e9790aa29c4c5c     <=
                                             I60de515e03218ac363566ce7b92f5034[SGN_MAX_SUM_WDTH] ?
                                             ~I60de515e03218ac363566ce7b92f5034 + 1 :
                                             I60de515e03218ac363566ce7b92f5034
                                             ;

            Icddb43f9b760a4597a0bb637fb405616  <=  I60de515e03218ac363566ce7b92f5034[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I16dcafa854ea9c67d8a080feb2ba9166     <=
                                             I9b75e7451fbf27c3645bebbdba234996[SGN_MAX_SUM_WDTH] ?
                                             ~I9b75e7451fbf27c3645bebbdba234996 + 1 :
                                             I9b75e7451fbf27c3645bebbdba234996
                                             ;

            Ic76e72b434b47c10ebac3fac4ea50bde  <=  I9b75e7451fbf27c3645bebbdba234996[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7f63338eee2663fbe61fffd248433310     <=
                                             I056c79002bbba10ddee2448e36dc7478[SGN_MAX_SUM_WDTH] ?
                                             ~I056c79002bbba10ddee2448e36dc7478 + 1 :
                                             I056c79002bbba10ddee2448e36dc7478
                                             ;

            I9eb87e62d23bc87d7cd82c0f329f247f  <=  I056c79002bbba10ddee2448e36dc7478[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icb1e3c56c8729c32d43c69710e345db2     <=
                                             Ia5db5f66b7fb04e2344abff9b4f75404[SGN_MAX_SUM_WDTH] ?
                                             ~Ia5db5f66b7fb04e2344abff9b4f75404 + 1 :
                                             Ia5db5f66b7fb04e2344abff9b4f75404
                                             ;

            I2eac5b39c6f485c9ae0bd341f894633d  <=  Ia5db5f66b7fb04e2344abff9b4f75404[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ece8e3c1e89613879336936f77d732f     <=
                                             I250898de23a8793f0c21eb333d61af53[SGN_MAX_SUM_WDTH] ?
                                             ~I250898de23a8793f0c21eb333d61af53 + 1 :
                                             I250898de23a8793f0c21eb333d61af53
                                             ;

            I76992221b1edff5684c482df7ac4693d  <=  I250898de23a8793f0c21eb333d61af53[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I72a646ae7e32a16af0f5930a6e95b36a     <=
                                             I1320273c298c7953b3227b58439b54c4[SGN_MAX_SUM_WDTH] ?
                                             ~I1320273c298c7953b3227b58439b54c4 + 1 :
                                             I1320273c298c7953b3227b58439b54c4
                                             ;

            Iada5bc4a51dc1bf57bb9cca11326bdff  <=  I1320273c298c7953b3227b58439b54c4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7e72d119dd93a6ab05a23fde0a865866     <=
                                             I49a036af196fb318309a43c150540a2c[SGN_MAX_SUM_WDTH] ?
                                             ~I49a036af196fb318309a43c150540a2c + 1 :
                                             I49a036af196fb318309a43c150540a2c
                                             ;

            I364ed3f83c49626bc3b939e53524d9c7  <=  I49a036af196fb318309a43c150540a2c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ied4fdf5805039cd2fcd042fd13755fdc     <=
                                             If115c3e5f121363c2b8a6c14905aebe7[SGN_MAX_SUM_WDTH] ?
                                             ~If115c3e5f121363c2b8a6c14905aebe7 + 1 :
                                             If115c3e5f121363c2b8a6c14905aebe7
                                             ;

            Ic2b000c3b2ca3beff2d427caab04701a  <=  If115c3e5f121363c2b8a6c14905aebe7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id44c2293b765cff450dd1d747c47c1f3     <=
                                             I5fcd95690fb291f9b95996e687de022c[SGN_MAX_SUM_WDTH] ?
                                             ~I5fcd95690fb291f9b95996e687de022c + 1 :
                                             I5fcd95690fb291f9b95996e687de022c
                                             ;

            I8e873fb2321eea82bb590a92411e2e2c  <=  I5fcd95690fb291f9b95996e687de022c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f4ed02f7aeb823b745040f7f3f43ac7     <=
                                             I5f6f8a4c5c5ab4cf1f9c496795c41ce8[SGN_MAX_SUM_WDTH] ?
                                             ~I5f6f8a4c5c5ab4cf1f9c496795c41ce8 + 1 :
                                             I5f6f8a4c5c5ab4cf1f9c496795c41ce8
                                             ;

            If4cb744ee52b6ae793431cd038069b57  <=  I5f6f8a4c5c5ab4cf1f9c496795c41ce8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6488b9b8f405d7d81a4874fab2678102     <=
                                             I775180b845280ec240e4adf20605b8fe[SGN_MAX_SUM_WDTH] ?
                                             ~I775180b845280ec240e4adf20605b8fe + 1 :
                                             I775180b845280ec240e4adf20605b8fe
                                             ;

            I7741e239c16828889d488cc87647c154  <=  I775180b845280ec240e4adf20605b8fe[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifff612d16828ec907a348479e19ddf31     <=
                                             I642fe2c7978d7229d660431061a6f781[SGN_MAX_SUM_WDTH] ?
                                             ~I642fe2c7978d7229d660431061a6f781 + 1 :
                                             I642fe2c7978d7229d660431061a6f781
                                             ;

            I7979161aa1e2262ebea862004c387697  <=  I642fe2c7978d7229d660431061a6f781[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I268262076f22bc6b1507bc8f91b98a0a     <=
                                             I3ce66aa6048542c81a89c28e80412e70[SGN_MAX_SUM_WDTH] ?
                                             ~I3ce66aa6048542c81a89c28e80412e70 + 1 :
                                             I3ce66aa6048542c81a89c28e80412e70
                                             ;

            Ic62fc602da3d16fe13d03a49a21269d0  <=  I3ce66aa6048542c81a89c28e80412e70[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If1f732841adb7c0cad1ba37c0f5fd517     <=
                                             I436fc89b03a41f35b8d2ab89464d07c0[SGN_MAX_SUM_WDTH] ?
                                             ~I436fc89b03a41f35b8d2ab89464d07c0 + 1 :
                                             I436fc89b03a41f35b8d2ab89464d07c0
                                             ;

            I94009bb7239be96243902ab0f0abea7e  <=  I436fc89b03a41f35b8d2ab89464d07c0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0df8a24f31c027756d248c3bd1b9bf7b     <=
                                             I67861da88ed0edc52bb876287fc60261[SGN_MAX_SUM_WDTH] ?
                                             ~I67861da88ed0edc52bb876287fc60261 + 1 :
                                             I67861da88ed0edc52bb876287fc60261
                                             ;

            Iae7b72abf4d3c536330a229e3836b441  <=  I67861da88ed0edc52bb876287fc60261[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8ef901e733b12e76412eb36684e2b575     <=
                                             If51bec96c3139419947f0442b0ad7281[SGN_MAX_SUM_WDTH] ?
                                             ~If51bec96c3139419947f0442b0ad7281 + 1 :
                                             If51bec96c3139419947f0442b0ad7281
                                             ;

            Ie5d9cc18b2dd300132470f206452ff17  <=  If51bec96c3139419947f0442b0ad7281[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia48916a02f68b1b8f5fc7fece04677bb     <=
                                             I5e126994711cd1782fcbd2fb3eec3cdc[SGN_MAX_SUM_WDTH] ?
                                             ~I5e126994711cd1782fcbd2fb3eec3cdc + 1 :
                                             I5e126994711cd1782fcbd2fb3eec3cdc
                                             ;

            I7c791c854d0bc28e8dd787545f8fbda0  <=  I5e126994711cd1782fcbd2fb3eec3cdc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia37409944d9fdd3b16e7007e13d82a79     <=
                                             I44d2fe323e921ba0fd66c82a792302e1[SGN_MAX_SUM_WDTH] ?
                                             ~I44d2fe323e921ba0fd66c82a792302e1 + 1 :
                                             I44d2fe323e921ba0fd66c82a792302e1
                                             ;

            I5b177dd5c14ad082516b47f550875682  <=  I44d2fe323e921ba0fd66c82a792302e1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idd65f149afe9d5f63ddaf34b82b11e95     <=
                                             I875b53feb16dc1ac263e9d1c2552dd38[SGN_MAX_SUM_WDTH] ?
                                             ~I875b53feb16dc1ac263e9d1c2552dd38 + 1 :
                                             I875b53feb16dc1ac263e9d1c2552dd38
                                             ;

            I55e4ad2d71a29ad63b4999d64ac0dc4f  <=  I875b53feb16dc1ac263e9d1c2552dd38[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If2886d560854faed32ebd8e33d868973     <=
                                             I651f168318d2ce4746ade3230e052ace[SGN_MAX_SUM_WDTH] ?
                                             ~I651f168318d2ce4746ade3230e052ace + 1 :
                                             I651f168318d2ce4746ade3230e052ace
                                             ;

            I59c5da6338f431a626c86a065a355c35  <=  I651f168318d2ce4746ade3230e052ace[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I77778118bb3ea900c080754ff4c49c26     <=
                                             I00a65dc6a94fa280ec3aac7b04fd4aba[SGN_MAX_SUM_WDTH] ?
                                             ~I00a65dc6a94fa280ec3aac7b04fd4aba + 1 :
                                             I00a65dc6a94fa280ec3aac7b04fd4aba
                                             ;

            Ia098bbeda8b755ece6b88eac83d03e55  <=  I00a65dc6a94fa280ec3aac7b04fd4aba[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7292ed752d8741594d757730950feea4     <=
                                             I38f5eb8d994476d2edb5fd71b7636452[SGN_MAX_SUM_WDTH] ?
                                             ~I38f5eb8d994476d2edb5fd71b7636452 + 1 :
                                             I38f5eb8d994476d2edb5fd71b7636452
                                             ;

            Ie7470dd75b54d14038de19e4d3043ba9  <=  I38f5eb8d994476d2edb5fd71b7636452[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I68cfd7868e061793ee8a41e69e80219b     <=
                                             If0d9102fbff225bd3ef4f4e1aab2811b[SGN_MAX_SUM_WDTH] ?
                                             ~If0d9102fbff225bd3ef4f4e1aab2811b + 1 :
                                             If0d9102fbff225bd3ef4f4e1aab2811b
                                             ;

            Ie95662d4faf6b5a4cd5ecfa41697b983  <=  If0d9102fbff225bd3ef4f4e1aab2811b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I667ead814b303fca64ef047bb8246b19     <=
                                             I09734a3840b1b01a467b075c65608f3e[SGN_MAX_SUM_WDTH] ?
                                             ~I09734a3840b1b01a467b075c65608f3e + 1 :
                                             I09734a3840b1b01a467b075c65608f3e
                                             ;

            Ia1b617e3d141263b51e58c5ef0bd7a89  <=  I09734a3840b1b01a467b075c65608f3e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4f25c7edb12e868cb5532e42b4ba5133     <=
                                             Icec563470fe1bec10dfa8d36561f6ed7[SGN_MAX_SUM_WDTH] ?
                                             ~Icec563470fe1bec10dfa8d36561f6ed7 + 1 :
                                             Icec563470fe1bec10dfa8d36561f6ed7
                                             ;

            If9a5d830e3ade0fd96b98f5949f165f0  <=  Icec563470fe1bec10dfa8d36561f6ed7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5aed2d82717f359bb5ac5a0ab91b7beb     <=
                                             Iaa82bbd78ea7acbc1949f7db44d339eb[SGN_MAX_SUM_WDTH] ?
                                             ~Iaa82bbd78ea7acbc1949f7db44d339eb + 1 :
                                             Iaa82bbd78ea7acbc1949f7db44d339eb
                                             ;

            Id3de87169c440f95d406693ef77cacd6  <=  Iaa82bbd78ea7acbc1949f7db44d339eb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I92835fd54631deaefa7b214e2c4b9bff     <=
                                             I1bf879a8671257cec876577804bd6ffb[SGN_MAX_SUM_WDTH] ?
                                             ~I1bf879a8671257cec876577804bd6ffb + 1 :
                                             I1bf879a8671257cec876577804bd6ffb
                                             ;

            I3751f191f5009322acb7c9be4f8d7129  <=  I1bf879a8671257cec876577804bd6ffb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I67e067da565635fcff166e3a7d0c446b     <=
                                             Ifdb571f08bb8fc78631b0af95d6f5b68[SGN_MAX_SUM_WDTH] ?
                                             ~Ifdb571f08bb8fc78631b0af95d6f5b68 + 1 :
                                             Ifdb571f08bb8fc78631b0af95d6f5b68
                                             ;

            Ic1927bb3335f6a28c0816eba12d3975e  <=  Ifdb571f08bb8fc78631b0af95d6f5b68[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifdb0f307b1b9458c0487a1574ccc094b     <=
                                             I06117d4a9cec69582f336796f82af871[SGN_MAX_SUM_WDTH] ?
                                             ~I06117d4a9cec69582f336796f82af871 + 1 :
                                             I06117d4a9cec69582f336796f82af871
                                             ;

            Ia659126b51468cfef48c97a135a71500  <=  I06117d4a9cec69582f336796f82af871[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5c6b7d143e42fd3b8bcdb7d7ed4da2c2     <=
                                             I23178a40d717727916e4c44fb8ea7de9[SGN_MAX_SUM_WDTH] ?
                                             ~I23178a40d717727916e4c44fb8ea7de9 + 1 :
                                             I23178a40d717727916e4c44fb8ea7de9
                                             ;

            I3c3c22bf63e55a81ae91b1dd1ef615a0  <=  I23178a40d717727916e4c44fb8ea7de9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie679a21d0136a08cc5e6526e9f8d1843     <=
                                             Idd1454bc7f85ca3c184a20fd0864c666[SGN_MAX_SUM_WDTH] ?
                                             ~Idd1454bc7f85ca3c184a20fd0864c666 + 1 :
                                             Idd1454bc7f85ca3c184a20fd0864c666
                                             ;

            Ia62832d325f86160285c4d1a790a32cb  <=  Idd1454bc7f85ca3c184a20fd0864c666[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I611942a72a5e12f6afaea6bde6699ef6     <=
                                             Iee01a4b6a910ede0b61e2465d7d5d696[SGN_MAX_SUM_WDTH] ?
                                             ~Iee01a4b6a910ede0b61e2465d7d5d696 + 1 :
                                             Iee01a4b6a910ede0b61e2465d7d5d696
                                             ;

            I83c7d177eec2dad0a924557cdc91ba77  <=  Iee01a4b6a910ede0b61e2465d7d5d696[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica9883c97f823a4491cbee5b45c43590     <=
                                             I383d6b1028ae1e4e2ea40cfa22043d72[SGN_MAX_SUM_WDTH] ?
                                             ~I383d6b1028ae1e4e2ea40cfa22043d72 + 1 :
                                             I383d6b1028ae1e4e2ea40cfa22043d72
                                             ;

            I7050adb9d06f767549b7f35c4679e391  <=  I383d6b1028ae1e4e2ea40cfa22043d72[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8e6addfc61f5bfb7af74fc2993639565     <=
                                             Ifde4b0c41d42daf9b134ee6c05db336a[SGN_MAX_SUM_WDTH] ?
                                             ~Ifde4b0c41d42daf9b134ee6c05db336a + 1 :
                                             Ifde4b0c41d42daf9b134ee6c05db336a
                                             ;

            I04aacd95d9e44657f616e01c9053f0fb  <=  Ifde4b0c41d42daf9b134ee6c05db336a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9d53619f10e2a426f7297bbf7c81158a     <=
                                             I9f0b1952f54a14726de1d31a2302a95f[SGN_MAX_SUM_WDTH] ?
                                             ~I9f0b1952f54a14726de1d31a2302a95f + 1 :
                                             I9f0b1952f54a14726de1d31a2302a95f
                                             ;

            I2ff317d57f59747c4524ef4278d51092  <=  I9f0b1952f54a14726de1d31a2302a95f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8a055c27778913287ad951183fa0d4d6     <=
                                             I3991c8d4f24af7dfb52a65f70c3ab2d5[SGN_MAX_SUM_WDTH] ?
                                             ~I3991c8d4f24af7dfb52a65f70c3ab2d5 + 1 :
                                             I3991c8d4f24af7dfb52a65f70c3ab2d5
                                             ;

            I8bd2a9d90074500698b302cb8db7f03a  <=  I3991c8d4f24af7dfb52a65f70c3ab2d5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f6ae5c80bb2f50084b5f5ee5ab0ffc3     <=
                                             Ie928ef6ba83900dca8b150428d713448[SGN_MAX_SUM_WDTH] ?
                                             ~Ie928ef6ba83900dca8b150428d713448 + 1 :
                                             Ie928ef6ba83900dca8b150428d713448
                                             ;

            I3b8cdfb1440732ce98cd1676e05a2af1  <=  Ie928ef6ba83900dca8b150428d713448[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3db8b3a342e8e2f13a448246aa001c2f     <=
                                             Ic085f1faeb81e3027f909a7bd890d359[SGN_MAX_SUM_WDTH] ?
                                             ~Ic085f1faeb81e3027f909a7bd890d359 + 1 :
                                             Ic085f1faeb81e3027f909a7bd890d359
                                             ;

            I671de3d408b5b783541663c7f1e3a6fa  <=  Ic085f1faeb81e3027f909a7bd890d359[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibbee0996ea0f5e16b1f711345be7f2ae     <=
                                             I159df37fedc1447f6766308aa58ff70c[SGN_MAX_SUM_WDTH] ?
                                             ~I159df37fedc1447f6766308aa58ff70c + 1 :
                                             I159df37fedc1447f6766308aa58ff70c
                                             ;

            I446857735e680cae93a24dccb59b1924  <=  I159df37fedc1447f6766308aa58ff70c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idb777f1eb4c3cbba103b9b43f948ccf9     <=
                                             I53491740a9877fcff56e6a3d8ac61643[SGN_MAX_SUM_WDTH] ?
                                             ~I53491740a9877fcff56e6a3d8ac61643 + 1 :
                                             I53491740a9877fcff56e6a3d8ac61643
                                             ;

            I77b05a8aa92c66a235195a66dc13c0cc  <=  I53491740a9877fcff56e6a3d8ac61643[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id5e46b1f8844c7587f99d22170581a24     <=
                                             If9eba70be918197cc0bb2974f04c0687[SGN_MAX_SUM_WDTH] ?
                                             ~If9eba70be918197cc0bb2974f04c0687 + 1 :
                                             If9eba70be918197cc0bb2974f04c0687
                                             ;

            Ie92110d19f4886cdfcfacd0920c06a4e  <=  If9eba70be918197cc0bb2974f04c0687[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I67aadabd3cf49456cace7392a1e7a35a     <=
                                             I2a30d44d2006f17582bb431e397d3874[SGN_MAX_SUM_WDTH] ?
                                             ~I2a30d44d2006f17582bb431e397d3874 + 1 :
                                             I2a30d44d2006f17582bb431e397d3874
                                             ;

            I36ba87b69b5b9dd919319230f697dfad  <=  I2a30d44d2006f17582bb431e397d3874[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id5635595d6b7b6dd7e6d510a27ad6702     <=
                                             I4b64bd561b279a17da4758a188a2f395[SGN_MAX_SUM_WDTH] ?
                                             ~I4b64bd561b279a17da4758a188a2f395 + 1 :
                                             I4b64bd561b279a17da4758a188a2f395
                                             ;

            Id20e72ac258d1d1b6cdca1e6c9e3596d  <=  I4b64bd561b279a17da4758a188a2f395[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ice783314a4868f0bba8bc3c5e3b65ae4     <=
                                             I93d5297fada8dfdcffed4b7b56ef9c43[SGN_MAX_SUM_WDTH] ?
                                             ~I93d5297fada8dfdcffed4b7b56ef9c43 + 1 :
                                             I93d5297fada8dfdcffed4b7b56ef9c43
                                             ;

            Ifc34f5d6b7a7d0533439794958959856  <=  I93d5297fada8dfdcffed4b7b56ef9c43[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib2d9b7f58cf571b904be02e6073f9b94     <=
                                             Ic6e5118343e784f89cd1d3ba03309f20[SGN_MAX_SUM_WDTH] ?
                                             ~Ic6e5118343e784f89cd1d3ba03309f20 + 1 :
                                             Ic6e5118343e784f89cd1d3ba03309f20
                                             ;

            I849ee5d34760be03d4285185136aa52e  <=  Ic6e5118343e784f89cd1d3ba03309f20[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I61b6effae91ae4bdcce4550eb5cf0796     <=
                                             Ic5d76ee2f693c012e26dc17acb0086e2[SGN_MAX_SUM_WDTH] ?
                                             ~Ic5d76ee2f693c012e26dc17acb0086e2 + 1 :
                                             Ic5d76ee2f693c012e26dc17acb0086e2
                                             ;

            Ia3559d98eb372b7307f30ad1f7c4c7cd  <=  Ic5d76ee2f693c012e26dc17acb0086e2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If5cf6e81b0e3b77f6a45f2555201acc2     <=
                                             Id4ad545c42b5e4c8d5383568ad1e2013[SGN_MAX_SUM_WDTH] ?
                                             ~Id4ad545c42b5e4c8d5383568ad1e2013 + 1 :
                                             Id4ad545c42b5e4c8d5383568ad1e2013
                                             ;

            I7332e088bbff69db19c62685e033d26a  <=  Id4ad545c42b5e4c8d5383568ad1e2013[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I62fae5bf51588f28c3521715b834909d     <=
                                             I3a6030885679b87e44a54cdac13681ad[SGN_MAX_SUM_WDTH] ?
                                             ~I3a6030885679b87e44a54cdac13681ad + 1 :
                                             I3a6030885679b87e44a54cdac13681ad
                                             ;

            I44daa5992b00e7af19adbee70bf01f2b  <=  I3a6030885679b87e44a54cdac13681ad[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If5cbdab78a4cf86b6285a400d0e0ac90     <=
                                             I0791083d118ca9bf64108ec397af3d04[SGN_MAX_SUM_WDTH] ?
                                             ~I0791083d118ca9bf64108ec397af3d04 + 1 :
                                             I0791083d118ca9bf64108ec397af3d04
                                             ;

            Ie517386cb5832e406fefc5e85eb2e7d1  <=  I0791083d118ca9bf64108ec397af3d04[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6e481cc49441c08bcd9fdcabbe90a000     <=
                                             Ic683598c8ec40f18eed02cb89e8a8270[SGN_MAX_SUM_WDTH] ?
                                             ~Ic683598c8ec40f18eed02cb89e8a8270 + 1 :
                                             Ic683598c8ec40f18eed02cb89e8a8270
                                             ;

            I9b096ce09467c10f448496fda13987d2  <=  Ic683598c8ec40f18eed02cb89e8a8270[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3aa663be3dd604564ef68b9a2b9d7319     <=
                                             I1fc9bb5cc8d38dd67592141a4dbf2532[SGN_MAX_SUM_WDTH] ?
                                             ~I1fc9bb5cc8d38dd67592141a4dbf2532 + 1 :
                                             I1fc9bb5cc8d38dd67592141a4dbf2532
                                             ;

            If1c0a3726041f70e508d68cbf6e40e04  <=  I1fc9bb5cc8d38dd67592141a4dbf2532[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8031632ee8700c63c207e2d6a6bdb630     <=
                                             I7ec34dc5c899abcd284ccd637fccf4ba[SGN_MAX_SUM_WDTH] ?
                                             ~I7ec34dc5c899abcd284ccd637fccf4ba + 1 :
                                             I7ec34dc5c899abcd284ccd637fccf4ba
                                             ;

            Iaf36ce8598a29573979c683a5e2cf9fd  <=  I7ec34dc5c899abcd284ccd637fccf4ba[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9be2701858da0bdffbf2dff7bcfd7e1     <=
                                             I2d43f4939c3509b6e7e540d3da880c35[SGN_MAX_SUM_WDTH] ?
                                             ~I2d43f4939c3509b6e7e540d3da880c35 + 1 :
                                             I2d43f4939c3509b6e7e540d3da880c35
                                             ;

            Ice82cfe55a5f226746e59e5c8beb46be  <=  I2d43f4939c3509b6e7e540d3da880c35[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ief209532f4cbf1c6a41bea414577f825     <=
                                             I385df2a645f7269a298cbadc418a54b9[SGN_MAX_SUM_WDTH] ?
                                             ~I385df2a645f7269a298cbadc418a54b9 + 1 :
                                             I385df2a645f7269a298cbadc418a54b9
                                             ;

            Iea1297491d1dfe98f395d8c73808a893  <=  I385df2a645f7269a298cbadc418a54b9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1c8953ad3f64f3c3cc506808aad29dab     <=
                                             I5f90162de7034f414b502958f5ec9b3a[SGN_MAX_SUM_WDTH] ?
                                             ~I5f90162de7034f414b502958f5ec9b3a + 1 :
                                             I5f90162de7034f414b502958f5ec9b3a
                                             ;

            If43dd31198c8a0da6fabd194cf13bb70  <=  I5f90162de7034f414b502958f5ec9b3a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1b519d88bbf86cfb080a50ea0480a128     <=
                                             I74353ed1bcc55b22f5d1f406b5069eaa[SGN_MAX_SUM_WDTH] ?
                                             ~I74353ed1bcc55b22f5d1f406b5069eaa + 1 :
                                             I74353ed1bcc55b22f5d1f406b5069eaa
                                             ;

            Ibeb8c72b90b50c6897224ca1a792fa56  <=  I74353ed1bcc55b22f5d1f406b5069eaa[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5b8258f35d889071109216b464abb2a4     <=
                                             I6c28ab1bc42131e4ff3fa98c97990c37[SGN_MAX_SUM_WDTH] ?
                                             ~I6c28ab1bc42131e4ff3fa98c97990c37 + 1 :
                                             I6c28ab1bc42131e4ff3fa98c97990c37
                                             ;

            I8e87530a131b5a73cad6df68b9e4967f  <=  I6c28ab1bc42131e4ff3fa98c97990c37[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id9681d4e0e4d375f9279de115a4337a3     <=
                                             Ia7c2ca9384d0415bbfe92f719a8a4a2f[SGN_MAX_SUM_WDTH] ?
                                             ~Ia7c2ca9384d0415bbfe92f719a8a4a2f + 1 :
                                             Ia7c2ca9384d0415bbfe92f719a8a4a2f
                                             ;

            Idf8d15c7bd7705b9aafbda09c3a5b46c  <=  Ia7c2ca9384d0415bbfe92f719a8a4a2f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib42144ece00b82debd70011724a29c91     <=
                                             Ice3a20a00f8742bbf47a043b84964ee3[SGN_MAX_SUM_WDTH] ?
                                             ~Ice3a20a00f8742bbf47a043b84964ee3 + 1 :
                                             Ice3a20a00f8742bbf47a043b84964ee3
                                             ;

            I2aea17846a53e2eb2968581ee2c48226  <=  Ice3a20a00f8742bbf47a043b84964ee3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic5717058a1815f63f164de1b1defe8cb     <=
                                             I22bdaa7e1b37f335d3fb2232df587cfd[SGN_MAX_SUM_WDTH] ?
                                             ~I22bdaa7e1b37f335d3fb2232df587cfd + 1 :
                                             I22bdaa7e1b37f335d3fb2232df587cfd
                                             ;

            I169d8f2bb5fde5b202b4239b7a7f1ed5  <=  I22bdaa7e1b37f335d3fb2232df587cfd[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iea41672f012f225d64d9c75b198c812f     <=
                                             I1c41347158d76f8b81dfa334e99d07ed[SGN_MAX_SUM_WDTH] ?
                                             ~I1c41347158d76f8b81dfa334e99d07ed + 1 :
                                             I1c41347158d76f8b81dfa334e99d07ed
                                             ;

            I40a223380fb4414a3f26a08cb90025ec  <=  I1c41347158d76f8b81dfa334e99d07ed[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7a070bd014e1d2c5e55e5fcba88a5664     <=
                                             I3464039cbf8ed089ae1894998c1e156b[SGN_MAX_SUM_WDTH] ?
                                             ~I3464039cbf8ed089ae1894998c1e156b + 1 :
                                             I3464039cbf8ed089ae1894998c1e156b
                                             ;

            Ie117f6ec475f5d6444998af151ce4e69  <=  I3464039cbf8ed089ae1894998c1e156b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4a0a8b28429b708363458c74230b0fc2     <=
                                             Ie7409851212f99a429d94460669686b8[SGN_MAX_SUM_WDTH] ?
                                             ~Ie7409851212f99a429d94460669686b8 + 1 :
                                             Ie7409851212f99a429d94460669686b8
                                             ;

            If7f3174da35dd39af7f4792aaa649bf1  <=  Ie7409851212f99a429d94460669686b8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If585e4075ac1740f3b141ae6a50200f7     <=
                                             Ia575bcac8f127884a151a3a323763614[SGN_MAX_SUM_WDTH] ?
                                             ~Ia575bcac8f127884a151a3a323763614 + 1 :
                                             Ia575bcac8f127884a151a3a323763614
                                             ;

            I719a892ad54e63b217c7271741b29cc5  <=  Ia575bcac8f127884a151a3a323763614[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie1a68cf09bb21a1629369fde87f51bea     <=
                                             I2a193624be6cb259f18ece3546c7ad21[SGN_MAX_SUM_WDTH] ?
                                             ~I2a193624be6cb259f18ece3546c7ad21 + 1 :
                                             I2a193624be6cb259f18ece3546c7ad21
                                             ;

            I4acf6d84471cd237f65c9b2391b7a20c  <=  I2a193624be6cb259f18ece3546c7ad21[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I72b8547125d0ad6c1ad39a68b55c818c     <=
                                             If40ad1197633c486c3aadfa277f9ab51[SGN_MAX_SUM_WDTH] ?
                                             ~If40ad1197633c486c3aadfa277f9ab51 + 1 :
                                             If40ad1197633c486c3aadfa277f9ab51
                                             ;

            I7a387a1f887c32e9d0f8e89912a8618c  <=  If40ad1197633c486c3aadfa277f9ab51[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie14ba4a8657740f9a8d057258db2cb09     <=
                                             I629ddfee3e7d36b93b743e69b4c817d6[SGN_MAX_SUM_WDTH] ?
                                             ~I629ddfee3e7d36b93b743e69b4c817d6 + 1 :
                                             I629ddfee3e7d36b93b743e69b4c817d6
                                             ;

            Ib862ac63c230ccde7fae0e62f9d047fe  <=  I629ddfee3e7d36b93b743e69b4c817d6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I27490a69fb2a1f6f298639254c37cf9e     <=
                                             I3469ef81705fd1534d6e5eb194f1e4b4[SGN_MAX_SUM_WDTH] ?
                                             ~I3469ef81705fd1534d6e5eb194f1e4b4 + 1 :
                                             I3469ef81705fd1534d6e5eb194f1e4b4
                                             ;

            I8f1a8a22637d37c3692e808d5eb3d543  <=  I3469ef81705fd1534d6e5eb194f1e4b4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I49b9c212fbe74a5dd8b087e417296186     <=
                                             I832d0a2832b2c665f1261b07ac6f9f2f[SGN_MAX_SUM_WDTH] ?
                                             ~I832d0a2832b2c665f1261b07ac6f9f2f + 1 :
                                             I832d0a2832b2c665f1261b07ac6f9f2f
                                             ;

            I6f420c64640dfb0c001f57df7e3b4504  <=  I832d0a2832b2c665f1261b07ac6f9f2f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0a8e6f5cc8b6ea599b7605abe6479bec     <=
                                             I3c2aa289ff967b044d6a37f75f048ec8[SGN_MAX_SUM_WDTH] ?
                                             ~I3c2aa289ff967b044d6a37f75f048ec8 + 1 :
                                             I3c2aa289ff967b044d6a37f75f048ec8
                                             ;

            I3600031716c2b4e21c9f577d34e033dc  <=  I3c2aa289ff967b044d6a37f75f048ec8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib6d94b34d3886717e4016fec196f277f     <=
                                             Id2ea09c8febd9e18d231a5b069beb3cf[SGN_MAX_SUM_WDTH] ?
                                             ~Id2ea09c8febd9e18d231a5b069beb3cf + 1 :
                                             Id2ea09c8febd9e18d231a5b069beb3cf
                                             ;

            I002820a37fa7c6c504c487df4368e2cf  <=  Id2ea09c8febd9e18d231a5b069beb3cf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id7e53d36da7171e036ebfc984dbcea6e     <=
                                             I7b80623d743adcc50430ab9c8591ff29[SGN_MAX_SUM_WDTH] ?
                                             ~I7b80623d743adcc50430ab9c8591ff29 + 1 :
                                             I7b80623d743adcc50430ab9c8591ff29
                                             ;

            I8a4c1f23212ff846400651b100add502  <=  I7b80623d743adcc50430ab9c8591ff29[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2ec254d80fd0683d782302cf3839559b     <=
                                             I05750cd7c98f3c9726b8bbf5cdc76844[SGN_MAX_SUM_WDTH] ?
                                             ~I05750cd7c98f3c9726b8bbf5cdc76844 + 1 :
                                             I05750cd7c98f3c9726b8bbf5cdc76844
                                             ;

            Ice1ce5b4c30841dd92268559ebadafcf  <=  I05750cd7c98f3c9726b8bbf5cdc76844[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibbedaef61051d5df82cd6d55e05c80da     <=
                                             I389c717754a30812dc8ae3c8dffa20fb[SGN_MAX_SUM_WDTH] ?
                                             ~I389c717754a30812dc8ae3c8dffa20fb + 1 :
                                             I389c717754a30812dc8ae3c8dffa20fb
                                             ;

            I3eeeb1949945032d6c1759875426b733  <=  I389c717754a30812dc8ae3c8dffa20fb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I501336bb7ba172c05dd5840036e6228c     <=
                                             I8f151f04b124fa5023d7be59c9a43519[SGN_MAX_SUM_WDTH] ?
                                             ~I8f151f04b124fa5023d7be59c9a43519 + 1 :
                                             I8f151f04b124fa5023d7be59c9a43519
                                             ;

            I384d5377ee6b8f7eb2db23a2e444ddbc  <=  I8f151f04b124fa5023d7be59c9a43519[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8e5c4c6c63e42054359cee697cc0d026     <=
                                             I29a6f7a5b1c0bcc988363bee48b6cdc9[SGN_MAX_SUM_WDTH] ?
                                             ~I29a6f7a5b1c0bcc988363bee48b6cdc9 + 1 :
                                             I29a6f7a5b1c0bcc988363bee48b6cdc9
                                             ;

            I30d615203b697787ead37394953925cc  <=  I29a6f7a5b1c0bcc988363bee48b6cdc9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id3daa6db921871b752bf92366446afcc     <=
                                             If35ed918a1a2b59c5e0ba5f3e0a1a6f0[SGN_MAX_SUM_WDTH] ?
                                             ~If35ed918a1a2b59c5e0ba5f3e0a1a6f0 + 1 :
                                             If35ed918a1a2b59c5e0ba5f3e0a1a6f0
                                             ;

            Ib16548d471f0a4f4625852ea04335dcc  <=  If35ed918a1a2b59c5e0ba5f3e0a1a6f0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id8367ec60787bfad0da8aa76c6ed8ddb     <=
                                             I0816b1444f89b9c61ccfee1d16a72c1a[SGN_MAX_SUM_WDTH] ?
                                             ~I0816b1444f89b9c61ccfee1d16a72c1a + 1 :
                                             I0816b1444f89b9c61ccfee1d16a72c1a
                                             ;

            I0987c561670b7b2b6683303c1be39561  <=  I0816b1444f89b9c61ccfee1d16a72c1a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I533649312ec995f1f9e514c59a8675b1     <=
                                             I4a292e7bcef3cdaa716ceb101685471e[SGN_MAX_SUM_WDTH] ?
                                             ~I4a292e7bcef3cdaa716ceb101685471e + 1 :
                                             I4a292e7bcef3cdaa716ceb101685471e
                                             ;

            I2bdf4736022e5da7294a0e851006a124  <=  I4a292e7bcef3cdaa716ceb101685471e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0621d0b2c83e70b4afd65eb9dca4b514     <=
                                             I1d6b3fdfa7d64dc0761ebcb6ad076bff[SGN_MAX_SUM_WDTH] ?
                                             ~I1d6b3fdfa7d64dc0761ebcb6ad076bff + 1 :
                                             I1d6b3fdfa7d64dc0761ebcb6ad076bff
                                             ;

            Ic6fd9592d2ffcb8f4ca83c6f0bd19975  <=  I1d6b3fdfa7d64dc0761ebcb6ad076bff[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2ae01892a3cd0432618d7280b31daddb     <=
                                             I3ce8fb414e9fa103854658db43291eb0[SGN_MAX_SUM_WDTH] ?
                                             ~I3ce8fb414e9fa103854658db43291eb0 + 1 :
                                             I3ce8fb414e9fa103854658db43291eb0
                                             ;

            I14bf11ad80890227e47fda26ae1b9c24  <=  I3ce8fb414e9fa103854658db43291eb0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ed8a2f30bd2ea269341c2267ae3fe83     <=
                                             I01d190427900b3cef55d978630d6e035[SGN_MAX_SUM_WDTH] ?
                                             ~I01d190427900b3cef55d978630d6e035 + 1 :
                                             I01d190427900b3cef55d978630d6e035
                                             ;

            I8ca17b6cf35e1b1f8f601604575d3f27  <=  I01d190427900b3cef55d978630d6e035[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2c819e7f62c0dc0aac650074b203163b     <=
                                             I59a613f178a100a88f479d85e5f01cbf[SGN_MAX_SUM_WDTH] ?
                                             ~I59a613f178a100a88f479d85e5f01cbf + 1 :
                                             I59a613f178a100a88f479d85e5f01cbf
                                             ;

            I275cd09649a750edb8ae8313e4e1e279  <=  I59a613f178a100a88f479d85e5f01cbf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I30e20b58913d6fbe5817e1956ba8e570     <=
                                             Ife0377dc8109d89213ab27df5304e1e0[SGN_MAX_SUM_WDTH] ?
                                             ~Ife0377dc8109d89213ab27df5304e1e0 + 1 :
                                             Ife0377dc8109d89213ab27df5304e1e0
                                             ;

            I7d6a6026eb3c4d06e682523424f9628f  <=  Ife0377dc8109d89213ab27df5304e1e0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1b922bed7f3c4a6705f3ce7a885a68cd     <=
                                             Idb55c5acb92ff1b590670da114d3c668[SGN_MAX_SUM_WDTH] ?
                                             ~Idb55c5acb92ff1b590670da114d3c668 + 1 :
                                             Idb55c5acb92ff1b590670da114d3c668
                                             ;

            Ia0c192e590d8c914555b434ce5a634a8  <=  Idb55c5acb92ff1b590670da114d3c668[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2f65f0917713ecc8585392d3b557c1bf     <=
                                             Iefdc7b1d3aea42c3ddf9645510803a98[SGN_MAX_SUM_WDTH] ?
                                             ~Iefdc7b1d3aea42c3ddf9645510803a98 + 1 :
                                             Iefdc7b1d3aea42c3ddf9645510803a98
                                             ;

            Ic98c8641d2022080297c54ff2539e75d  <=  Iefdc7b1d3aea42c3ddf9645510803a98[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3301533e7d9e527118a67c462f1b4357     <=
                                             Ieae82f715fb1dc2d6d173f82b1547c35[SGN_MAX_SUM_WDTH] ?
                                             ~Ieae82f715fb1dc2d6d173f82b1547c35 + 1 :
                                             Ieae82f715fb1dc2d6d173f82b1547c35
                                             ;

            I87f34821cd0b58f8855b25c75f2dd32d  <=  Ieae82f715fb1dc2d6d173f82b1547c35[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I52a88bdb1f03da82730f7579b7b5305d     <=
                                             I18a9e19a2c41be29621e5da6a2b08e3e[SGN_MAX_SUM_WDTH] ?
                                             ~I18a9e19a2c41be29621e5da6a2b08e3e + 1 :
                                             I18a9e19a2c41be29621e5da6a2b08e3e
                                             ;

            I87211ac14d832ad3205d47fb83cf256a  <=  I18a9e19a2c41be29621e5da6a2b08e3e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I644c730662b3725d26cd46fb46106104     <=
                                             If4bfa23dd5ba282c7c9445769eb865f2[SGN_MAX_SUM_WDTH] ?
                                             ~If4bfa23dd5ba282c7c9445769eb865f2 + 1 :
                                             If4bfa23dd5ba282c7c9445769eb865f2
                                             ;

            Ib81431cfb3b281555fa7e5b4582a2524  <=  If4bfa23dd5ba282c7c9445769eb865f2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3da3e36c76c4123bec6879bccb39e933     <=
                                             Id9717e06ce4a9b03b8430559671918d7[SGN_MAX_SUM_WDTH] ?
                                             ~Id9717e06ce4a9b03b8430559671918d7 + 1 :
                                             Id9717e06ce4a9b03b8430559671918d7
                                             ;

            I835b902949c2c4c09b757d4d35574a76  <=  Id9717e06ce4a9b03b8430559671918d7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iebde55cddc8170f7dd8855ea55eff0ce     <=
                                             Ie54acd665004eec584ab9ff50df3961c[SGN_MAX_SUM_WDTH] ?
                                             ~Ie54acd665004eec584ab9ff50df3961c + 1 :
                                             Ie54acd665004eec584ab9ff50df3961c
                                             ;

            I8510240df7dc41f85ad58a39868a1fd7  <=  Ie54acd665004eec584ab9ff50df3961c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie673e2d92a7090b2fa1c5e14a2e03be3     <=
                                             I16c418af5cc92780b28cd56e8baa825a[SGN_MAX_SUM_WDTH] ?
                                             ~I16c418af5cc92780b28cd56e8baa825a + 1 :
                                             I16c418af5cc92780b28cd56e8baa825a
                                             ;

            I1b6abc8fbab3849b285e9f88a4fe867b  <=  I16c418af5cc92780b28cd56e8baa825a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If90afe75714f8660ad0eb9f9ea06cd6b     <=
                                             Iddb359180e3925dcf7081ba0560c27da[SGN_MAX_SUM_WDTH] ?
                                             ~Iddb359180e3925dcf7081ba0560c27da + 1 :
                                             Iddb359180e3925dcf7081ba0560c27da
                                             ;

            Ied638fee34f8baed4154b0b72e43a21e  <=  Iddb359180e3925dcf7081ba0560c27da[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifd96e3a6e0050c30a4308328cfecb21f     <=
                                             I354ac9e0f361928cf5cc7aaf22fd9622[SGN_MAX_SUM_WDTH] ?
                                             ~I354ac9e0f361928cf5cc7aaf22fd9622 + 1 :
                                             I354ac9e0f361928cf5cc7aaf22fd9622
                                             ;

            I14fa7aebb608d4a3d67176ba27d34d9a  <=  I354ac9e0f361928cf5cc7aaf22fd9622[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I68b92cc2d83e9a718edd2aea82314016     <=
                                             Ibf2b259738d54319e3af570db254a79f[SGN_MAX_SUM_WDTH] ?
                                             ~Ibf2b259738d54319e3af570db254a79f + 1 :
                                             Ibf2b259738d54319e3af570db254a79f
                                             ;

            Iad90879acba3fc2101829549264960f3  <=  Ibf2b259738d54319e3af570db254a79f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6bdbb92363f0e072ed04654e9aad17a5     <=
                                             I07150b2eb1a5818fe98aa210cb6e8221[SGN_MAX_SUM_WDTH] ?
                                             ~I07150b2eb1a5818fe98aa210cb6e8221 + 1 :
                                             I07150b2eb1a5818fe98aa210cb6e8221
                                             ;

            Ife0952b85f14a960007b67646b0cd969  <=  I07150b2eb1a5818fe98aa210cb6e8221[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I87a4267db59b97ef1b9bca8743cb0322     <=
                                             I5dea5fdbd4e09be8fd264360ae399b32[SGN_MAX_SUM_WDTH] ?
                                             ~I5dea5fdbd4e09be8fd264360ae399b32 + 1 :
                                             I5dea5fdbd4e09be8fd264360ae399b32
                                             ;

            If876ca6a14ffb4323503ed46666bc25f  <=  I5dea5fdbd4e09be8fd264360ae399b32[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I44eacb2bea725efab7c0dd560279f0f8     <=
                                             I9c52550c142c131371199bbf8bc08c01[SGN_MAX_SUM_WDTH] ?
                                             ~I9c52550c142c131371199bbf8bc08c01 + 1 :
                                             I9c52550c142c131371199bbf8bc08c01
                                             ;

            If2dfcbf493b761fb5d7c622e739b23f3  <=  I9c52550c142c131371199bbf8bc08c01[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I87a2736466c5ee62b7cc55f17e715ffa     <=
                                             I72d86068a1d9bdfe04f6ebe9afcf980f[SGN_MAX_SUM_WDTH] ?
                                             ~I72d86068a1d9bdfe04f6ebe9afcf980f + 1 :
                                             I72d86068a1d9bdfe04f6ebe9afcf980f
                                             ;

            I2c8f4a147b363d9c5ef0e080d9a9ed40  <=  I72d86068a1d9bdfe04f6ebe9afcf980f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7a66c7713ba126fdc24940cd92f7e10b     <=
                                             I412dfb474dbd41f407bbd57b0dd75a4e[SGN_MAX_SUM_WDTH] ?
                                             ~I412dfb474dbd41f407bbd57b0dd75a4e + 1 :
                                             I412dfb474dbd41f407bbd57b0dd75a4e
                                             ;

            I485f9d1104a965d5d035feef912a2ca8  <=  I412dfb474dbd41f407bbd57b0dd75a4e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1f11c579f34c41aade41c53f53468057     <=
                                             Ie759523643b0c4becb96025e66635b3b[SGN_MAX_SUM_WDTH] ?
                                             ~Ie759523643b0c4becb96025e66635b3b + 1 :
                                             Ie759523643b0c4becb96025e66635b3b
                                             ;

            I10fca5f2cbf5e2bc3433c0dda579a051  <=  Ie759523643b0c4becb96025e66635b3b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I651a438f70583d476ae10f066e035435     <=
                                             I1ef0aa04ba8b896c7ca95c10513b0ecf[SGN_MAX_SUM_WDTH] ?
                                             ~I1ef0aa04ba8b896c7ca95c10513b0ecf + 1 :
                                             I1ef0aa04ba8b896c7ca95c10513b0ecf
                                             ;

            If8572800d5d80cc92dd917b60447b63b  <=  I1ef0aa04ba8b896c7ca95c10513b0ecf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibdf17fa73794c846e15fe0a915b071e5     <=
                                             I880964445bdadb87455b7f8a865fa0e8[SGN_MAX_SUM_WDTH] ?
                                             ~I880964445bdadb87455b7f8a865fa0e8 + 1 :
                                             I880964445bdadb87455b7f8a865fa0e8
                                             ;

            I24645082ef16129eed1c574f5fc601ca  <=  I880964445bdadb87455b7f8a865fa0e8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I76d3221fbcefc0ee08655f7ba4919f3c     <=
                                             I145bec82b2f3234d2299ea32c9cd32ef[SGN_MAX_SUM_WDTH] ?
                                             ~I145bec82b2f3234d2299ea32c9cd32ef + 1 :
                                             I145bec82b2f3234d2299ea32c9cd32ef
                                             ;

            I207a0f6184a0b3be71766a8b47ea5535  <=  I145bec82b2f3234d2299ea32c9cd32ef[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3458f69c90ea8b20b3d1f67e9a13ec2e     <=
                                             Ib045b4ad82a55c17dd36f29467d49f36[SGN_MAX_SUM_WDTH] ?
                                             ~Ib045b4ad82a55c17dd36f29467d49f36 + 1 :
                                             Ib045b4ad82a55c17dd36f29467d49f36
                                             ;

            I5cac08dabbb6de3b01c821d4db93a8e3  <=  Ib045b4ad82a55c17dd36f29467d49f36[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia2d6e9e1e92a30c7028af50ddfbb9bf9     <=
                                             I7a195d3fb06596483191024720bfae2c[SGN_MAX_SUM_WDTH] ?
                                             ~I7a195d3fb06596483191024720bfae2c + 1 :
                                             I7a195d3fb06596483191024720bfae2c
                                             ;

            Ibe6b8c57d7ff47b6fdad5fadf1f6b841  <=  I7a195d3fb06596483191024720bfae2c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I66c91b5133d9812a03daecc0b14211f8     <=
                                             Ib84c4b8d94ce1e35ab220224ffedf4e5[SGN_MAX_SUM_WDTH] ?
                                             ~Ib84c4b8d94ce1e35ab220224ffedf4e5 + 1 :
                                             Ib84c4b8d94ce1e35ab220224ffedf4e5
                                             ;

            I477326720157df2503149125a43ee987  <=  Ib84c4b8d94ce1e35ab220224ffedf4e5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifb5986949e88167526d9fcfe07b417ca     <=
                                             Idd54eedf955c30f097484bd789eaa3d1[SGN_MAX_SUM_WDTH] ?
                                             ~Idd54eedf955c30f097484bd789eaa3d1 + 1 :
                                             Idd54eedf955c30f097484bd789eaa3d1
                                             ;

            I2c741a5fed7d88e9bdd6b7459feac649  <=  Idd54eedf955c30f097484bd789eaa3d1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedada801ca6cd173ee523ef335e91ff6     <=
                                             I123677fa899ce173a83101d91990014a[SGN_MAX_SUM_WDTH] ?
                                             ~I123677fa899ce173a83101d91990014a + 1 :
                                             I123677fa899ce173a83101d91990014a
                                             ;

            I17a6511072c7fb4846be5844decf17d6  <=  I123677fa899ce173a83101d91990014a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4e2722e547586da7565b2d91a7fc91e7     <=
                                             I26617d3c93a1f4069ee6fb732264d935[SGN_MAX_SUM_WDTH] ?
                                             ~I26617d3c93a1f4069ee6fb732264d935 + 1 :
                                             I26617d3c93a1f4069ee6fb732264d935
                                             ;

            I5ebc3047985651f4b9a957d502a97e95  <=  I26617d3c93a1f4069ee6fb732264d935[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib321a8ceda62c64ab25dc1c718301bda     <=
                                             I00410cf0d9a85b1fa2f70212bed15642[SGN_MAX_SUM_WDTH] ?
                                             ~I00410cf0d9a85b1fa2f70212bed15642 + 1 :
                                             I00410cf0d9a85b1fa2f70212bed15642
                                             ;

            Ifa09fc1b009d073d5a9973b430c63469  <=  I00410cf0d9a85b1fa2f70212bed15642[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I58daeebec4873e6c1c07c090ff81235c     <=
                                             I28f355e643584a4ab8d55777aa26fa78[SGN_MAX_SUM_WDTH] ?
                                             ~I28f355e643584a4ab8d55777aa26fa78 + 1 :
                                             I28f355e643584a4ab8d55777aa26fa78
                                             ;

            Ie6212a29c7c6b035cfff4c869f945b68  <=  I28f355e643584a4ab8d55777aa26fa78[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3f103fbbe49c86c9db46129bd4632cab     <=
                                             Id21bc865cd2de83bced952fb9c25f11a[SGN_MAX_SUM_WDTH] ?
                                             ~Id21bc865cd2de83bced952fb9c25f11a + 1 :
                                             Id21bc865cd2de83bced952fb9c25f11a
                                             ;

            If343015b4815b01dae88bbb6f2017b3d  <=  Id21bc865cd2de83bced952fb9c25f11a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id6697ca17f1bd6ddd112951b9d89a8ea     <=
                                             Ib6fbb4e2ef502ae86dc697dccfe035a8[SGN_MAX_SUM_WDTH] ?
                                             ~Ib6fbb4e2ef502ae86dc697dccfe035a8 + 1 :
                                             Ib6fbb4e2ef502ae86dc697dccfe035a8
                                             ;

            Ia0116a3cebf94318ed5b287960957ad6  <=  Ib6fbb4e2ef502ae86dc697dccfe035a8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I445ede2983c7470b4418a2ec0cbbd5e1     <=
                                             I2b0c304769c917cc6acc0855ada30c54[SGN_MAX_SUM_WDTH] ?
                                             ~I2b0c304769c917cc6acc0855ada30c54 + 1 :
                                             I2b0c304769c917cc6acc0855ada30c54
                                             ;

            Id75c23e80cdf25d883806ed20d4ae783  <=  I2b0c304769c917cc6acc0855ada30c54[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I034e56cd77ee400ed81b78177b202930     <=
                                             Iba61bc5c2e1230784d619375b7c756b4[SGN_MAX_SUM_WDTH] ?
                                             ~Iba61bc5c2e1230784d619375b7c756b4 + 1 :
                                             Iba61bc5c2e1230784d619375b7c756b4
                                             ;

            I1b43f29e0ddb72467befd6f3a9c1c829  <=  Iba61bc5c2e1230784d619375b7c756b4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I08edadbd9366786f96b44268d096b4aa     <=
                                             I613acad8a236e9deeb6967de9c067a48[SGN_MAX_SUM_WDTH] ?
                                             ~I613acad8a236e9deeb6967de9c067a48 + 1 :
                                             I613acad8a236e9deeb6967de9c067a48
                                             ;

            I3fd0fa3b774d30a267d61e9427d09f3f  <=  I613acad8a236e9deeb6967de9c067a48[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f86a7af86eb04c5df18e09888cdce7b     <=
                                             I427eb014c821ba5108aaa6ebbd8bc23c[SGN_MAX_SUM_WDTH] ?
                                             ~I427eb014c821ba5108aaa6ebbd8bc23c + 1 :
                                             I427eb014c821ba5108aaa6ebbd8bc23c
                                             ;

            I2eb08ebaa07a1004638cdd61a7209b7d  <=  I427eb014c821ba5108aaa6ebbd8bc23c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic00d037a11f8a27ab34e4daab8c9c2e6     <=
                                             I9b3fc0250b26e6faa2b7b44e863ff3f0[SGN_MAX_SUM_WDTH] ?
                                             ~I9b3fc0250b26e6faa2b7b44e863ff3f0 + 1 :
                                             I9b3fc0250b26e6faa2b7b44e863ff3f0
                                             ;

            I258c45897919cec5c6acaddee7f3a41b  <=  I9b3fc0250b26e6faa2b7b44e863ff3f0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4d95ceccc6c3ad37f13c98339c59e5c4     <=
                                             I79c12183f8bb94f4a3ce466570eadb80[SGN_MAX_SUM_WDTH] ?
                                             ~I79c12183f8bb94f4a3ce466570eadb80 + 1 :
                                             I79c12183f8bb94f4a3ce466570eadb80
                                             ;

            Ib42d37576e3aff3d205f1f8822cc58b5  <=  I79c12183f8bb94f4a3ce466570eadb80[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1ea967d377f462a0e06d7d0d4d95b342     <=
                                             Id4ba2f12931de7439cd52eb15b0241eb[SGN_MAX_SUM_WDTH] ?
                                             ~Id4ba2f12931de7439cd52eb15b0241eb + 1 :
                                             Id4ba2f12931de7439cd52eb15b0241eb
                                             ;

            I1c2ee281cd47a8414851c5e1c758ea65  <=  Id4ba2f12931de7439cd52eb15b0241eb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib0feec63123e66bd6ad6935e9b7fa6bf     <=
                                             I430558329b5398ffd51855414df8ba17[SGN_MAX_SUM_WDTH] ?
                                             ~I430558329b5398ffd51855414df8ba17 + 1 :
                                             I430558329b5398ffd51855414df8ba17
                                             ;

            Ie644d131c4f2c603e8e64c5581fdf822  <=  I430558329b5398ffd51855414df8ba17[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7d120060ddae9ff8f7206b3ef63eda50     <=
                                             I4eacf5b6fddf6cb1dad592392eeef166[SGN_MAX_SUM_WDTH] ?
                                             ~I4eacf5b6fddf6cb1dad592392eeef166 + 1 :
                                             I4eacf5b6fddf6cb1dad592392eeef166
                                             ;

            I9b76f0121a3f7e887e7121db50024ab4  <=  I4eacf5b6fddf6cb1dad592392eeef166[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib47f8f72386e2e65a88fbadd3a705225     <=
                                             I64921a58b87a14a3d6d02647f5c4a496[SGN_MAX_SUM_WDTH] ?
                                             ~I64921a58b87a14a3d6d02647f5c4a496 + 1 :
                                             I64921a58b87a14a3d6d02647f5c4a496
                                             ;

            I9eaf4e9ebe07717503ff69b51f0e1905  <=  I64921a58b87a14a3d6d02647f5c4a496[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4e0efc35346e2934f5bb4c34a4bc5f90     <=
                                             I9a93abf3585f9f937118adfdacdd8736[SGN_MAX_SUM_WDTH] ?
                                             ~I9a93abf3585f9f937118adfdacdd8736 + 1 :
                                             I9a93abf3585f9f937118adfdacdd8736
                                             ;

            Icb0841ecf142687c3aa23e68f01c927c  <=  I9a93abf3585f9f937118adfdacdd8736[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3ca1014802f58087e3434a1e0df19c01     <=
                                             Ib368c9afabdccf356ff389540397e3e9[SGN_MAX_SUM_WDTH] ?
                                             ~Ib368c9afabdccf356ff389540397e3e9 + 1 :
                                             Ib368c9afabdccf356ff389540397e3e9
                                             ;

            Ie8c0fac00a9de74870e59cbf9e87a39b  <=  Ib368c9afabdccf356ff389540397e3e9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I688a3879b7be1544e6f94b4221c03213     <=
                                             I939d31990dc2265d78b3d5b9a031f0df[SGN_MAX_SUM_WDTH] ?
                                             ~I939d31990dc2265d78b3d5b9a031f0df + 1 :
                                             I939d31990dc2265d78b3d5b9a031f0df
                                             ;

            Iae5d6faac1f5685cb1d400ee2b1d85e0  <=  I939d31990dc2265d78b3d5b9a031f0df[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic22988138610c8671ec342f65f34c7ae     <=
                                             I3ded8a67a0163feb95cafacb2c539412[SGN_MAX_SUM_WDTH] ?
                                             ~I3ded8a67a0163feb95cafacb2c539412 + 1 :
                                             I3ded8a67a0163feb95cafacb2c539412
                                             ;

            Ib62b02ddf0f57bee49838d19783ef6c3  <=  I3ded8a67a0163feb95cafacb2c539412[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b85fdd83569e5cbb7d71eed50cb32fd     <=
                                             I20c10afd04ed128ce31162ca3c1a89fa[SGN_MAX_SUM_WDTH] ?
                                             ~I20c10afd04ed128ce31162ca3c1a89fa + 1 :
                                             I20c10afd04ed128ce31162ca3c1a89fa
                                             ;

            Ibd59d0e5a062f149bd0e91ba76985a13  <=  I20c10afd04ed128ce31162ca3c1a89fa[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idf55390c11e5b41ebc2a28e0af109913     <=
                                             I71db9043fb2adee1e96818330469e51d[SGN_MAX_SUM_WDTH] ?
                                             ~I71db9043fb2adee1e96818330469e51d + 1 :
                                             I71db9043fb2adee1e96818330469e51d
                                             ;

            I876fdba97e755b74532f7ab191fbac14  <=  I71db9043fb2adee1e96818330469e51d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6b48935ea25672ee9a42f49eae9e519f     <=
                                             I64112bb2686f6348b7caaf3e0cf6a4aa[SGN_MAX_SUM_WDTH] ?
                                             ~I64112bb2686f6348b7caaf3e0cf6a4aa + 1 :
                                             I64112bb2686f6348b7caaf3e0cf6a4aa
                                             ;

            I8edf1a08ef943f06ee28771c6e140e28  <=  I64112bb2686f6348b7caaf3e0cf6a4aa[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6a9e6c39c20e45773dab7823a7ff9486     <=
                                             Ib4d8b49de697e1a70b07e76e836872b5[SGN_MAX_SUM_WDTH] ?
                                             ~Ib4d8b49de697e1a70b07e76e836872b5 + 1 :
                                             Ib4d8b49de697e1a70b07e76e836872b5
                                             ;

            I7e12ad8a8ef857e02f4563b2f3a7f0ca  <=  Ib4d8b49de697e1a70b07e76e836872b5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I42907182010c5889ddb7a700ead16525     <=
                                             I67dd716c2039d45a57fe94847cf2eef5[SGN_MAX_SUM_WDTH] ?
                                             ~I67dd716c2039d45a57fe94847cf2eef5 + 1 :
                                             I67dd716c2039d45a57fe94847cf2eef5
                                             ;

            I17b3a9df6752da6cc987e902e6bbad48  <=  I67dd716c2039d45a57fe94847cf2eef5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib6c26f3e3358cc2ed6fbda83eabd4bd3     <=
                                             I60558c2a8261a6c4a06491a95c40dfec[SGN_MAX_SUM_WDTH] ?
                                             ~I60558c2a8261a6c4a06491a95c40dfec + 1 :
                                             I60558c2a8261a6c4a06491a95c40dfec
                                             ;

            I487496233a32f657171b3789590d0522  <=  I60558c2a8261a6c4a06491a95c40dfec[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia50d85808790790450f87a5246874b3f     <=
                                             I37e4ed1440968cf86567341f4febf6a7[SGN_MAX_SUM_WDTH] ?
                                             ~I37e4ed1440968cf86567341f4febf6a7 + 1 :
                                             I37e4ed1440968cf86567341f4febf6a7
                                             ;

            Ie34534dfd435b3d1cf35e82ca71e83ba  <=  I37e4ed1440968cf86567341f4febf6a7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id4a1744702d7808a80bc40697c864765     <=
                                             I369a541788e6ec2dbf5a29a93b8e9379[SGN_MAX_SUM_WDTH] ?
                                             ~I369a541788e6ec2dbf5a29a93b8e9379 + 1 :
                                             I369a541788e6ec2dbf5a29a93b8e9379
                                             ;

            I0e8679271ba733bb87c44b6b9f0b6ed2  <=  I369a541788e6ec2dbf5a29a93b8e9379[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0cf3d2f3e6793a2dcf15949da16ad28d     <=
                                             I7fcf3847a6884d9e2cb216ac22cc6eea[SGN_MAX_SUM_WDTH] ?
                                             ~I7fcf3847a6884d9e2cb216ac22cc6eea + 1 :
                                             I7fcf3847a6884d9e2cb216ac22cc6eea
                                             ;

            Ic14760b65c6fe150c3c48e64389a41d8  <=  I7fcf3847a6884d9e2cb216ac22cc6eea[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I90bd9107f4c931fa1ccb92998ea8cdeb     <=
                                             Ifc34e5240f1440c3a0415cc944241208[SGN_MAX_SUM_WDTH] ?
                                             ~Ifc34e5240f1440c3a0415cc944241208 + 1 :
                                             Ifc34e5240f1440c3a0415cc944241208
                                             ;

            Ied6c684cdd280b41ffab93a026d27282  <=  Ifc34e5240f1440c3a0415cc944241208[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ida1c729e6bfcec2c31a92aa9002f2c68     <=
                                             I7e7a9c6ba8c0e7b945fc5cbc7def9c6b[SGN_MAX_SUM_WDTH] ?
                                             ~I7e7a9c6ba8c0e7b945fc5cbc7def9c6b + 1 :
                                             I7e7a9c6ba8c0e7b945fc5cbc7def9c6b
                                             ;

            Id0f4dbb72da33748d8baf723c5a32567  <=  I7e7a9c6ba8c0e7b945fc5cbc7def9c6b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib848feeccd0ea78ebc8ba8368534c3d1     <=
                                             I8ea9c190206ea186295c33528d45551c[SGN_MAX_SUM_WDTH] ?
                                             ~I8ea9c190206ea186295c33528d45551c + 1 :
                                             I8ea9c190206ea186295c33528d45551c
                                             ;

            Ib0bb71b1f8829347b3a9a7543f9dd964  <=  I8ea9c190206ea186295c33528d45551c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icc11970bbae3adcfa33a0e5dba3e78f4     <=
                                             I70f9d851136c9e8fb264fb43d6ebeb61[SGN_MAX_SUM_WDTH] ?
                                             ~I70f9d851136c9e8fb264fb43d6ebeb61 + 1 :
                                             I70f9d851136c9e8fb264fb43d6ebeb61
                                             ;

            I47cbb92d2284aef7b9e56e88f0ba6f7e  <=  I70f9d851136c9e8fb264fb43d6ebeb61[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I86bb4ef4bdd7af8861280ef30fbeeeea     <=
                                             Iea50b0ab0e00bfce47e6fdb129ea4cae[SGN_MAX_SUM_WDTH] ?
                                             ~Iea50b0ab0e00bfce47e6fdb129ea4cae + 1 :
                                             Iea50b0ab0e00bfce47e6fdb129ea4cae
                                             ;

            Ic69094123b75ae36e3e54f179a9f2cb5  <=  Iea50b0ab0e00bfce47e6fdb129ea4cae[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7e0c259c6c7bacdff5edc44a22e005ba     <=
                                             Ie74b8877e9a7df32f3f5674aab1300af[SGN_MAX_SUM_WDTH] ?
                                             ~Ie74b8877e9a7df32f3f5674aab1300af + 1 :
                                             Ie74b8877e9a7df32f3f5674aab1300af
                                             ;

            I07abbbd75d91018ac53f53e64cffafb9  <=  Ie74b8877e9a7df32f3f5674aab1300af[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I897ddba059b27f7ed009b0cb70cfb46f     <=
                                             Iaa3d8acf714f23e5059aa21cc1c36dd4[SGN_MAX_SUM_WDTH] ?
                                             ~Iaa3d8acf714f23e5059aa21cc1c36dd4 + 1 :
                                             Iaa3d8acf714f23e5059aa21cc1c36dd4
                                             ;

            Ib02268d5048c7c8e83118070e927453f  <=  Iaa3d8acf714f23e5059aa21cc1c36dd4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4496243eb0542a514b551b4d09bffd7d     <=
                                             Ic98698807ac6942eaa491de5a2a523c0[SGN_MAX_SUM_WDTH] ?
                                             ~Ic98698807ac6942eaa491de5a2a523c0 + 1 :
                                             Ic98698807ac6942eaa491de5a2a523c0
                                             ;

            Idc2a9c6dd8d2aa912548c918c8a488f4  <=  Ic98698807ac6942eaa491de5a2a523c0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic931fb08b2e8441321ebdeed84576a0d     <=
                                             I3579622172c0ccdf3eeb3bd490b2e6db[SGN_MAX_SUM_WDTH] ?
                                             ~I3579622172c0ccdf3eeb3bd490b2e6db + 1 :
                                             I3579622172c0ccdf3eeb3bd490b2e6db
                                             ;

            I5ad7eb9d3ce7c712515254f892d1670d  <=  I3579622172c0ccdf3eeb3bd490b2e6db[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ieb6af5390b98e893ee05a939c16d2ffd     <=
                                             I1369d79bd170cc9b7ed0352e0701261b[SGN_MAX_SUM_WDTH] ?
                                             ~I1369d79bd170cc9b7ed0352e0701261b + 1 :
                                             I1369d79bd170cc9b7ed0352e0701261b
                                             ;

            Ife25829fb3c5023b7d69bbaadf9cf77e  <=  I1369d79bd170cc9b7ed0352e0701261b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2a54bad4c5a8885dd24b8687c6db0de     <=
                                             I16196f7cfe21843797e1f3ef19b09048[SGN_MAX_SUM_WDTH] ?
                                             ~I16196f7cfe21843797e1f3ef19b09048 + 1 :
                                             I16196f7cfe21843797e1f3ef19b09048
                                             ;

            I8b2a79aa4ac88e6b4ca8188a7852022e  <=  I16196f7cfe21843797e1f3ef19b09048[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ecbad763d2b48b78a0584beaefc78ee     <=
                                             I20e403ad09d5eeb59020f7fe3b683432[SGN_MAX_SUM_WDTH] ?
                                             ~I20e403ad09d5eeb59020f7fe3b683432 + 1 :
                                             I20e403ad09d5eeb59020f7fe3b683432
                                             ;

            I081e2595b18f306a74d070203447ecf6  <=  I20e403ad09d5eeb59020f7fe3b683432[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I20556d23c873c71c7ebc8a961bf40251     <=
                                             I8d6ef29e41c3ef0fe66820e77c486591[SGN_MAX_SUM_WDTH] ?
                                             ~I8d6ef29e41c3ef0fe66820e77c486591 + 1 :
                                             I8d6ef29e41c3ef0fe66820e77c486591
                                             ;

            I68b152a599887c0039dd9d45c528c219  <=  I8d6ef29e41c3ef0fe66820e77c486591[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I79012e6351e6320c22437aa216ea4df1     <=
                                             I77fcee77b0cb1c65ca313526461231e4[SGN_MAX_SUM_WDTH] ?
                                             ~I77fcee77b0cb1c65ca313526461231e4 + 1 :
                                             I77fcee77b0cb1c65ca313526461231e4
                                             ;

            Id051f1d5454802e0eb37e22248efe8ca  <=  I77fcee77b0cb1c65ca313526461231e4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibf74ab9af877d27c3a6f3881f00ddaf1     <=
                                             I40c64a3c54b15800ed725dfce5144f17[SGN_MAX_SUM_WDTH] ?
                                             ~I40c64a3c54b15800ed725dfce5144f17 + 1 :
                                             I40c64a3c54b15800ed725dfce5144f17
                                             ;

            Ic4c6f707f461cebbc4c93f2ba664ae7b  <=  I40c64a3c54b15800ed725dfce5144f17[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I843d35db35d7b42a87ce78d3772cec2f     <=
                                             I57bddc5d3b9daf16fa9c2eaa3a148a03[SGN_MAX_SUM_WDTH] ?
                                             ~I57bddc5d3b9daf16fa9c2eaa3a148a03 + 1 :
                                             I57bddc5d3b9daf16fa9c2eaa3a148a03
                                             ;

            Ia538dadbd6ae3711740595a18c89b65d  <=  I57bddc5d3b9daf16fa9c2eaa3a148a03[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2b1398b4bfd374d7221b0a68da28e979     <=
                                             I5d3dc544f4e02f31e8dbc2b399afa89e[SGN_MAX_SUM_WDTH] ?
                                             ~I5d3dc544f4e02f31e8dbc2b399afa89e + 1 :
                                             I5d3dc544f4e02f31e8dbc2b399afa89e
                                             ;

            Ie7d9730b191781c78391141d95d4f8bd  <=  I5d3dc544f4e02f31e8dbc2b399afa89e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6f615d6e74b0c02f8e4265523ad16404     <=
                                             I0bc53eebdddc25c9c1423068bbe7a2a1[SGN_MAX_SUM_WDTH] ?
                                             ~I0bc53eebdddc25c9c1423068bbe7a2a1 + 1 :
                                             I0bc53eebdddc25c9c1423068bbe7a2a1
                                             ;

            I12f2f886517647044cc251861721bbb9  <=  I0bc53eebdddc25c9c1423068bbe7a2a1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iae8a98dd4a7cbfbc56c1404b6a2020af     <=
                                             I23429a89ac40e62e5b13ec75e348e432[SGN_MAX_SUM_WDTH] ?
                                             ~I23429a89ac40e62e5b13ec75e348e432 + 1 :
                                             I23429a89ac40e62e5b13ec75e348e432
                                             ;

            I615053b36a1851a06125e2ed5ec7f880  <=  I23429a89ac40e62e5b13ec75e348e432[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iad53375a54d01c559c74981bf279dfb5     <=
                                             I417ae67e3ed05fb6ac8b24bcba692a83[SGN_MAX_SUM_WDTH] ?
                                             ~I417ae67e3ed05fb6ac8b24bcba692a83 + 1 :
                                             I417ae67e3ed05fb6ac8b24bcba692a83
                                             ;

            Ifbc6aa14cd448bbe416897a3671ba857  <=  I417ae67e3ed05fb6ac8b24bcba692a83[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5db1307f922e0c742d7d9f3a79a4a4f3     <=
                                             I5edf732eb5451f0f84087b8ccccab387[SGN_MAX_SUM_WDTH] ?
                                             ~I5edf732eb5451f0f84087b8ccccab387 + 1 :
                                             I5edf732eb5451f0f84087b8ccccab387
                                             ;

            Ie596289582a73e37f78f4ca4cab21e3c  <=  I5edf732eb5451f0f84087b8ccccab387[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9f78172ed5bf73752196f9a8810005f3     <=
                                             I26833c93cc1b8be86febb45560ae4707[SGN_MAX_SUM_WDTH] ?
                                             ~I26833c93cc1b8be86febb45560ae4707 + 1 :
                                             I26833c93cc1b8be86febb45560ae4707
                                             ;

            Ifad8c7bacf72583f91be27fbe5b7a1e1  <=  I26833c93cc1b8be86febb45560ae4707[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If85a22d670d47f491dd7568d0453ba1d     <=
                                             Iab7fe9d9176e8ceb00b7d04116dc0236[SGN_MAX_SUM_WDTH] ?
                                             ~Iab7fe9d9176e8ceb00b7d04116dc0236 + 1 :
                                             Iab7fe9d9176e8ceb00b7d04116dc0236
                                             ;

            Ie74c72742807ae4243748fd27d80d626  <=  Iab7fe9d9176e8ceb00b7d04116dc0236[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9e529170b2896e930a839295796fd31     <=
                                             Ie66e4f53df7e0bb44442a3c74883ab30[SGN_MAX_SUM_WDTH] ?
                                             ~Ie66e4f53df7e0bb44442a3c74883ab30 + 1 :
                                             Ie66e4f53df7e0bb44442a3c74883ab30
                                             ;

            Ie7a68c2b368a295f95571bc4a109b9f1  <=  Ie66e4f53df7e0bb44442a3c74883ab30[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7af536846bac40c1f221d1f72c6c25c     <=
                                             I591dd226d239200c681a1aac16849d31[SGN_MAX_SUM_WDTH] ?
                                             ~I591dd226d239200c681a1aac16849d31 + 1 :
                                             I591dd226d239200c681a1aac16849d31
                                             ;

            Id88a7edf897eea1b4a137141789a04f5  <=  I591dd226d239200c681a1aac16849d31[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib0eb61a2cb831dd35ce9850994e7c2da     <=
                                             Ic572d19feb1b9d45cb81aa0aeee01340[SGN_MAX_SUM_WDTH] ?
                                             ~Ic572d19feb1b9d45cb81aa0aeee01340 + 1 :
                                             Ic572d19feb1b9d45cb81aa0aeee01340
                                             ;

            Ib13436ad16a37d656d6b1ee95b9aee20  <=  Ic572d19feb1b9d45cb81aa0aeee01340[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I89d338f59960af7a47595d6afa206abc     <=
                                             I31306ed55c012f4e3f3da72bc404d6ba[SGN_MAX_SUM_WDTH] ?
                                             ~I31306ed55c012f4e3f3da72bc404d6ba + 1 :
                                             I31306ed55c012f4e3f3da72bc404d6ba
                                             ;

            Idc07dc30c0a957e474546ac7a60df38f  <=  I31306ed55c012f4e3f3da72bc404d6ba[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib3c1176eb8991e3e85855a9fe845c303     <=
                                             I374c888e91b747a2a6b58649c4a1969b[SGN_MAX_SUM_WDTH] ?
                                             ~I374c888e91b747a2a6b58649c4a1969b + 1 :
                                             I374c888e91b747a2a6b58649c4a1969b
                                             ;

            I595665d8128bb87ab62741d7ac520a4b  <=  I374c888e91b747a2a6b58649c4a1969b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I93073d05d509b821a743998cf32c58ee     <=
                                             Ic71fea427a788b416d088a44f2600c51[SGN_MAX_SUM_WDTH] ?
                                             ~Ic71fea427a788b416d088a44f2600c51 + 1 :
                                             Ic71fea427a788b416d088a44f2600c51
                                             ;

            I256050251d23250854ff337bef28e460  <=  Ic71fea427a788b416d088a44f2600c51[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iab6dac1909c1564c3890ffecc13418df     <=
                                             Ib6fec22f8466773bb13224a90a4e3c2d[SGN_MAX_SUM_WDTH] ?
                                             ~Ib6fec22f8466773bb13224a90a4e3c2d + 1 :
                                             Ib6fec22f8466773bb13224a90a4e3c2d
                                             ;

            I82f0e5a32d1bcd761a74f1f9ce8c88ba  <=  Ib6fec22f8466773bb13224a90a4e3c2d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1b75eeb29167a171d89f6e67039436d5     <=
                                             Id30dc8c00fd07e9ad68a8fc3c740557f[SGN_MAX_SUM_WDTH] ?
                                             ~Id30dc8c00fd07e9ad68a8fc3c740557f + 1 :
                                             Id30dc8c00fd07e9ad68a8fc3c740557f
                                             ;

            I98febac90cccb5fc1f3d966b6e38c4d3  <=  Id30dc8c00fd07e9ad68a8fc3c740557f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3a31adc52a1405555017b2ddf219b407     <=
                                             I85777d4d61b8e6fc99706bbe7fbfad8c[SGN_MAX_SUM_WDTH] ?
                                             ~I85777d4d61b8e6fc99706bbe7fbfad8c + 1 :
                                             I85777d4d61b8e6fc99706bbe7fbfad8c
                                             ;

            Ib534288c2cf976b6ec85db743bc2a823  <=  I85777d4d61b8e6fc99706bbe7fbfad8c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iaadba89c6a370240fc0758029f7d8db0     <=
                                             I707e0745e78aef8c802c0fd5a7b58ae5[SGN_MAX_SUM_WDTH] ?
                                             ~I707e0745e78aef8c802c0fd5a7b58ae5 + 1 :
                                             I707e0745e78aef8c802c0fd5a7b58ae5
                                             ;

            If988b82b86db1f4ff6d3695f7b0197e4  <=  I707e0745e78aef8c802c0fd5a7b58ae5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4f4a64fb3ced7d9f7ee4513178e9655a     <=
                                             I513c23daa981e69789b074975a589954[SGN_MAX_SUM_WDTH] ?
                                             ~I513c23daa981e69789b074975a589954 + 1 :
                                             I513c23daa981e69789b074975a589954
                                             ;

            I6ef260ef75e47b011a46ba2080ac3684  <=  I513c23daa981e69789b074975a589954[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0c76ca58f69c91758e755cd581241284     <=
                                             I3b0ea0ad1bf5f5820e582b0c1f97d949[SGN_MAX_SUM_WDTH] ?
                                             ~I3b0ea0ad1bf5f5820e582b0c1f97d949 + 1 :
                                             I3b0ea0ad1bf5f5820e582b0c1f97d949
                                             ;

            Ifc1da524e7670772834d521a6fc4c96f  <=  I3b0ea0ad1bf5f5820e582b0c1f97d949[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2312bce18958346149c868846e04643b     <=
                                             I857759675a04284a230c6e09e993db26[SGN_MAX_SUM_WDTH] ?
                                             ~I857759675a04284a230c6e09e993db26 + 1 :
                                             I857759675a04284a230c6e09e993db26
                                             ;

            I852d5295a32984af00c95f6d9389555e  <=  I857759675a04284a230c6e09e993db26[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3e154098cb0a48f1c23234f46613f406     <=
                                             I943326eaa918c39cb3fe412c77d8b131[SGN_MAX_SUM_WDTH] ?
                                             ~I943326eaa918c39cb3fe412c77d8b131 + 1 :
                                             I943326eaa918c39cb3fe412c77d8b131
                                             ;

            I3c0a621dbef864fd1f566bc2e47f32c6  <=  I943326eaa918c39cb3fe412c77d8b131[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1645c1c588bcbf15dd62d47e08b8e139     <=
                                             I9dcf55a3343d214ab70cbde50a34da4d[SGN_MAX_SUM_WDTH] ?
                                             ~I9dcf55a3343d214ab70cbde50a34da4d + 1 :
                                             I9dcf55a3343d214ab70cbde50a34da4d
                                             ;

            Ic04828ba2db8239b093043c27476d345  <=  I9dcf55a3343d214ab70cbde50a34da4d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4c25de66590e1745d37112e08d8c8e2c     <=
                                             I1fe6a30dcbcbdcfc0b3d6bbe38e9c3bc[SGN_MAX_SUM_WDTH] ?
                                             ~I1fe6a30dcbcbdcfc0b3d6bbe38e9c3bc + 1 :
                                             I1fe6a30dcbcbdcfc0b3d6bbe38e9c3bc
                                             ;

            I319012bc6fe93d78de57bcace0caaef5  <=  I1fe6a30dcbcbdcfc0b3d6bbe38e9c3bc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia03092ac621b8dd1c206fea1e8b0215f     <=
                                             I39216b818931b9d2fb6a93e5eda743aa[SGN_MAX_SUM_WDTH] ?
                                             ~I39216b818931b9d2fb6a93e5eda743aa + 1 :
                                             I39216b818931b9d2fb6a93e5eda743aa
                                             ;

            Ibb35bace971548c9fc98d773d1aff712  <=  I39216b818931b9d2fb6a93e5eda743aa[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5c9bdb033436dc9f6069baca31f24c2d     <=
                                             I24238e5bba0bf63288ad44c5dd3545f3[SGN_MAX_SUM_WDTH] ?
                                             ~I24238e5bba0bf63288ad44c5dd3545f3 + 1 :
                                             I24238e5bba0bf63288ad44c5dd3545f3
                                             ;

            I90023493600924a76d2192080cf6194e  <=  I24238e5bba0bf63288ad44c5dd3545f3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f07cf4865480f18ad6945974ec2231c     <=
                                             Ic0a34c6b56cc30ddec7e5b755e18a27d[SGN_MAX_SUM_WDTH] ?
                                             ~Ic0a34c6b56cc30ddec7e5b755e18a27d + 1 :
                                             Ic0a34c6b56cc30ddec7e5b755e18a27d
                                             ;

            Ia9f5ce4603af279bbd9b486b67016482  <=  Ic0a34c6b56cc30ddec7e5b755e18a27d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4a7119e8862fe4a6a4100dd9ac67dd24     <=
                                             I45e63318c784a30395ca1bbc692d1402[SGN_MAX_SUM_WDTH] ?
                                             ~I45e63318c784a30395ca1bbc692d1402 + 1 :
                                             I45e63318c784a30395ca1bbc692d1402
                                             ;

            I05721e06a1acdcc0571907c7d853f18c  <=  I45e63318c784a30395ca1bbc692d1402[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id78fcfc6724a05f46d44d7c3e7d0c756     <=
                                             Iae0e9a6d88b4fba34944cd2f0dd5c9ed[SGN_MAX_SUM_WDTH] ?
                                             ~Iae0e9a6d88b4fba34944cd2f0dd5c9ed + 1 :
                                             Iae0e9a6d88b4fba34944cd2f0dd5c9ed
                                             ;

            Ibfcfd3151af0d82bfce293ada44059b3  <=  Iae0e9a6d88b4fba34944cd2f0dd5c9ed[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7cbd9d619623cbabf8ed6b1fece8f012     <=
                                             I91d8bc9088850978c17bfa5f0bf93b26[SGN_MAX_SUM_WDTH] ?
                                             ~I91d8bc9088850978c17bfa5f0bf93b26 + 1 :
                                             I91d8bc9088850978c17bfa5f0bf93b26
                                             ;

            I9539fcc40d26b13015a864718b116d5b  <=  I91d8bc9088850978c17bfa5f0bf93b26[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I58951165d251e370b0f3b3fb537aed18     <=
                                             I014cecda30cbc4e25a1265a65ed0f0d4[SGN_MAX_SUM_WDTH] ?
                                             ~I014cecda30cbc4e25a1265a65ed0f0d4 + 1 :
                                             I014cecda30cbc4e25a1265a65ed0f0d4
                                             ;

            I5490039998187a1a2efc3549e3dee7d6  <=  I014cecda30cbc4e25a1265a65ed0f0d4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I21daac106f526d84cb8fa5239c19499d     <=
                                             I845250d1ee6395d022a0a20698eea330[SGN_MAX_SUM_WDTH] ?
                                             ~I845250d1ee6395d022a0a20698eea330 + 1 :
                                             I845250d1ee6395d022a0a20698eea330
                                             ;

            I2b97a79c90f6578c8b2f321f8d598cc8  <=  I845250d1ee6395d022a0a20698eea330[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I178029cec3a5d6141abdfa91b91fdbf4     <=
                                             I5d36a24496d96371aba3f0407c21e34d[SGN_MAX_SUM_WDTH] ?
                                             ~I5d36a24496d96371aba3f0407c21e34d + 1 :
                                             I5d36a24496d96371aba3f0407c21e34d
                                             ;

            I0c616f736879c28a5222de3d6f49a587  <=  I5d36a24496d96371aba3f0407c21e34d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I96dfb2efbb55a644616e3474ed07c364     <=
                                             If2f7a871f45dc098b3ebe056153235c7[SGN_MAX_SUM_WDTH] ?
                                             ~If2f7a871f45dc098b3ebe056153235c7 + 1 :
                                             If2f7a871f45dc098b3ebe056153235c7
                                             ;

            I5590d801fd7fb496019d4c31b7c6d898  <=  If2f7a871f45dc098b3ebe056153235c7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7a17d8f0e2d16c441044db68ee037731     <=
                                             Ib49df5d97f0ba140b6ec5f80aae719d6[SGN_MAX_SUM_WDTH] ?
                                             ~Ib49df5d97f0ba140b6ec5f80aae719d6 + 1 :
                                             Ib49df5d97f0ba140b6ec5f80aae719d6
                                             ;

            I27e1d2e0e980216b27b90ea48c061025  <=  Ib49df5d97f0ba140b6ec5f80aae719d6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2ced9bb3ae6bdc5b5ef2865fb46abf07     <=
                                             Ib25900518732253ccc4800716f3d772d[SGN_MAX_SUM_WDTH] ?
                                             ~Ib25900518732253ccc4800716f3d772d + 1 :
                                             Ib25900518732253ccc4800716f3d772d
                                             ;

            I474f6bd977f4197742d0bddb3bece684  <=  Ib25900518732253ccc4800716f3d772d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I89a93384020d93cf4d26b3902e06cd9e     <=
                                             I9d9b410818773fca2bc21ed678683369[SGN_MAX_SUM_WDTH] ?
                                             ~I9d9b410818773fca2bc21ed678683369 + 1 :
                                             I9d9b410818773fca2bc21ed678683369
                                             ;

            Iaa1e981134f5a5c02983c49562683bc5  <=  I9d9b410818773fca2bc21ed678683369[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibbb47d29b9a45559c13ffa3b046c66f5     <=
                                             Ia003b700205a0b2faf1cefa2c85c4df0[SGN_MAX_SUM_WDTH] ?
                                             ~Ia003b700205a0b2faf1cefa2c85c4df0 + 1 :
                                             Ia003b700205a0b2faf1cefa2c85c4df0
                                             ;

            Ib051eb1091a85f85a1e50007f1b27cab  <=  Ia003b700205a0b2faf1cefa2c85c4df0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0034177eb1049577a3578b371527f34b     <=
                                             I3b98b4efc159ac3eb3c7ea322459b666[SGN_MAX_SUM_WDTH] ?
                                             ~I3b98b4efc159ac3eb3c7ea322459b666 + 1 :
                                             I3b98b4efc159ac3eb3c7ea322459b666
                                             ;

            I6b5645cdde4b35a16fe3e91d90caaa4e  <=  I3b98b4efc159ac3eb3c7ea322459b666[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I22d9ea7bb5a1a3405bcd04b9af40fa62     <=
                                             Ibfe30b79869ff3125c248f623c494d09[SGN_MAX_SUM_WDTH] ?
                                             ~Ibfe30b79869ff3125c248f623c494d09 + 1 :
                                             Ibfe30b79869ff3125c248f623c494d09
                                             ;

            I8850ab26807dcd55fefadf6310729ca7  <=  Ibfe30b79869ff3125c248f623c494d09[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8a632e7a911bf5726fee587189cb6f16     <=
                                             Ice88c3ab21612bbd46676c650d9f4dbc[SGN_MAX_SUM_WDTH] ?
                                             ~Ice88c3ab21612bbd46676c650d9f4dbc + 1 :
                                             Ice88c3ab21612bbd46676c650d9f4dbc
                                             ;

            Ic5cb81c821716a8aabf8cc2283ff73ba  <=  Ice88c3ab21612bbd46676c650d9f4dbc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3765afc490b34e8a310998a4ebcff8cb     <=
                                             Ideadf767ef2ab66a1495ead1806ffe47[SGN_MAX_SUM_WDTH] ?
                                             ~Ideadf767ef2ab66a1495ead1806ffe47 + 1 :
                                             Ideadf767ef2ab66a1495ead1806ffe47
                                             ;

            I9a6923c6368526a53ef70e16471386ef  <=  Ideadf767ef2ab66a1495ead1806ffe47[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7607e800ae46a96e016b303120da4247     <=
                                             I28749b0f4f83f99b9082f7004e72aa70[SGN_MAX_SUM_WDTH] ?
                                             ~I28749b0f4f83f99b9082f7004e72aa70 + 1 :
                                             I28749b0f4f83f99b9082f7004e72aa70
                                             ;

            I620b8ecdcaccc1ec80ebcf9fa6af0017  <=  I28749b0f4f83f99b9082f7004e72aa70[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29b2f1fddee5e32f217d25410bcfce4f     <=
                                             I71ef3d84207d8995c13e88c16a0bacf8[SGN_MAX_SUM_WDTH] ?
                                             ~I71ef3d84207d8995c13e88c16a0bacf8 + 1 :
                                             I71ef3d84207d8995c13e88c16a0bacf8
                                             ;

            I141cda06bae0c5666e3bc61c6fe5ad66  <=  I71ef3d84207d8995c13e88c16a0bacf8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iba5f8a31a81f6aa06f5e38c03dc6db54     <=
                                             I630979d7924b3c17fe0aeaa04507ed03[SGN_MAX_SUM_WDTH] ?
                                             ~I630979d7924b3c17fe0aeaa04507ed03 + 1 :
                                             I630979d7924b3c17fe0aeaa04507ed03
                                             ;

            Ia9c273b32d0701c7f185ab2de9e57829  <=  I630979d7924b3c17fe0aeaa04507ed03[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifcb5c907ad503331317599e4e0ce7be8     <=
                                             I50a84fa93d73bfe0287f3297707b1901[SGN_MAX_SUM_WDTH] ?
                                             ~I50a84fa93d73bfe0287f3297707b1901 + 1 :
                                             I50a84fa93d73bfe0287f3297707b1901
                                             ;

            Ic3fb524ab434e80b3289c9241b65d224  <=  I50a84fa93d73bfe0287f3297707b1901[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I62d6f2ab4ec8b6ecfa544ad4d90eb30b     <=
                                             I19d6383f6319e9ed4b4f16fdf7a40cef[SGN_MAX_SUM_WDTH] ?
                                             ~I19d6383f6319e9ed4b4f16fdf7a40cef + 1 :
                                             I19d6383f6319e9ed4b4f16fdf7a40cef
                                             ;

            I23c8b64e433af0bd00cef44e38df99f8  <=  I19d6383f6319e9ed4b4f16fdf7a40cef[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ide65414c51b3cb182c0f2f238903d60a     <=
                                             I3515fa4f304e4b1537c612ca0212b4bc[SGN_MAX_SUM_WDTH] ?
                                             ~I3515fa4f304e4b1537c612ca0212b4bc + 1 :
                                             I3515fa4f304e4b1537c612ca0212b4bc
                                             ;

            If6a5dc79c0f6ce348956286737a369d8  <=  I3515fa4f304e4b1537c612ca0212b4bc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I03a8dc2288eaeb619e746990e20cc868     <=
                                             Ia154b83a5a01bf0ea74fcc873e45d980[SGN_MAX_SUM_WDTH] ?
                                             ~Ia154b83a5a01bf0ea74fcc873e45d980 + 1 :
                                             Ia154b83a5a01bf0ea74fcc873e45d980
                                             ;

            I34e6e9d2153e4a70ee36ab85e72d5318  <=  Ia154b83a5a01bf0ea74fcc873e45d980[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id81c1b44d16ddbcd466382c60fe84986     <=
                                             If021572d95ea7fcbae1454447dbbe212[SGN_MAX_SUM_WDTH] ?
                                             ~If021572d95ea7fcbae1454447dbbe212 + 1 :
                                             If021572d95ea7fcbae1454447dbbe212
                                             ;

            Ifdabf743a8cb46b7053000ff48ea0c60  <=  If021572d95ea7fcbae1454447dbbe212[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I503d72f4a2fd20dbf35aa27321d2ede7     <=
                                             Ib6c860f3146839d2c0e925007ac02d67[SGN_MAX_SUM_WDTH] ?
                                             ~Ib6c860f3146839d2c0e925007ac02d67 + 1 :
                                             Ib6c860f3146839d2c0e925007ac02d67
                                             ;

            I22f5bb821a2571d1764978fd76c8f1d0  <=  Ib6c860f3146839d2c0e925007ac02d67[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id6595a4cf33062d1f05cbcee2d0685f1     <=
                                             I21ae48e98044dcc69386800f72cc5fb7[SGN_MAX_SUM_WDTH] ?
                                             ~I21ae48e98044dcc69386800f72cc5fb7 + 1 :
                                             I21ae48e98044dcc69386800f72cc5fb7
                                             ;

            I1b695aa715615662eff7065c742b0859  <=  I21ae48e98044dcc69386800f72cc5fb7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I83ebdd7331ca8fbcf5250851b346c0b0     <=
                                             I4f436764c02c61027d89854865770734[SGN_MAX_SUM_WDTH] ?
                                             ~I4f436764c02c61027d89854865770734 + 1 :
                                             I4f436764c02c61027d89854865770734
                                             ;

            Iec91b3ca3b54010755d57f8b8ea4a544  <=  I4f436764c02c61027d89854865770734[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7f6ea26cdfe5986065e7b5aa6842cc1c     <=
                                             If213a0715834eb56c9c8862dcd643f36[SGN_MAX_SUM_WDTH] ?
                                             ~If213a0715834eb56c9c8862dcd643f36 + 1 :
                                             If213a0715834eb56c9c8862dcd643f36
                                             ;

            I06ad520cb02e46d34c45f207d42a9243  <=  If213a0715834eb56c9c8862dcd643f36[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idab1ec32c20f93c4cc1acb38158f92d5     <=
                                             If1eced44ede97a4e0ec55c26df8d6935[SGN_MAX_SUM_WDTH] ?
                                             ~If1eced44ede97a4e0ec55c26df8d6935 + 1 :
                                             If1eced44ede97a4e0ec55c26df8d6935
                                             ;

            I9d18ff3465afd8cae63abba68487542e  <=  If1eced44ede97a4e0ec55c26df8d6935[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0738add83419502e73674ded2f1ad6c7     <=
                                             Ibe579be01c1b2925be397ab7d202c200[SGN_MAX_SUM_WDTH] ?
                                             ~Ibe579be01c1b2925be397ab7d202c200 + 1 :
                                             Ibe579be01c1b2925be397ab7d202c200
                                             ;

            I914dedc1d5e5e21c9b8d07ec0ecc01f9  <=  Ibe579be01c1b2925be397ab7d202c200[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6c93e63a8e5a2dbd598f1565c7323b39     <=
                                             I675731b8fceb36c9a103803dea3700bc[SGN_MAX_SUM_WDTH] ?
                                             ~I675731b8fceb36c9a103803dea3700bc + 1 :
                                             I675731b8fceb36c9a103803dea3700bc
                                             ;

            I3375fff5ee0d4b4b12c5a70fbdee59fe  <=  I675731b8fceb36c9a103803dea3700bc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4aa57a9d46371f1680d5f95596f60b5d     <=
                                             I01374171f18d419d149433d7c789f1ef[SGN_MAX_SUM_WDTH] ?
                                             ~I01374171f18d419d149433d7c789f1ef + 1 :
                                             I01374171f18d419d149433d7c789f1ef
                                             ;

            Ia8e304ca12c82e41cb8e4de7be199394  <=  I01374171f18d419d149433d7c789f1ef[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5369a7203b78951a3c006c2d3b22507c     <=
                                             I9f66291cd8f80896cf27fa0b8382f465[SGN_MAX_SUM_WDTH] ?
                                             ~I9f66291cd8f80896cf27fa0b8382f465 + 1 :
                                             I9f66291cd8f80896cf27fa0b8382f465
                                             ;

            I3566f2779e860008b1a5d305366a07c9  <=  I9f66291cd8f80896cf27fa0b8382f465[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie72a79a6966cf198687b7c8a8bcdeb13     <=
                                             I73341b7d2d30f5fe7ce2d8659331de3b[SGN_MAX_SUM_WDTH] ?
                                             ~I73341b7d2d30f5fe7ce2d8659331de3b + 1 :
                                             I73341b7d2d30f5fe7ce2d8659331de3b
                                             ;

            Ie68b31360c12a83c6095254b6f14603c  <=  I73341b7d2d30f5fe7ce2d8659331de3b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie917ae4c44ab0f9c2f1747ff0d2a754e     <=
                                             Ieb9c6cc947f6e0429770118119be79e1[SGN_MAX_SUM_WDTH] ?
                                             ~Ieb9c6cc947f6e0429770118119be79e1 + 1 :
                                             Ieb9c6cc947f6e0429770118119be79e1
                                             ;

            I42ae0c42360c977b35429ce290516a6f  <=  Ieb9c6cc947f6e0429770118119be79e1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b1a31ccb34a742552c11b1945e23dd8     <=
                                             I2c58e39ab3b79963fa0eddc7180070dc[SGN_MAX_SUM_WDTH] ?
                                             ~I2c58e39ab3b79963fa0eddc7180070dc + 1 :
                                             I2c58e39ab3b79963fa0eddc7180070dc
                                             ;

            Ibe01835305315fab50269c72ef849b61  <=  I2c58e39ab3b79963fa0eddc7180070dc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9a65a845cf2eced39050e8481665f557     <=
                                             I789b342281d9ed8dbc03af5c0c508062[SGN_MAX_SUM_WDTH] ?
                                             ~I789b342281d9ed8dbc03af5c0c508062 + 1 :
                                             I789b342281d9ed8dbc03af5c0c508062
                                             ;

            Id806a2df1c4519bbbe811791cb4072f9  <=  I789b342281d9ed8dbc03af5c0c508062[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3b402b35d38a9fde312c89b82297c1a5     <=
                                             I95b62a2fcb0af75048d095dde733ddbc[SGN_MAX_SUM_WDTH] ?
                                             ~I95b62a2fcb0af75048d095dde733ddbc + 1 :
                                             I95b62a2fcb0af75048d095dde733ddbc
                                             ;

            Ifb70a30f8bade95f402e71f95fe6644b  <=  I95b62a2fcb0af75048d095dde733ddbc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I309fa33562370e339c19e2377e6a6a7a     <=
                                             I1e9d61b53dd7ce47230b341cc1b4e8b4[SGN_MAX_SUM_WDTH] ?
                                             ~I1e9d61b53dd7ce47230b341cc1b4e8b4 + 1 :
                                             I1e9d61b53dd7ce47230b341cc1b4e8b4
                                             ;

            I592a495aecc800236c3470ff8e6adbb5  <=  I1e9d61b53dd7ce47230b341cc1b4e8b4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7d06aed81222a030837cad2074c68e19     <=
                                             If5d6db7c002ad813677ca165380839b0[SGN_MAX_SUM_WDTH] ?
                                             ~If5d6db7c002ad813677ca165380839b0 + 1 :
                                             If5d6db7c002ad813677ca165380839b0
                                             ;

            I1c8024aa9d81704d2dcf63e34853f8cf  <=  If5d6db7c002ad813677ca165380839b0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I835cc6af0cd8189035f2441c2e0d3100     <=
                                             I0f7ceff0b6160697dbd097293de15156[SGN_MAX_SUM_WDTH] ?
                                             ~I0f7ceff0b6160697dbd097293de15156 + 1 :
                                             I0f7ceff0b6160697dbd097293de15156
                                             ;

            Ief03713f5cf37200373a20d42c7fc9eb  <=  I0f7ceff0b6160697dbd097293de15156[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If6f768d12f04087246a0d65de1aef99b     <=
                                             I2e142efe8de226e1a283576d1ae9ced9[SGN_MAX_SUM_WDTH] ?
                                             ~I2e142efe8de226e1a283576d1ae9ced9 + 1 :
                                             I2e142efe8de226e1a283576d1ae9ced9
                                             ;

            Ic3cb34aae74c5f1a870b3635f8a40764  <=  I2e142efe8de226e1a283576d1ae9ced9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie4b180e1e2cadb865b0eaf6509f99dbb     <=
                                             I88e4b172c1b5c2733bf050fa442964ce[SGN_MAX_SUM_WDTH] ?
                                             ~I88e4b172c1b5c2733bf050fa442964ce + 1 :
                                             I88e4b172c1b5c2733bf050fa442964ce
                                             ;

            Ifa3df8b249467cc1e827c69925ef415f  <=  I88e4b172c1b5c2733bf050fa442964ce[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie329a11fc3f6f59f6f1790612fde3250     <=
                                             Ie1f997dc210ff90c7ff78737d1240c30[SGN_MAX_SUM_WDTH] ?
                                             ~Ie1f997dc210ff90c7ff78737d1240c30 + 1 :
                                             Ie1f997dc210ff90c7ff78737d1240c30
                                             ;

            Icf3ad912aaeaa0c5cd1ab0edb898d6e8  <=  Ie1f997dc210ff90c7ff78737d1240c30[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idb7ddbee4076f7bf49177e69f5e4d112     <=
                                             I31307a02f9909905fd672eeaf54422a6[SGN_MAX_SUM_WDTH] ?
                                             ~I31307a02f9909905fd672eeaf54422a6 + 1 :
                                             I31307a02f9909905fd672eeaf54422a6
                                             ;

            Ib774f380e3d7cfd1f5f064e93d8134b4  <=  I31307a02f9909905fd672eeaf54422a6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I614d66a7dca2d08efdfdc157ca803d5c     <=
                                             I1e2dbb3cd67d96f046b39fd52947ff4e[SGN_MAX_SUM_WDTH] ?
                                             ~I1e2dbb3cd67d96f046b39fd52947ff4e + 1 :
                                             I1e2dbb3cd67d96f046b39fd52947ff4e
                                             ;

            Ic07c650e6e49892a41cfaf3a37471426  <=  I1e2dbb3cd67d96f046b39fd52947ff4e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iea16eb0ab70ebb1bc47ae55e11ced62d     <=
                                             Icad3b8650e3c4b3a425e1a1c7da14c1a[SGN_MAX_SUM_WDTH] ?
                                             ~Icad3b8650e3c4b3a425e1a1c7da14c1a + 1 :
                                             Icad3b8650e3c4b3a425e1a1c7da14c1a
                                             ;

            Ib1073489d63ea33d7f3892f4ff875358  <=  Icad3b8650e3c4b3a425e1a1c7da14c1a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifa8db43284d5bbebaed4f72d65cf9f92     <=
                                             I40acfb6473e56562b5bc1e7bfdeed8a6[SGN_MAX_SUM_WDTH] ?
                                             ~I40acfb6473e56562b5bc1e7bfdeed8a6 + 1 :
                                             I40acfb6473e56562b5bc1e7bfdeed8a6
                                             ;

            I174b6c36f2af82f8047cc76543a3b4ee  <=  I40acfb6473e56562b5bc1e7bfdeed8a6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I365d9f3e8b2a9890427f07386deeb093     <=
                                             I06a6d7c6a5be68cb75d83b2d8a1d3217[SGN_MAX_SUM_WDTH] ?
                                             ~I06a6d7c6a5be68cb75d83b2d8a1d3217 + 1 :
                                             I06a6d7c6a5be68cb75d83b2d8a1d3217
                                             ;

            I953b975a89adcc88039284970e9b3404  <=  I06a6d7c6a5be68cb75d83b2d8a1d3217[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I466aaa0b6cde2ade1901797b8c11e32c     <=
                                             I3d3ebea1cf84cec93ff60459177fdd18[SGN_MAX_SUM_WDTH] ?
                                             ~I3d3ebea1cf84cec93ff60459177fdd18 + 1 :
                                             I3d3ebea1cf84cec93ff60459177fdd18
                                             ;

            If2b40d249c531e10cc22d1335f350441  <=  I3d3ebea1cf84cec93ff60459177fdd18[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7057e329a65ab240ed6cfa824307af65     <=
                                             I59868ed1411b6439564cc73edf55297d[SGN_MAX_SUM_WDTH] ?
                                             ~I59868ed1411b6439564cc73edf55297d + 1 :
                                             I59868ed1411b6439564cc73edf55297d
                                             ;

            I44ccc3ae897109dd51f9afeef93daca4  <=  I59868ed1411b6439564cc73edf55297d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I624e50e3457d33d12680eaf8e7c34aa3     <=
                                             I97ae3d6c75edf1fd87347a8fd50fd27d[SGN_MAX_SUM_WDTH] ?
                                             ~I97ae3d6c75edf1fd87347a8fd50fd27d + 1 :
                                             I97ae3d6c75edf1fd87347a8fd50fd27d
                                             ;

            Ie9236599cea94cfb603c6b977fdbb44a  <=  I97ae3d6c75edf1fd87347a8fd50fd27d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9f356fd6820c33fdb5baff05a781e192     <=
                                             If98ad7df6cb49466733052834b458bb1[SGN_MAX_SUM_WDTH] ?
                                             ~If98ad7df6cb49466733052834b458bb1 + 1 :
                                             If98ad7df6cb49466733052834b458bb1
                                             ;

            I25f1ee9cee4d04bd8fec1fe601d016d7  <=  If98ad7df6cb49466733052834b458bb1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I39b9c7c664fe7017731877d145d55b44     <=
                                             I2ea63dcc06519b46da5b70cf36b68c76[SGN_MAX_SUM_WDTH] ?
                                             ~I2ea63dcc06519b46da5b70cf36b68c76 + 1 :
                                             I2ea63dcc06519b46da5b70cf36b68c76
                                             ;

            I5ec1e530b9007a75a778af4d82ab427b  <=  I2ea63dcc06519b46da5b70cf36b68c76[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic62ffbb9e58e0d08b0dec24bba1dc6f2     <=
                                             I979c3adad47ed2b8488aa7beaab7a565[SGN_MAX_SUM_WDTH] ?
                                             ~I979c3adad47ed2b8488aa7beaab7a565 + 1 :
                                             I979c3adad47ed2b8488aa7beaab7a565
                                             ;

            I8a9e516aa824260998d10db758642bb0  <=  I979c3adad47ed2b8488aa7beaab7a565[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8da2a532288fb817e7dc0cb7b4e3761c     <=
                                             Idc93f47a3946c69fc0c956ec3e4d4c28[SGN_MAX_SUM_WDTH] ?
                                             ~Idc93f47a3946c69fc0c956ec3e4d4c28 + 1 :
                                             Idc93f47a3946c69fc0c956ec3e4d4c28
                                             ;

            I70dd1350d65155ee7b562f4c79024a3d  <=  Idc93f47a3946c69fc0c956ec3e4d4c28[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6a6e559f5c98f846014e8107fea5a5d9     <=
                                             I3d57c80540bbdb043ce47c688950fd18[SGN_MAX_SUM_WDTH] ?
                                             ~I3d57c80540bbdb043ce47c688950fd18 + 1 :
                                             I3d57c80540bbdb043ce47c688950fd18
                                             ;

            Ic9146d8b3dd0c612073b70b8a8791e8c  <=  I3d57c80540bbdb043ce47c688950fd18[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibef9219f577b1a62dfdd77296fbfb24d     <=
                                             Id2083cbcf2aaa813c72071314c13ae6f[SGN_MAX_SUM_WDTH] ?
                                             ~Id2083cbcf2aaa813c72071314c13ae6f + 1 :
                                             Id2083cbcf2aaa813c72071314c13ae6f
                                             ;

            I857d3155df0b6dd704514b039c66fa97  <=  Id2083cbcf2aaa813c72071314c13ae6f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I52e6688b5bfff75529d18e20b22832ce     <=
                                             Iea95f61532bffc857f39331b244188d0[SGN_MAX_SUM_WDTH] ?
                                             ~Iea95f61532bffc857f39331b244188d0 + 1 :
                                             Iea95f61532bffc857f39331b244188d0
                                             ;

            Idc1b8aa2f81a7fbd87e4f5821d14bf01  <=  Iea95f61532bffc857f39331b244188d0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iff22c49354eefca0ea3c5959c14b782c     <=
                                             I42dd514d52d448707c7dcc5c799ee7f1[SGN_MAX_SUM_WDTH] ?
                                             ~I42dd514d52d448707c7dcc5c799ee7f1 + 1 :
                                             I42dd514d52d448707c7dcc5c799ee7f1
                                             ;

            I68b585571699a57bc6ba5e8955467119  <=  I42dd514d52d448707c7dcc5c799ee7f1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie5377bbdb4111ed00356d5b7737102f3     <=
                                             Ib6ee76ae9fed974530f73fb401405e27[SGN_MAX_SUM_WDTH] ?
                                             ~Ib6ee76ae9fed974530f73fb401405e27 + 1 :
                                             Ib6ee76ae9fed974530f73fb401405e27
                                             ;

            Ib70e99c3acc76286a6811bcacc9284de  <=  Ib6ee76ae9fed974530f73fb401405e27[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I55bf0f3379a8c44634b8f0a3d06c049e     <=
                                             I3aea3d7d9965e4cde24ba83120af804e[SGN_MAX_SUM_WDTH] ?
                                             ~I3aea3d7d9965e4cde24ba83120af804e + 1 :
                                             I3aea3d7d9965e4cde24ba83120af804e
                                             ;

            Iee17ece482d04964d3c21a092ec955a4  <=  I3aea3d7d9965e4cde24ba83120af804e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9bc9541607f4f6aedb686cdde297bcda     <=
                                             I3b1550f5b3e421d44005a01b0075bf33[SGN_MAX_SUM_WDTH] ?
                                             ~I3b1550f5b3e421d44005a01b0075bf33 + 1 :
                                             I3b1550f5b3e421d44005a01b0075bf33
                                             ;

            I5a247475beb737d470f03507e55f5b24  <=  I3b1550f5b3e421d44005a01b0075bf33[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia4620554fbb1d81a71a15a846e4be2f5     <=
                                             I00bc9cf3ab66e198dd7bf2cc930aa2c5[SGN_MAX_SUM_WDTH] ?
                                             ~I00bc9cf3ab66e198dd7bf2cc930aa2c5 + 1 :
                                             I00bc9cf3ab66e198dd7bf2cc930aa2c5
                                             ;

            I13b0c9578f7b6b3b7e6704d7b44079c4  <=  I00bc9cf3ab66e198dd7bf2cc930aa2c5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibb31b35388ba8ba2ecf98449308ee67d     <=
                                             I79d4eac1731095e588b7003d1c83aba7[SGN_MAX_SUM_WDTH] ?
                                             ~I79d4eac1731095e588b7003d1c83aba7 + 1 :
                                             I79d4eac1731095e588b7003d1c83aba7
                                             ;

            I41eff06fe1dea8be4613945de596d3ca  <=  I79d4eac1731095e588b7003d1c83aba7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia20410fb3d56587f89a54c00b943b305     <=
                                             I6512194d646b949c1f8037e3911a8720[SGN_MAX_SUM_WDTH] ?
                                             ~I6512194d646b949c1f8037e3911a8720 + 1 :
                                             I6512194d646b949c1f8037e3911a8720
                                             ;

            I08f22261d5713c0636d77c7938f592d6  <=  I6512194d646b949c1f8037e3911a8720[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9d268f3da12e35b9a4229b7340c0f018     <=
                                             Ief2dcb1d14d5065729e66207068d0519[SGN_MAX_SUM_WDTH] ?
                                             ~Ief2dcb1d14d5065729e66207068d0519 + 1 :
                                             Ief2dcb1d14d5065729e66207068d0519
                                             ;

            I1c7e41b9cb1bdb6f649c88c0ed3f4100  <=  Ief2dcb1d14d5065729e66207068d0519[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2fce29bd666082eedb2fb3ec8b5ae4dd     <=
                                             Ib343818dd2f04189d56a6fc40c8da197[SGN_MAX_SUM_WDTH] ?
                                             ~Ib343818dd2f04189d56a6fc40c8da197 + 1 :
                                             Ib343818dd2f04189d56a6fc40c8da197
                                             ;

            Idd59a5357d4c835379ed180ac0924bf1  <=  Ib343818dd2f04189d56a6fc40c8da197[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia1e8b61e2579a90f5c88ded11c7322c2     <=
                                             Ie38501f8b5cd9e64ed80bed953adbb48[SGN_MAX_SUM_WDTH] ?
                                             ~Ie38501f8b5cd9e64ed80bed953adbb48 + 1 :
                                             Ie38501f8b5cd9e64ed80bed953adbb48
                                             ;

            Ibe7e5c2cb9c50eca34a3859d13e83a92  <=  Ie38501f8b5cd9e64ed80bed953adbb48[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8cf3718ba65b7fed72e3955f190e34d1     <=
                                             Id50a8c0b1739857f19228131b51f7937[SGN_MAX_SUM_WDTH] ?
                                             ~Id50a8c0b1739857f19228131b51f7937 + 1 :
                                             Id50a8c0b1739857f19228131b51f7937
                                             ;

            Ibf5c141c5cc0a6a20c05b52bf8282476  <=  Id50a8c0b1739857f19228131b51f7937[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7e802d300af54d394b4ee041798c0513     <=
                                             I8946d670fb58546b8854b34dad0e8430[SGN_MAX_SUM_WDTH] ?
                                             ~I8946d670fb58546b8854b34dad0e8430 + 1 :
                                             I8946d670fb58546b8854b34dad0e8430
                                             ;

            I0038305f94aaefe2cd1a243580d95932  <=  I8946d670fb58546b8854b34dad0e8430[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id4fd5a4b97cfa1e176a26f3a823c5516     <=
                                             I122129edde3336f22ba613499bfabfc0[SGN_MAX_SUM_WDTH] ?
                                             ~I122129edde3336f22ba613499bfabfc0 + 1 :
                                             I122129edde3336f22ba613499bfabfc0
                                             ;

            I5364deb983adc2ae505ed2b8c57f876d  <=  I122129edde3336f22ba613499bfabfc0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icbf8d4e75fc66c05eb49c5075696fb07     <=
                                             I2ce23daae62346911511cfea5bed788f[SGN_MAX_SUM_WDTH] ?
                                             ~I2ce23daae62346911511cfea5bed788f + 1 :
                                             I2ce23daae62346911511cfea5bed788f
                                             ;

            Ifdb5589982db805a0416e1c01276249a  <=  I2ce23daae62346911511cfea5bed788f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I746a7e90adb2f213b75ae12a161aca0d     <=
                                             I5496ff29bde6957c01c5d7e5f2d8cbac[SGN_MAX_SUM_WDTH] ?
                                             ~I5496ff29bde6957c01c5d7e5f2d8cbac + 1 :
                                             I5496ff29bde6957c01c5d7e5f2d8cbac
                                             ;

            I8bb5522183b65583fda83067990b3e94  <=  I5496ff29bde6957c01c5d7e5f2d8cbac[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icb1029aaaaed8c698862ea9c5e22132c     <=
                                             I66fe45afee3cd240ed3ef77262387f40[SGN_MAX_SUM_WDTH] ?
                                             ~I66fe45afee3cd240ed3ef77262387f40 + 1 :
                                             I66fe45afee3cd240ed3ef77262387f40
                                             ;

            I1e77fe6aeaba852aba34ed37dd53add6  <=  I66fe45afee3cd240ed3ef77262387f40[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib93ea7028c172373b53cdafecae32a67     <=
                                             Id08a0b67ee6d6e08628238b1e5ac0dc8[SGN_MAX_SUM_WDTH] ?
                                             ~Id08a0b67ee6d6e08628238b1e5ac0dc8 + 1 :
                                             Id08a0b67ee6d6e08628238b1e5ac0dc8
                                             ;

            I9171019227f35760d02d0c8ce786f4d3  <=  Id08a0b67ee6d6e08628238b1e5ac0dc8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9628275b000e418f3903daebfdace92     <=
                                             I2b94a5c3e2ee6f13fae5ec588be73ba0[SGN_MAX_SUM_WDTH] ?
                                             ~I2b94a5c3e2ee6f13fae5ec588be73ba0 + 1 :
                                             I2b94a5c3e2ee6f13fae5ec588be73ba0
                                             ;

            I6e92a48aaab94074a555efa9bd1e7243  <=  I2b94a5c3e2ee6f13fae5ec588be73ba0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I830202fb6f08f98c7f71893a881bd555     <=
                                             I8b6ce93d2c7b309d4d043e938ef6cb12[SGN_MAX_SUM_WDTH] ?
                                             ~I8b6ce93d2c7b309d4d043e938ef6cb12 + 1 :
                                             I8b6ce93d2c7b309d4d043e938ef6cb12
                                             ;

            I3bc094d67805664859fdcb66f1360e64  <=  I8b6ce93d2c7b309d4d043e938ef6cb12[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6f38bc9359562f57c1603355e9ee312b     <=
                                             I46d88449ca1db5f462e0442932bc5f53[SGN_MAX_SUM_WDTH] ?
                                             ~I46d88449ca1db5f462e0442932bc5f53 + 1 :
                                             I46d88449ca1db5f462e0442932bc5f53
                                             ;

            I2518ccf385b3b677d95983bc550282e8  <=  I46d88449ca1db5f462e0442932bc5f53[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4701b732d59c26e3790a63c1936f9a24     <=
                                             I402417fdf22d1b9e08e905e3206a6edc[SGN_MAX_SUM_WDTH] ?
                                             ~I402417fdf22d1b9e08e905e3206a6edc + 1 :
                                             I402417fdf22d1b9e08e905e3206a6edc
                                             ;

            I7547c56b32513ad45d775b4502596d9d  <=  I402417fdf22d1b9e08e905e3206a6edc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib5d28d8f73d17ab6df6a1291e50c04ab     <=
                                             I287e3042873300b74530542044f57277[SGN_MAX_SUM_WDTH] ?
                                             ~I287e3042873300b74530542044f57277 + 1 :
                                             I287e3042873300b74530542044f57277
                                             ;

            I013d84bfd582acc7accf07ec522961fa  <=  I287e3042873300b74530542044f57277[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I81259f391db792339824ad5dd1a0057b     <=
                                             I4c6118afff7012ebdec7b6168f1ba067[SGN_MAX_SUM_WDTH] ?
                                             ~I4c6118afff7012ebdec7b6168f1ba067 + 1 :
                                             I4c6118afff7012ebdec7b6168f1ba067
                                             ;

            I0ec27b590ee6dcdd9c1086105e3b6c23  <=  I4c6118afff7012ebdec7b6168f1ba067[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6f09ac63effe67a86798b9b4e1690664     <=
                                             I444e2151e66af9ec6c1e984ad706b7a0[SGN_MAX_SUM_WDTH] ?
                                             ~I444e2151e66af9ec6c1e984ad706b7a0 + 1 :
                                             I444e2151e66af9ec6c1e984ad706b7a0
                                             ;

            I4cdc955fa9afc75c2c977de4ec540e1e  <=  I444e2151e66af9ec6c1e984ad706b7a0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I370b4b3a0048a93ba374a40e170c75a3     <=
                                             I3c800d94a189c70fb956298deb686700[SGN_MAX_SUM_WDTH] ?
                                             ~I3c800d94a189c70fb956298deb686700 + 1 :
                                             I3c800d94a189c70fb956298deb686700
                                             ;

            Ieefbb5d6f4ac1e586832c5c0f513c5a2  <=  I3c800d94a189c70fb956298deb686700[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3f8476d0aa0ea2439b67ea1a4adf36c5     <=
                                             I0b3393ffccd4b2a9b42a68f185b074f8[SGN_MAX_SUM_WDTH] ?
                                             ~I0b3393ffccd4b2a9b42a68f185b074f8 + 1 :
                                             I0b3393ffccd4b2a9b42a68f185b074f8
                                             ;

            Ic828cdd5dfde844df4c150921af2a443  <=  I0b3393ffccd4b2a9b42a68f185b074f8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35b52dba10a8a5b22b518388fecac82d     <=
                                             Ie1996578a600cbb605703974fcd3494a[SGN_MAX_SUM_WDTH] ?
                                             ~Ie1996578a600cbb605703974fcd3494a + 1 :
                                             Ie1996578a600cbb605703974fcd3494a
                                             ;

            Idf1ecab26889c4adcb835fda6b1cb368  <=  Ie1996578a600cbb605703974fcd3494a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic7db274ed18e6fdecf30381a31238777     <=
                                             Ib912bf53b3fc6753b228a488d9d25520[SGN_MAX_SUM_WDTH] ?
                                             ~Ib912bf53b3fc6753b228a488d9d25520 + 1 :
                                             Ib912bf53b3fc6753b228a488d9d25520
                                             ;

            I00d3f14b20e1ea7d726533386e0eba27  <=  Ib912bf53b3fc6753b228a488d9d25520[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2c4e538a8db759e9799541d9178ec61e     <=
                                             I77f81eeb736f7ad4abcd88fa9b952bc0[SGN_MAX_SUM_WDTH] ?
                                             ~I77f81eeb736f7ad4abcd88fa9b952bc0 + 1 :
                                             I77f81eeb736f7ad4abcd88fa9b952bc0
                                             ;

            I7f720a18542528f0c9bfb14f699ff4da  <=  I77f81eeb736f7ad4abcd88fa9b952bc0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ief6d4c3f5ef8663e111ef99347b023f5     <=
                                             Ic09db56c2b021b09e0cf4fe501f2a5ec[SGN_MAX_SUM_WDTH] ?
                                             ~Ic09db56c2b021b09e0cf4fe501f2a5ec + 1 :
                                             Ic09db56c2b021b09e0cf4fe501f2a5ec
                                             ;

            Ia98a6f01e4eb5bc74d50d350e79be426  <=  Ic09db56c2b021b09e0cf4fe501f2a5ec[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id95e964e5faecb52c72669b0d28a4bf5     <=
                                             I576cf92938eb1c168e0f9ee1b6bf0be7[SGN_MAX_SUM_WDTH] ?
                                             ~I576cf92938eb1c168e0f9ee1b6bf0be7 + 1 :
                                             I576cf92938eb1c168e0f9ee1b6bf0be7
                                             ;

            I182b43872d50de6f7afb700f178b160e  <=  I576cf92938eb1c168e0f9ee1b6bf0be7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0fcef4538102ac6d24aa7090d5405afa     <=
                                             Ia1d7ca394ee29ff9cc463c525fbf7947[SGN_MAX_SUM_WDTH] ?
                                             ~Ia1d7ca394ee29ff9cc463c525fbf7947 + 1 :
                                             Ia1d7ca394ee29ff9cc463c525fbf7947
                                             ;

            Ic9b72b2a91d951cf08cf54ed215ecaa8  <=  Ia1d7ca394ee29ff9cc463c525fbf7947[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I055019e38eec6badd1739033d43d7d97     <=
                                             I7fff588b55c99166b13cd816d6a5c166[SGN_MAX_SUM_WDTH] ?
                                             ~I7fff588b55c99166b13cd816d6a5c166 + 1 :
                                             I7fff588b55c99166b13cd816d6a5c166
                                             ;

            I93084ccf5b5e4efaee968b497bb2a775  <=  I7fff588b55c99166b13cd816d6a5c166[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I35c20a6e823da77a870b421eef2e0a95     <=
                                             I755d06b657ce02dabc6dbb6d44e619e6[SGN_MAX_SUM_WDTH] ?
                                             ~I755d06b657ce02dabc6dbb6d44e619e6 + 1 :
                                             I755d06b657ce02dabc6dbb6d44e619e6
                                             ;

            Id38852415486e6989b89a0d85ad6771b  <=  I755d06b657ce02dabc6dbb6d44e619e6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I32cc12cdacef1a4ef64577e0fa977f46     <=
                                             If86871aa91ead2d985e915f4d58408f3[SGN_MAX_SUM_WDTH] ?
                                             ~If86871aa91ead2d985e915f4d58408f3 + 1 :
                                             If86871aa91ead2d985e915f4d58408f3
                                             ;

            I17cf58ef5326978c62c03c56090a299f  <=  If86871aa91ead2d985e915f4d58408f3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I26b3f2360ca4a8caee61b2f3a3a08267     <=
                                             Ie53d1075a122b58f8ee4282b91322ccc[SGN_MAX_SUM_WDTH] ?
                                             ~Ie53d1075a122b58f8ee4282b91322ccc + 1 :
                                             Ie53d1075a122b58f8ee4282b91322ccc
                                             ;

            Ie41ca18c7d11a47e274f9c33f75393ec  <=  Ie53d1075a122b58f8ee4282b91322ccc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ef9b7dc0c63e9ca6a5fb5f7ffa06041     <=
                                             I54acee9cb56584f9876867492fabe469[SGN_MAX_SUM_WDTH] ?
                                             ~I54acee9cb56584f9876867492fabe469 + 1 :
                                             I54acee9cb56584f9876867492fabe469
                                             ;

            I7b80b4902fe98c10dd72c9eb082346e5  <=  I54acee9cb56584f9876867492fabe469[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If881473b05090f40a027d7eeee7f7ed9     <=
                                             Ia4e992a0d0c4f89e3bbaba81b6be3c41[SGN_MAX_SUM_WDTH] ?
                                             ~Ia4e992a0d0c4f89e3bbaba81b6be3c41 + 1 :
                                             Ia4e992a0d0c4f89e3bbaba81b6be3c41
                                             ;

            I20ffba20af04b99954bf719589e90d1a  <=  Ia4e992a0d0c4f89e3bbaba81b6be3c41[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I23bd59ab5b038935301396aaf2acefc1     <=
                                             I8c215a65ea37a535fc9230a0141d209f[SGN_MAX_SUM_WDTH] ?
                                             ~I8c215a65ea37a535fc9230a0141d209f + 1 :
                                             I8c215a65ea37a535fc9230a0141d209f
                                             ;

            If8fe5af7e5c3c97b5a713f6bcf919f1f  <=  I8c215a65ea37a535fc9230a0141d209f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I874386d94dacf84e699d159af1a49836     <=
                                             I564374188b8065f6a46972355d27b0a9[SGN_MAX_SUM_WDTH] ?
                                             ~I564374188b8065f6a46972355d27b0a9 + 1 :
                                             I564374188b8065f6a46972355d27b0a9
                                             ;

            Idc5fb0f3a04ab32948e249e088a11b11  <=  I564374188b8065f6a46972355d27b0a9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95bfe51a759bf4165168e5e3b99d6b34     <=
                                             Ide9ea9ced1a2398876700b19dd25a080[SGN_MAX_SUM_WDTH] ?
                                             ~Ide9ea9ced1a2398876700b19dd25a080 + 1 :
                                             Ide9ea9ced1a2398876700b19dd25a080
                                             ;

            Ia9f1e580e8f441394d719d52a7bad688  <=  Ide9ea9ced1a2398876700b19dd25a080[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4ba5b2f9b7ec0937ecd2c9945cf6de87     <=
                                             I999b0d3276b81801b5a6a5af4d98e6fc[SGN_MAX_SUM_WDTH] ?
                                             ~I999b0d3276b81801b5a6a5af4d98e6fc + 1 :
                                             I999b0d3276b81801b5a6a5af4d98e6fc
                                             ;

            I02849282dd1bd663fd39baccf41762f9  <=  I999b0d3276b81801b5a6a5af4d98e6fc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b08fb8db0e8a1de3d416907c87fe700     <=
                                             I94b6767c45b74142ab2d457b5fe3b64e[SGN_MAX_SUM_WDTH] ?
                                             ~I94b6767c45b74142ab2d457b5fe3b64e + 1 :
                                             I94b6767c45b74142ab2d457b5fe3b64e
                                             ;

            Ie4cda4648f6ceb76b8fb74f290ab6439  <=  I94b6767c45b74142ab2d457b5fe3b64e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie030d12e5acf9ef4975a17c83b2481c1     <=
                                             I2062510b4d8249d8a9b75377d4513266[SGN_MAX_SUM_WDTH] ?
                                             ~I2062510b4d8249d8a9b75377d4513266 + 1 :
                                             I2062510b4d8249d8a9b75377d4513266
                                             ;

            I24135210c23b2422a42c90ee25594191  <=  I2062510b4d8249d8a9b75377d4513266[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia7a0e852d3dfcef950804ea0ebb0c80a     <=
                                             Iba97ce79b40d24270208680c74b41799[SGN_MAX_SUM_WDTH] ?
                                             ~Iba97ce79b40d24270208680c74b41799 + 1 :
                                             Iba97ce79b40d24270208680c74b41799
                                             ;

            Ib08897f9216599042f7b97b137e07fe1  <=  Iba97ce79b40d24270208680c74b41799[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iaa4c38d030eab2b7899399aa0d7886d9     <=
                                             I35b405f29c891a3ccaf0b64443d114e9[SGN_MAX_SUM_WDTH] ?
                                             ~I35b405f29c891a3ccaf0b64443d114e9 + 1 :
                                             I35b405f29c891a3ccaf0b64443d114e9
                                             ;

            I51e14ece9ab6607f83e6ba27f3f046a9  <=  I35b405f29c891a3ccaf0b64443d114e9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icce7ff1d652d4d9c2be5ecf679059bbe     <=
                                             Ib44c2f3a3916b3eaa7452f0126f934ab[SGN_MAX_SUM_WDTH] ?
                                             ~Ib44c2f3a3916b3eaa7452f0126f934ab + 1 :
                                             Ib44c2f3a3916b3eaa7452f0126f934ab
                                             ;

            I7a626ec321bf963a5401892a7e3891c7  <=  Ib44c2f3a3916b3eaa7452f0126f934ab[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If816bc5eacaea23443602e575ddf60b8     <=
                                             I2f0d79178e118fb89f9504e5f75fd612[SGN_MAX_SUM_WDTH] ?
                                             ~I2f0d79178e118fb89f9504e5f75fd612 + 1 :
                                             I2f0d79178e118fb89f9504e5f75fd612
                                             ;

            If76f04fe0baf171d7df2c0cd849aea2b  <=  I2f0d79178e118fb89f9504e5f75fd612[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3b224a4ded05446cc5300d430bdd1947     <=
                                             I1e5f655fd8601930d7c9307aab545391[SGN_MAX_SUM_WDTH] ?
                                             ~I1e5f655fd8601930d7c9307aab545391 + 1 :
                                             I1e5f655fd8601930d7c9307aab545391
                                             ;

            Ia9c8cc5e3becf3d48feedec8fa2c93a4  <=  I1e5f655fd8601930d7c9307aab545391[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia5fc5cfb0e52237b407b37a3858fccb5     <=
                                             I77691bc302dff581968daeeeaf44e9a9[SGN_MAX_SUM_WDTH] ?
                                             ~I77691bc302dff581968daeeeaf44e9a9 + 1 :
                                             I77691bc302dff581968daeeeaf44e9a9
                                             ;

            If3b77c41fabcdb283f2c6fdacaa5e9a4  <=  I77691bc302dff581968daeeeaf44e9a9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I92f8ba6e7f8e9b30fb5b6973eb8fd03e     <=
                                             Ic0f0982cdd813ef3da99d8534e23c9e7[SGN_MAX_SUM_WDTH] ?
                                             ~Ic0f0982cdd813ef3da99d8534e23c9e7 + 1 :
                                             Ic0f0982cdd813ef3da99d8534e23c9e7
                                             ;

            Ie5373b01a92f2ff85be8077cfef2175a  <=  Ic0f0982cdd813ef3da99d8534e23c9e7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icdfa60d2a024dd934f7e6639c6cb2c28     <=
                                             I449f136e29d92eedd2273b58bd34431c[SGN_MAX_SUM_WDTH] ?
                                             ~I449f136e29d92eedd2273b58bd34431c + 1 :
                                             I449f136e29d92eedd2273b58bd34431c
                                             ;

            I5109afc4dc91780e05704ea5e1399e3e  <=  I449f136e29d92eedd2273b58bd34431c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifff70b976513eaa42b6bd4b80c98611e     <=
                                             I0906f557008adaf488966d5aa989e6ae[SGN_MAX_SUM_WDTH] ?
                                             ~I0906f557008adaf488966d5aa989e6ae + 1 :
                                             I0906f557008adaf488966d5aa989e6ae
                                             ;

            I3e0b41bee4c76eb5f3340ad23bfa01ad  <=  I0906f557008adaf488966d5aa989e6ae[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica12fa8b631b70a6bbe9f6e92bf73ea0     <=
                                             Ic0b69b2b6f55b4613bac3aad8e864c9f[SGN_MAX_SUM_WDTH] ?
                                             ~Ic0b69b2b6f55b4613bac3aad8e864c9f + 1 :
                                             Ic0b69b2b6f55b4613bac3aad8e864c9f
                                             ;

            Ic0732810fd355d59a3168be896a0f9ac  <=  Ic0b69b2b6f55b4613bac3aad8e864c9f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie69c255335760f706c644b115887269b     <=
                                             I6ccadd50ca8d59878cf089a35319b6c0[SGN_MAX_SUM_WDTH] ?
                                             ~I6ccadd50ca8d59878cf089a35319b6c0 + 1 :
                                             I6ccadd50ca8d59878cf089a35319b6c0
                                             ;

            I220e32641265b46527ca61111f7ebf1b  <=  I6ccadd50ca8d59878cf089a35319b6c0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idb06676b41de19bc86eae34c292183d9     <=
                                             Ia5aabf0fe6a5d3731b363c80a7238a14[SGN_MAX_SUM_WDTH] ?
                                             ~Ia5aabf0fe6a5d3731b363c80a7238a14 + 1 :
                                             Ia5aabf0fe6a5d3731b363c80a7238a14
                                             ;

            Ice59d2af73d0b0f2ae91a2ef0c2b7f04  <=  Ia5aabf0fe6a5d3731b363c80a7238a14[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib21d2306d5ded3406fac754e69a10d20     <=
                                             I217dc03c6c19195b3c2f478b2b8b0bb8[SGN_MAX_SUM_WDTH] ?
                                             ~I217dc03c6c19195b3c2f478b2b8b0bb8 + 1 :
                                             I217dc03c6c19195b3c2f478b2b8b0bb8
                                             ;

            Ic308610ea8bb62ecb6094192e02dbdba  <=  I217dc03c6c19195b3c2f478b2b8b0bb8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib41d1aa2dcf81879976fb8964cbf6f79     <=
                                             I70c592140d0fd63e2b9b8ab9b619df9a[SGN_MAX_SUM_WDTH] ?
                                             ~I70c592140d0fd63e2b9b8ab9b619df9a + 1 :
                                             I70c592140d0fd63e2b9b8ab9b619df9a
                                             ;

            I33ee415d85e2bcd8f975d34b880f6ea7  <=  I70c592140d0fd63e2b9b8ab9b619df9a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5f8f5e246f008b8d8c75f72828337bab     <=
                                             I4d9ac478c0c0b7191a0ffeb3c6d7c521[SGN_MAX_SUM_WDTH] ?
                                             ~I4d9ac478c0c0b7191a0ffeb3c6d7c521 + 1 :
                                             I4d9ac478c0c0b7191a0ffeb3c6d7c521
                                             ;

            Ie61f299252b8fecfd3e8634b64df5a90  <=  I4d9ac478c0c0b7191a0ffeb3c6d7c521[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id6625e78da0e14d2eeb19cc8ac6520e0     <=
                                             I8bb214c6ec5a16858101699241a1b4bb[SGN_MAX_SUM_WDTH] ?
                                             ~I8bb214c6ec5a16858101699241a1b4bb + 1 :
                                             I8bb214c6ec5a16858101699241a1b4bb
                                             ;

            Icc67656ad2dd3fffae4e5abe02f8fff9  <=  I8bb214c6ec5a16858101699241a1b4bb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6d9ddc6afa559ac35c042df1a9390ce9     <=
                                             Iff81d398838ac6181e09d95903bf57a9[SGN_MAX_SUM_WDTH] ?
                                             ~Iff81d398838ac6181e09d95903bf57a9 + 1 :
                                             Iff81d398838ac6181e09d95903bf57a9
                                             ;

            I0c47ccef4b55410286248884a7249703  <=  Iff81d398838ac6181e09d95903bf57a9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9334055c7833676469670372d3c5cc31     <=
                                             I710eb104c64c7eb72a55cbfc11bff827[SGN_MAX_SUM_WDTH] ?
                                             ~I710eb104c64c7eb72a55cbfc11bff827 + 1 :
                                             I710eb104c64c7eb72a55cbfc11bff827
                                             ;

            I94e4041b482064334fd0ed92b91bde89  <=  I710eb104c64c7eb72a55cbfc11bff827[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0c97d772c737c6ff85b584bf69ccaf93     <=
                                             I9f2d9117540a1d6902b1a7ec3e9d5ab4[SGN_MAX_SUM_WDTH] ?
                                             ~I9f2d9117540a1d6902b1a7ec3e9d5ab4 + 1 :
                                             I9f2d9117540a1d6902b1a7ec3e9d5ab4
                                             ;

            I39d3bce4060032a81e6b6a1c1805cfe8  <=  I9f2d9117540a1d6902b1a7ec3e9d5ab4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic6ce97ae85d91dd8a79f3f9d0da375a2     <=
                                             Ie3204e2e502d2c192994f3c74f1ea38f[SGN_MAX_SUM_WDTH] ?
                                             ~Ie3204e2e502d2c192994f3c74f1ea38f + 1 :
                                             Ie3204e2e502d2c192994f3c74f1ea38f
                                             ;

            Ifb422c30663eb4824caa72326b238df6  <=  Ie3204e2e502d2c192994f3c74f1ea38f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I83ff9a2750b298b0f7c9b6ce13f574af     <=
                                             I97f03a2baec02107032233e68c0b146b[SGN_MAX_SUM_WDTH] ?
                                             ~I97f03a2baec02107032233e68c0b146b + 1 :
                                             I97f03a2baec02107032233e68c0b146b
                                             ;

            I41ab6fb6ec6ef7ffff70e50f25f217b6  <=  I97f03a2baec02107032233e68c0b146b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I85699a2a05c343a6a9e828af6d445e9e     <=
                                             I860ccc9f56a3376ea0e8137a045fe650[SGN_MAX_SUM_WDTH] ?
                                             ~I860ccc9f56a3376ea0e8137a045fe650 + 1 :
                                             I860ccc9f56a3376ea0e8137a045fe650
                                             ;

            I3ce10718a2211184999663c3c2493cc1  <=  I860ccc9f56a3376ea0e8137a045fe650[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I51f6e39b24b2554884e381be79f47ff2     <=
                                             I7b00537ae91be6f2ad8be0776e29da79[SGN_MAX_SUM_WDTH] ?
                                             ~I7b00537ae91be6f2ad8be0776e29da79 + 1 :
                                             I7b00537ae91be6f2ad8be0776e29da79
                                             ;

            I877e8d94236c3d8b0a31858a98fba5d6  <=  I7b00537ae91be6f2ad8be0776e29da79[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9f65fd05c6929300860c8cbbde5607f2     <=
                                             I68413adceb35fe859824c32bb76d9906[SGN_MAX_SUM_WDTH] ?
                                             ~I68413adceb35fe859824c32bb76d9906 + 1 :
                                             I68413adceb35fe859824c32bb76d9906
                                             ;

            Iff2f1716cbd73b406d8f07c22dc79fc8  <=  I68413adceb35fe859824c32bb76d9906[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If09761d8f06051d4287ee29ac9c9fa19     <=
                                             Ib61183063f591e5845ca8ce70f598c79[SGN_MAX_SUM_WDTH] ?
                                             ~Ib61183063f591e5845ca8ce70f598c79 + 1 :
                                             Ib61183063f591e5845ca8ce70f598c79
                                             ;

            Ibc48fabc172f27ebce18d0a9b5120dc5  <=  Ib61183063f591e5845ca8ce70f598c79[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I33bfbe0bcca6d32c86b9576577e3f265     <=
                                             Ia7a97e75655c4eaa8652f43c27d5ae50[SGN_MAX_SUM_WDTH] ?
                                             ~Ia7a97e75655c4eaa8652f43c27d5ae50 + 1 :
                                             Ia7a97e75655c4eaa8652f43c27d5ae50
                                             ;

            Ie562ebb336e476a81f20a652d4cb20f1  <=  Ia7a97e75655c4eaa8652f43c27d5ae50[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If2921210b1c05ecbf00af3a2bcb96ef4     <=
                                             I0402af748fe9d48a514d23691a2cb6b8[SGN_MAX_SUM_WDTH] ?
                                             ~I0402af748fe9d48a514d23691a2cb6b8 + 1 :
                                             I0402af748fe9d48a514d23691a2cb6b8
                                             ;

            Ib5ee5a6ffc45ed1fece0822dc4619b57  <=  I0402af748fe9d48a514d23691a2cb6b8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib074e38e280474a782da831a3e0028b4     <=
                                             I5e9d62da7f6aeaa717f5a394e2531210[SGN_MAX_SUM_WDTH] ?
                                             ~I5e9d62da7f6aeaa717f5a394e2531210 + 1 :
                                             I5e9d62da7f6aeaa717f5a394e2531210
                                             ;

            I86ba73ee348f80e2f9891d2ebc8a02ed  <=  I5e9d62da7f6aeaa717f5a394e2531210[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I507449dde0bc0c8f53a10759436ec731     <=
                                             Idb3666a01522d57729513cd3f18c9798[SGN_MAX_SUM_WDTH] ?
                                             ~Idb3666a01522d57729513cd3f18c9798 + 1 :
                                             Idb3666a01522d57729513cd3f18c9798
                                             ;

            I1e96d5af3d0e3fdce39530dfd0131a7d  <=  Idb3666a01522d57729513cd3f18c9798[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id55a3e3f2d75baeba71a345fad695c69     <=
                                             Ifb6e917336ab665d9bfea6dcfe21bc8c[SGN_MAX_SUM_WDTH] ?
                                             ~Ifb6e917336ab665d9bfea6dcfe21bc8c + 1 :
                                             Ifb6e917336ab665d9bfea6dcfe21bc8c
                                             ;

            I38352b363fa37f6f822fbc1a39100968  <=  Ifb6e917336ab665d9bfea6dcfe21bc8c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I20984f43d22671639a7a178ad15aec04     <=
                                             I0adf84fd4ea2e882b59a42dad6683707[SGN_MAX_SUM_WDTH] ?
                                             ~I0adf84fd4ea2e882b59a42dad6683707 + 1 :
                                             I0adf84fd4ea2e882b59a42dad6683707
                                             ;

            I4ba41864bb1d2130c6971e0b2903027a  <=  I0adf84fd4ea2e882b59a42dad6683707[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I59f88336d6bdd50ded87d353fb5ce3e9     <=
                                             I1d0e0cb3903cece98c3a65f920e5ab21[SGN_MAX_SUM_WDTH] ?
                                             ~I1d0e0cb3903cece98c3a65f920e5ab21 + 1 :
                                             I1d0e0cb3903cece98c3a65f920e5ab21
                                             ;

            Ib68deeb7bec4ca3585d1a4dcbf8793f1  <=  I1d0e0cb3903cece98c3a65f920e5ab21[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I488635e3f7ed77ea88199f5bffd4b1d6     <=
                                             I8b12d3b1f65fad05577cf25e8d7950a5[SGN_MAX_SUM_WDTH] ?
                                             ~I8b12d3b1f65fad05577cf25e8d7950a5 + 1 :
                                             I8b12d3b1f65fad05577cf25e8d7950a5
                                             ;

            Ida3d808d100e0bba290f96ed9e744e65  <=  I8b12d3b1f65fad05577cf25e8d7950a5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie6893017d21c050ba10d206854f4a9f4     <=
                                             Ifb24658924186dba2d1a85ee28fc0313[SGN_MAX_SUM_WDTH] ?
                                             ~Ifb24658924186dba2d1a85ee28fc0313 + 1 :
                                             Ifb24658924186dba2d1a85ee28fc0313
                                             ;

            I4d4901ff372f6820ca9c8c29cefa664a  <=  Ifb24658924186dba2d1a85ee28fc0313[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id3f68b4dc0ab60673208b7d2081f3533     <=
                                             I067250d29597d7c71da50f8cf557eb61[SGN_MAX_SUM_WDTH] ?
                                             ~I067250d29597d7c71da50f8cf557eb61 + 1 :
                                             I067250d29597d7c71da50f8cf557eb61
                                             ;

            Ib99e1b93fb7fbda260d93eea3d24c3e9  <=  I067250d29597d7c71da50f8cf557eb61[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I433756b944e061a824a89bda241e879f     <=
                                             Ic86c9a00eacc20772706da9399aab4ba[SGN_MAX_SUM_WDTH] ?
                                             ~Ic86c9a00eacc20772706da9399aab4ba + 1 :
                                             Ic86c9a00eacc20772706da9399aab4ba
                                             ;

            I019e399a1cef87745e025a7d74e94db0  <=  Ic86c9a00eacc20772706da9399aab4ba[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2eb60a922aa4f7482dd92b9351d53a2d     <=
                                             I8271913876a2729269e844dc4809a25f[SGN_MAX_SUM_WDTH] ?
                                             ~I8271913876a2729269e844dc4809a25f + 1 :
                                             I8271913876a2729269e844dc4809a25f
                                             ;

            Ia8974083bfd064f2c27dcd421490fcfd  <=  I8271913876a2729269e844dc4809a25f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0867979e1b159c8ceae548930376f482     <=
                                             I3af8e500702e46e7330796cb23979266[SGN_MAX_SUM_WDTH] ?
                                             ~I3af8e500702e46e7330796cb23979266 + 1 :
                                             I3af8e500702e46e7330796cb23979266
                                             ;

            I8fd5787ebf758919e7cb75d7419441e8  <=  I3af8e500702e46e7330796cb23979266[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4accfbeae8a5ee0dbeab23ef3a116145     <=
                                             Ice852e353c55faedcde1922d0179b30a[SGN_MAX_SUM_WDTH] ?
                                             ~Ice852e353c55faedcde1922d0179b30a + 1 :
                                             Ice852e353c55faedcde1922d0179b30a
                                             ;

            Id14074d5230885c38b89b09b130ecf68  <=  Ice852e353c55faedcde1922d0179b30a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic7570b0b7c5bef5758f68562ae4c90f6     <=
                                             Ibb9864cd5bcd1ef1fc7bfd822db3150b[SGN_MAX_SUM_WDTH] ?
                                             ~Ibb9864cd5bcd1ef1fc7bfd822db3150b + 1 :
                                             Ibb9864cd5bcd1ef1fc7bfd822db3150b
                                             ;

            I86fefad34d3c864dd0e725133f303b4f  <=  Ibb9864cd5bcd1ef1fc7bfd822db3150b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iceadadc4456881fdeea85934a9bf4d6c     <=
                                             I13f58835ab9e6362ffddf06976c97207[SGN_MAX_SUM_WDTH] ?
                                             ~I13f58835ab9e6362ffddf06976c97207 + 1 :
                                             I13f58835ab9e6362ffddf06976c97207
                                             ;

            I1ca188bcdebbf41d84f7a5220bd1d195  <=  I13f58835ab9e6362ffddf06976c97207[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7b2b617ae67424f54961eebce42de77e     <=
                                             I35bfac2d8d88c61e93a27db564f9ecef[SGN_MAX_SUM_WDTH] ?
                                             ~I35bfac2d8d88c61e93a27db564f9ecef + 1 :
                                             I35bfac2d8d88c61e93a27db564f9ecef
                                             ;

            Ifc640243288c9b37b7eb9e00351b23f0  <=  I35bfac2d8d88c61e93a27db564f9ecef[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I953f0f8af76f89b2d9ab4abf19fb411d     <=
                                             I7ecdf9f7726df27510f35fe6c1b5b4be[SGN_MAX_SUM_WDTH] ?
                                             ~I7ecdf9f7726df27510f35fe6c1b5b4be + 1 :
                                             I7ecdf9f7726df27510f35fe6c1b5b4be
                                             ;

            I3d149293f106ae8680c7f4702daa0bd6  <=  I7ecdf9f7726df27510f35fe6c1b5b4be[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I915b4736dcb20f831d02e48f4e79f008     <=
                                             I7327385650ea109a8bb07f1c92252d28[SGN_MAX_SUM_WDTH] ?
                                             ~I7327385650ea109a8bb07f1c92252d28 + 1 :
                                             I7327385650ea109a8bb07f1c92252d28
                                             ;

            Ie232799bd6c4ec99e24c78f3ad798265  <=  I7327385650ea109a8bb07f1c92252d28[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7eec587348ae1ca1f00c0a3ad10ad27     <=
                                             Ib5d66de65bb7bc9e1f7b3f05e4bd703b[SGN_MAX_SUM_WDTH] ?
                                             ~Ib5d66de65bb7bc9e1f7b3f05e4bd703b + 1 :
                                             Ib5d66de65bb7bc9e1f7b3f05e4bd703b
                                             ;

            Ifebcf64858d5e2d07ad7894d6182eb11  <=  Ib5d66de65bb7bc9e1f7b3f05e4bd703b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I001a212686304248c8359e5fc01227c0     <=
                                             Ifca73a480a501ea2636c47e487987167[SGN_MAX_SUM_WDTH] ?
                                             ~Ifca73a480a501ea2636c47e487987167 + 1 :
                                             Ifca73a480a501ea2636c47e487987167
                                             ;

            Ibab55499323660588ec82ebd07ab0572  <=  Ifca73a480a501ea2636c47e487987167[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibb7554e012c0fc1223c29b759c900666     <=
                                             I75a3f16cb4ddc4b0478fb1c07c10aba8[SGN_MAX_SUM_WDTH] ?
                                             ~I75a3f16cb4ddc4b0478fb1c07c10aba8 + 1 :
                                             I75a3f16cb4ddc4b0478fb1c07c10aba8
                                             ;

            I89af7644c48a80d7d22f50b008d35841  <=  I75a3f16cb4ddc4b0478fb1c07c10aba8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9aeb9c42b54a05be6bf9b7b88b6860ba     <=
                                             I5603979fb76ebb2bab9a8764c4833b52[SGN_MAX_SUM_WDTH] ?
                                             ~I5603979fb76ebb2bab9a8764c4833b52 + 1 :
                                             I5603979fb76ebb2bab9a8764c4833b52
                                             ;

            I0152dc6e6a7acd72a2144623e63998ef  <=  I5603979fb76ebb2bab9a8764c4833b52[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6a5a5966965b0790b906c6fda71aef80     <=
                                             I939430bcba9f8bb28f5782040a4c76e7[SGN_MAX_SUM_WDTH] ?
                                             ~I939430bcba9f8bb28f5782040a4c76e7 + 1 :
                                             I939430bcba9f8bb28f5782040a4c76e7
                                             ;

            I951dedd7af44c3865a8f36888432d0c9  <=  I939430bcba9f8bb28f5782040a4c76e7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic943083ca65ace6c42d73f4234739a06     <=
                                             I71ed74fcff44b1a6ec1ddf7b18cf8a31[SGN_MAX_SUM_WDTH] ?
                                             ~I71ed74fcff44b1a6ec1ddf7b18cf8a31 + 1 :
                                             I71ed74fcff44b1a6ec1ddf7b18cf8a31
                                             ;

            I8188dd7cb03854c6f709de06ff785d91  <=  I71ed74fcff44b1a6ec1ddf7b18cf8a31[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id0b321686d4c39621024cf0dd99822dc     <=
                                             Icc204071ef0dd850f42840be901a1c8c[SGN_MAX_SUM_WDTH] ?
                                             ~Icc204071ef0dd850f42840be901a1c8c + 1 :
                                             Icc204071ef0dd850f42840be901a1c8c
                                             ;

            I3b30b4ab00a49e10a75587aa324d6132  <=  Icc204071ef0dd850f42840be901a1c8c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0839dd3787442f1b79b87e02436bfdce     <=
                                             Ie8187be889aa7f205231e2e60cb827e3[SGN_MAX_SUM_WDTH] ?
                                             ~Ie8187be889aa7f205231e2e60cb827e3 + 1 :
                                             Ie8187be889aa7f205231e2e60cb827e3
                                             ;

            Ie50aca688b3433fad7565998cb900155  <=  Ie8187be889aa7f205231e2e60cb827e3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I89e6a9fd97d8aa4dd3b832c3be4697b2     <=
                                             I18c57ba0c68acdec8308c2ba40482668[SGN_MAX_SUM_WDTH] ?
                                             ~I18c57ba0c68acdec8308c2ba40482668 + 1 :
                                             I18c57ba0c68acdec8308c2ba40482668
                                             ;

            I3342fe0c5d3ee5021892d53eb45bde21  <=  I18c57ba0c68acdec8308c2ba40482668[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I93d4157f48b132642752220059861e98     <=
                                             If45f0a6203e1a6ef6e0d86ccccab3920[SGN_MAX_SUM_WDTH] ?
                                             ~If45f0a6203e1a6ef6e0d86ccccab3920 + 1 :
                                             If45f0a6203e1a6ef6e0d86ccccab3920
                                             ;

            I5134b762ac428bed07ce102d8927a418  <=  If45f0a6203e1a6ef6e0d86ccccab3920[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8fc4faa2891d7fd3479ac1f788f481dc     <=
                                             I834626bbcdd99143f36052aa6e77de49[SGN_MAX_SUM_WDTH] ?
                                             ~I834626bbcdd99143f36052aa6e77de49 + 1 :
                                             I834626bbcdd99143f36052aa6e77de49
                                             ;

            Ic14f948884da19a272a4760ffaab9ea9  <=  I834626bbcdd99143f36052aa6e77de49[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I440f30e9cb4bc89233b46ea00b4cbeb4     <=
                                             I58860aa281debf67db1369b2e22b9f5b[SGN_MAX_SUM_WDTH] ?
                                             ~I58860aa281debf67db1369b2e22b9f5b + 1 :
                                             I58860aa281debf67db1369b2e22b9f5b
                                             ;

            I46e1047bca2b38e62b4de80d1d2249de  <=  I58860aa281debf67db1369b2e22b9f5b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6568bfd8780c11e0b1b049a01f92abd8     <=
                                             I885d19716778193c3288c8322cfd32ae[SGN_MAX_SUM_WDTH] ?
                                             ~I885d19716778193c3288c8322cfd32ae + 1 :
                                             I885d19716778193c3288c8322cfd32ae
                                             ;

            I866b30a63b3b5fb708934a1cbb0e1d9a  <=  I885d19716778193c3288c8322cfd32ae[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibf7dc4da07f9955d5d4c7e1f63f1ad68     <=
                                             I19a6d51c460b600130966b5be281d23e[SGN_MAX_SUM_WDTH] ?
                                             ~I19a6d51c460b600130966b5be281d23e + 1 :
                                             I19a6d51c460b600130966b5be281d23e
                                             ;

            Iaddc1f2e822fd2fe9d9046d759a82cb4  <=  I19a6d51c460b600130966b5be281d23e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7ec1a328587b72a39c462083efea0ee0     <=
                                             I7a4326b2355162700b8647861c80f43f[SGN_MAX_SUM_WDTH] ?
                                             ~I7a4326b2355162700b8647861c80f43f + 1 :
                                             I7a4326b2355162700b8647861c80f43f
                                             ;

            If9285bf7611bcc5ea6432215c349e021  <=  I7a4326b2355162700b8647861c80f43f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iaf028e7ab4dc77a7649f15d603834b5f     <=
                                             I40ce63d36b1aa901d29c0ecc3ad20a66[SGN_MAX_SUM_WDTH] ?
                                             ~I40ce63d36b1aa901d29c0ecc3ad20a66 + 1 :
                                             I40ce63d36b1aa901d29c0ecc3ad20a66
                                             ;

            Id277f5f05551eeb5dec1701056330da1  <=  I40ce63d36b1aa901d29c0ecc3ad20a66[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I58db79a8e9f0cd1ded379897ba2f27ae     <=
                                             I32230b8893dd9fd1da4ce1f2553b5550[SGN_MAX_SUM_WDTH] ?
                                             ~I32230b8893dd9fd1da4ce1f2553b5550 + 1 :
                                             I32230b8893dd9fd1da4ce1f2553b5550
                                             ;

            I9963d0b24763ed8038b1f3922b8f9548  <=  I32230b8893dd9fd1da4ce1f2553b5550[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6d3cb4ccb4e51c7e6603d0abd1a082c4     <=
                                             If7fb4fa70b6803a7e4c64a834669dbfa[SGN_MAX_SUM_WDTH] ?
                                             ~If7fb4fa70b6803a7e4c64a834669dbfa + 1 :
                                             If7fb4fa70b6803a7e4c64a834669dbfa
                                             ;

            Ia98de3691917dfb63bebdc3f8655c8be  <=  If7fb4fa70b6803a7e4c64a834669dbfa[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I79f75f49ea8a29d684af396014b2f3ab     <=
                                             Iaf1e5c8b7267eca64468227734dcfbdb[SGN_MAX_SUM_WDTH] ?
                                             ~Iaf1e5c8b7267eca64468227734dcfbdb + 1 :
                                             Iaf1e5c8b7267eca64468227734dcfbdb
                                             ;

            I0bce960fcc58938e6a1e01b912eabbf2  <=  Iaf1e5c8b7267eca64468227734dcfbdb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9c5ecd86bedb189fada40fae9d751a68     <=
                                             I5ab38b4a054c50fced80e9323f4a9ddf[SGN_MAX_SUM_WDTH] ?
                                             ~I5ab38b4a054c50fced80e9323f4a9ddf + 1 :
                                             I5ab38b4a054c50fced80e9323f4a9ddf
                                             ;

            Ice5f7168aeb940d48093cc9df7cba36b  <=  I5ab38b4a054c50fced80e9323f4a9ddf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iad5f06e1989ead7d306c70a3b02cb8f4     <=
                                             I779f57a085e170d2ab7e7b5f046e42e6[SGN_MAX_SUM_WDTH] ?
                                             ~I779f57a085e170d2ab7e7b5f046e42e6 + 1 :
                                             I779f57a085e170d2ab7e7b5f046e42e6
                                             ;

            I859d795a7d141eb777c1f3c038203794  <=  I779f57a085e170d2ab7e7b5f046e42e6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If6d1a410df5a4aea6a01337a6074fbd9     <=
                                             I120e630331e23d75054584a44aafaf63[SGN_MAX_SUM_WDTH] ?
                                             ~I120e630331e23d75054584a44aafaf63 + 1 :
                                             I120e630331e23d75054584a44aafaf63
                                             ;

            I0dccb8eaad52ce4d780696a8485420f1  <=  I120e630331e23d75054584a44aafaf63[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3bc40a4db14566b5099b14cee5f61135     <=
                                             I3f690a6c75649328d7cccf08cc6ca81b[SGN_MAX_SUM_WDTH] ?
                                             ~I3f690a6c75649328d7cccf08cc6ca81b + 1 :
                                             I3f690a6c75649328d7cccf08cc6ca81b
                                             ;

            I6d4fc81ced37c159303c243af04d345e  <=  I3f690a6c75649328d7cccf08cc6ca81b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7e683fd8235d7cfbf4ff407a286f07de     <=
                                             I2105fce588dc6840254a1eaf02b549c9[SGN_MAX_SUM_WDTH] ?
                                             ~I2105fce588dc6840254a1eaf02b549c9 + 1 :
                                             I2105fce588dc6840254a1eaf02b549c9
                                             ;

            Iefdb8bd28839af9413a3906cbfe715e6  <=  I2105fce588dc6840254a1eaf02b549c9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I97afcedf05e588b7976d6005191dc916     <=
                                             Ic0b28cd43f561513b63ff20e31038f37[SGN_MAX_SUM_WDTH] ?
                                             ~Ic0b28cd43f561513b63ff20e31038f37 + 1 :
                                             Ic0b28cd43f561513b63ff20e31038f37
                                             ;

            I0615acb0f7cf79b5f6ae8e91cb525dc9  <=  Ic0b28cd43f561513b63ff20e31038f37[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib8d8eec0aaa662adf2837c9b705fce7e     <=
                                             Ib4e0926a64eaefff0e36fdde4783e923[SGN_MAX_SUM_WDTH] ?
                                             ~Ib4e0926a64eaefff0e36fdde4783e923 + 1 :
                                             Ib4e0926a64eaefff0e36fdde4783e923
                                             ;

            Ieed4c810a5bb69de112522dcf00b16ed  <=  Ib4e0926a64eaefff0e36fdde4783e923[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icbd765be950123705955e2c5d7ace84b     <=
                                             Ieb485d7a868decbc901fad618f56412a[SGN_MAX_SUM_WDTH] ?
                                             ~Ieb485d7a868decbc901fad618f56412a + 1 :
                                             Ieb485d7a868decbc901fad618f56412a
                                             ;

            If533578cacb685a95afbb8e1c05d3c07  <=  Ieb485d7a868decbc901fad618f56412a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I706e8f5617cfae1e6fc83db18c8b5fe3     <=
                                             I71853033c5b7e4e98414209075b4d708[SGN_MAX_SUM_WDTH] ?
                                             ~I71853033c5b7e4e98414209075b4d708 + 1 :
                                             I71853033c5b7e4e98414209075b4d708
                                             ;

            Ia858ff5551286beffd4cf82f876d30ac  <=  I71853033c5b7e4e98414209075b4d708[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1dd8f8c7f1b673898096b1f3ae383197     <=
                                             I37621b4bc9c88a42a47d3123465fa4d5[SGN_MAX_SUM_WDTH] ?
                                             ~I37621b4bc9c88a42a47d3123465fa4d5 + 1 :
                                             I37621b4bc9c88a42a47d3123465fa4d5
                                             ;

            I4c66570630a650fa7b9bec543f685487  <=  I37621b4bc9c88a42a47d3123465fa4d5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I10ca8978cf4659265ed25a27d09acc1c     <=
                                             Ied0d483617ee30ac0539009fba84a684[SGN_MAX_SUM_WDTH] ?
                                             ~Ied0d483617ee30ac0539009fba84a684 + 1 :
                                             Ied0d483617ee30ac0539009fba84a684
                                             ;

            If10f33385e236eaba56cbab8c2883399  <=  Ied0d483617ee30ac0539009fba84a684[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iec4656b32460def4a608b6b0f6486af9     <=
                                             I574d31b300f16225a707bbae0918c445[SGN_MAX_SUM_WDTH] ?
                                             ~I574d31b300f16225a707bbae0918c445 + 1 :
                                             I574d31b300f16225a707bbae0918c445
                                             ;

            I7cb58e4c486e683faa4acad4756815d5  <=  I574d31b300f16225a707bbae0918c445[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5f4475897d1d58965da1b35fe0ef8c01     <=
                                             I9fef812393d8a5f87abc46add3371777[SGN_MAX_SUM_WDTH] ?
                                             ~I9fef812393d8a5f87abc46add3371777 + 1 :
                                             I9fef812393d8a5f87abc46add3371777
                                             ;

            I452e51cca9acec44e36e4efd21b43034  <=  I9fef812393d8a5f87abc46add3371777[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ife61469306df3cf220666b187f1496a9     <=
                                             I64a11eacbd9a28d7e65c56c38127876b[SGN_MAX_SUM_WDTH] ?
                                             ~I64a11eacbd9a28d7e65c56c38127876b + 1 :
                                             I64a11eacbd9a28d7e65c56c38127876b
                                             ;

            Ice0234f25de4ab1f03a3cb01a2d61dbf  <=  I64a11eacbd9a28d7e65c56c38127876b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib49319b9dfa4914f92f423ceaf840014     <=
                                             Id11f93a74e2de2ea1e27e9d2858a472f[SGN_MAX_SUM_WDTH] ?
                                             ~Id11f93a74e2de2ea1e27e9d2858a472f + 1 :
                                             Id11f93a74e2de2ea1e27e9d2858a472f
                                             ;

            I12a18a1f8d4416e9bc8abee6ac3dacfc  <=  Id11f93a74e2de2ea1e27e9d2858a472f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I93ff2f879233cac9b9f0dd2f4c082c09     <=
                                             Ibd0708af1cccb49fded84694d6ffd6f7[SGN_MAX_SUM_WDTH] ?
                                             ~Ibd0708af1cccb49fded84694d6ffd6f7 + 1 :
                                             Ibd0708af1cccb49fded84694d6ffd6f7
                                             ;

            Id17ada8dae3f9810d1892d34f2288859  <=  Ibd0708af1cccb49fded84694d6ffd6f7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I44597d694e9c5d29280e503d72a27c8d     <=
                                             I18edce191243df3a622232f681b7e3f9[SGN_MAX_SUM_WDTH] ?
                                             ~I18edce191243df3a622232f681b7e3f9 + 1 :
                                             I18edce191243df3a622232f681b7e3f9
                                             ;

            Ia2c5fe53cb5b318fa63d09881609655f  <=  I18edce191243df3a622232f681b7e3f9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I04a19448c5e75af8021ad02d1a708bb0     <=
                                             Ib68ae994fc94acf008e424d8f8c8eb4b[SGN_MAX_SUM_WDTH] ?
                                             ~Ib68ae994fc94acf008e424d8f8c8eb4b + 1 :
                                             Ib68ae994fc94acf008e424d8f8c8eb4b
                                             ;

            I579c7926e7b78f4ffc606adc10522f53  <=  Ib68ae994fc94acf008e424d8f8c8eb4b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I71a3093121c2f19dcd1412b468652fa8     <=
                                             Icb6bc0221ed78051fa10967f5cce4a7f[SGN_MAX_SUM_WDTH] ?
                                             ~Icb6bc0221ed78051fa10967f5cce4a7f + 1 :
                                             Icb6bc0221ed78051fa10967f5cce4a7f
                                             ;

            Iffa06a336949f56f4e5a88a06d8b7e60  <=  Icb6bc0221ed78051fa10967f5cce4a7f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3ae09c82029c617034fe6aacbe9e94e6     <=
                                             I3abb9a64f85be533ac16eafaf85c5ad1[SGN_MAX_SUM_WDTH] ?
                                             ~I3abb9a64f85be533ac16eafaf85c5ad1 + 1 :
                                             I3abb9a64f85be533ac16eafaf85c5ad1
                                             ;

            Iaf82668eb49248709540f2f529f1b3e4  <=  I3abb9a64f85be533ac16eafaf85c5ad1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie7af6b3b441f910b000a333afad6c76f     <=
                                             If6badde34faca49e04b3dde9b11c0556[SGN_MAX_SUM_WDTH] ?
                                             ~If6badde34faca49e04b3dde9b11c0556 + 1 :
                                             If6badde34faca49e04b3dde9b11c0556
                                             ;

            I90b3708abdf742370f06cc513ee307e1  <=  If6badde34faca49e04b3dde9b11c0556[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4d71dfea8407aa5b5cbb991bc4fea963     <=
                                             I09d6aa4053f5e1280d70556ad1cc89a4[SGN_MAX_SUM_WDTH] ?
                                             ~I09d6aa4053f5e1280d70556ad1cc89a4 + 1 :
                                             I09d6aa4053f5e1280d70556ad1cc89a4
                                             ;

            Ia17906696bd0e095d7a5297da2e049ea  <=  I09d6aa4053f5e1280d70556ad1cc89a4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1a082caecc831a90e74674ba35da4183     <=
                                             I9d1f949ca74fcf76431906a3a95d4866[SGN_MAX_SUM_WDTH] ?
                                             ~I9d1f949ca74fcf76431906a3a95d4866 + 1 :
                                             I9d1f949ca74fcf76431906a3a95d4866
                                             ;

            I180d4f3b23b518271d7cb8189fbeadc5  <=  I9d1f949ca74fcf76431906a3a95d4866[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iec1de44616a2354a56ab1f681059d4c5     <=
                                             I10221054a7689d49c97a1e908e2fb44b[SGN_MAX_SUM_WDTH] ?
                                             ~I10221054a7689d49c97a1e908e2fb44b + 1 :
                                             I10221054a7689d49c97a1e908e2fb44b
                                             ;

            Id79636d195efff260c430978f0bcee9c  <=  I10221054a7689d49c97a1e908e2fb44b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie3c2318e64d0e218c3db557404c4aac8     <=
                                             I4ec67f577ac5c95d8a93f21935a4fb7f[SGN_MAX_SUM_WDTH] ?
                                             ~I4ec67f577ac5c95d8a93f21935a4fb7f + 1 :
                                             I4ec67f577ac5c95d8a93f21935a4fb7f
                                             ;

            Idbf4ad11ab2a27044193448c8739fec6  <=  I4ec67f577ac5c95d8a93f21935a4fb7f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9a251d50f41e51b1a5cc2475f267e8a0     <=
                                             I069f6a3e5c61b47031648ed6e7ab0330[SGN_MAX_SUM_WDTH] ?
                                             ~I069f6a3e5c61b47031648ed6e7ab0330 + 1 :
                                             I069f6a3e5c61b47031648ed6e7ab0330
                                             ;

            I3051f561a5e1131ebf167cb6ccb5adf4  <=  I069f6a3e5c61b47031648ed6e7ab0330[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9b5767a49f7b9dcb8fdaea924835033c     <=
                                             I4b15910b07c427bfb666057cf4700947[SGN_MAX_SUM_WDTH] ?
                                             ~I4b15910b07c427bfb666057cf4700947 + 1 :
                                             I4b15910b07c427bfb666057cf4700947
                                             ;

            I9322a2a61900943075bbc23c72a3f65d  <=  I4b15910b07c427bfb666057cf4700947[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ca1e6700a19d03621a193c7240bff54     <=
                                             I5694aa90f55816a9ca217470b70f29a6[SGN_MAX_SUM_WDTH] ?
                                             ~I5694aa90f55816a9ca217470b70f29a6 + 1 :
                                             I5694aa90f55816a9ca217470b70f29a6
                                             ;

            Iedc463e359dd3003d9f7e50f3e858e93  <=  I5694aa90f55816a9ca217470b70f29a6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I931c597ff12bffce581f653346202f83     <=
                                             Ia1d3638756959bfb67f32a37c58fe190[SGN_MAX_SUM_WDTH] ?
                                             ~Ia1d3638756959bfb67f32a37c58fe190 + 1 :
                                             Ia1d3638756959bfb67f32a37c58fe190
                                             ;

            Ie7cfdd25541414ff3f8d6e5d7677fbe5  <=  Ia1d3638756959bfb67f32a37c58fe190[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia3a2c5d59f6340917ca3933c05ba4678     <=
                                             I3e81666362b0209c98c5337a74dcbfa9[SGN_MAX_SUM_WDTH] ?
                                             ~I3e81666362b0209c98c5337a74dcbfa9 + 1 :
                                             I3e81666362b0209c98c5337a74dcbfa9
                                             ;

            I1e93f0470d2818249f1c28ef2a399a0e  <=  I3e81666362b0209c98c5337a74dcbfa9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie83d0a8ee5ed214bc7577467748aaa04     <=
                                             Iaa723368e8f531ae9bf99c9b99fdf0f7[SGN_MAX_SUM_WDTH] ?
                                             ~Iaa723368e8f531ae9bf99c9b99fdf0f7 + 1 :
                                             Iaa723368e8f531ae9bf99c9b99fdf0f7
                                             ;

            I5d6e576b0fa7e3219aaf9ccc345085b8  <=  Iaa723368e8f531ae9bf99c9b99fdf0f7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iaac29552e5fc65aaf4f0116f917b707c     <=
                                             I3713f644fba6dd9d4bb4dc3b4c91fe77[SGN_MAX_SUM_WDTH] ?
                                             ~I3713f644fba6dd9d4bb4dc3b4c91fe77 + 1 :
                                             I3713f644fba6dd9d4bb4dc3b4c91fe77
                                             ;

            Id962beade26396738ba0e97f67d5e261  <=  I3713f644fba6dd9d4bb4dc3b4c91fe77[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie2c8eac7204b98139c03b6fbfff9af36     <=
                                             I5a3e3131db6fdd74e5c822fde6a8f2c1[SGN_MAX_SUM_WDTH] ?
                                             ~I5a3e3131db6fdd74e5c822fde6a8f2c1 + 1 :
                                             I5a3e3131db6fdd74e5c822fde6a8f2c1
                                             ;

            Id0ab747d92288f23cef793567b2363d1  <=  I5a3e3131db6fdd74e5c822fde6a8f2c1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ied7fcdaec662cb3c2f89f131986fa102     <=
                                             If18033df3d6ee029fdecf3323ad8d62d[SGN_MAX_SUM_WDTH] ?
                                             ~If18033df3d6ee029fdecf3323ad8d62d + 1 :
                                             If18033df3d6ee029fdecf3323ad8d62d
                                             ;

            Ie536879e6fa9be65376d7f00e0fc40d0  <=  If18033df3d6ee029fdecf3323ad8d62d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib16a17d6430570b45a304d847ee2b11c     <=
                                             I7514cd65da98bd214b4e1da34ac358f1[SGN_MAX_SUM_WDTH] ?
                                             ~I7514cd65da98bd214b4e1da34ac358f1 + 1 :
                                             I7514cd65da98bd214b4e1da34ac358f1
                                             ;

            Ibf312ae4f51fbc44b43848f9df62a45f  <=  I7514cd65da98bd214b4e1da34ac358f1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I42169e454756fe4d1c5f17f2eeb2e091     <=
                                             Id947f3ca55c826ef94d1ac4ad2a227bf[SGN_MAX_SUM_WDTH] ?
                                             ~Id947f3ca55c826ef94d1ac4ad2a227bf + 1 :
                                             Id947f3ca55c826ef94d1ac4ad2a227bf
                                             ;

            Icfc03646b36b971b9fa57d04a26dbfc4  <=  Id947f3ca55c826ef94d1ac4ad2a227bf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6fde38a3a92e06fa77123e3279813c41     <=
                                             Ia6f83033bc647143bbf5377056c7072f[SGN_MAX_SUM_WDTH] ?
                                             ~Ia6f83033bc647143bbf5377056c7072f + 1 :
                                             Ia6f83033bc647143bbf5377056c7072f
                                             ;

            I4f134c0669b5a6a8c7e03be7eee30c6c  <=  Ia6f83033bc647143bbf5377056c7072f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id8ee16437e8d6d6da6d37440e04097b6     <=
                                             I21dd15d84c5abe8d2ac53f65236f587c[SGN_MAX_SUM_WDTH] ?
                                             ~I21dd15d84c5abe8d2ac53f65236f587c + 1 :
                                             I21dd15d84c5abe8d2ac53f65236f587c
                                             ;

            I6c765e677f42fe600b848698c8a78349  <=  I21dd15d84c5abe8d2ac53f65236f587c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibf249d8e5acced9b064132575f40e001     <=
                                             Ia88c70253514b080daa27d2df0aef202[SGN_MAX_SUM_WDTH] ?
                                             ~Ia88c70253514b080daa27d2df0aef202 + 1 :
                                             Ia88c70253514b080daa27d2df0aef202
                                             ;

            I284b23051c85300c2a1e3afe8f25e99e  <=  Ia88c70253514b080daa27d2df0aef202[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I580659084e3d17b48de6b1c66154fcf5     <=
                                             I3cd11d85b17ce4c2181dfd2430ff4595[SGN_MAX_SUM_WDTH] ?
                                             ~I3cd11d85b17ce4c2181dfd2430ff4595 + 1 :
                                             I3cd11d85b17ce4c2181dfd2430ff4595
                                             ;

            I9b560d9baf8a7422b0dd84720e924ced  <=  I3cd11d85b17ce4c2181dfd2430ff4595[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7a14e45d43ab77b265501902152c8616     <=
                                             I9817361d029cc98d7407cf3b8b020567[SGN_MAX_SUM_WDTH] ?
                                             ~I9817361d029cc98d7407cf3b8b020567 + 1 :
                                             I9817361d029cc98d7407cf3b8b020567
                                             ;

            I457ae11ad90c8478751eb4b42764e158  <=  I9817361d029cc98d7407cf3b8b020567[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I81ba868784103e0eb05a44d981d4d666     <=
                                             I47a6f2033a2356ac604133d12d7e0c0e[SGN_MAX_SUM_WDTH] ?
                                             ~I47a6f2033a2356ac604133d12d7e0c0e + 1 :
                                             I47a6f2033a2356ac604133d12d7e0c0e
                                             ;

            I2b7822d5d77aaed61eee87570564df76  <=  I47a6f2033a2356ac604133d12d7e0c0e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic6b88783957cbaf253648a30b22f6b1c     <=
                                             I3da1998324eb1853e5ec747b112095aa[SGN_MAX_SUM_WDTH] ?
                                             ~I3da1998324eb1853e5ec747b112095aa + 1 :
                                             I3da1998324eb1853e5ec747b112095aa
                                             ;

            Ibdad0ab78e4404c852e60a2b04c3a5f6  <=  I3da1998324eb1853e5ec747b112095aa[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4103c218a85a1d08db5c4f4b5686b2e5     <=
                                             Ic729cdba5f8a3933121a0ef35da99f8c[SGN_MAX_SUM_WDTH] ?
                                             ~Ic729cdba5f8a3933121a0ef35da99f8c + 1 :
                                             Ic729cdba5f8a3933121a0ef35da99f8c
                                             ;

            Ic4efba3932e598784f5b9ad6ad04772d  <=  Ic729cdba5f8a3933121a0ef35da99f8c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0e6c0958af503e4a120a49d02a432863     <=
                                             Id7542fd1fe3a099d7274f15c008f1cc5[SGN_MAX_SUM_WDTH] ?
                                             ~Id7542fd1fe3a099d7274f15c008f1cc5 + 1 :
                                             Id7542fd1fe3a099d7274f15c008f1cc5
                                             ;

            Ia03836a4e93d2f36513227d1dfaea0fa  <=  Id7542fd1fe3a099d7274f15c008f1cc5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f76b31e8f15c0e5fe24dcb723418111     <=
                                             I1a91347d29cd64af8941a3e042228a52[SGN_MAX_SUM_WDTH] ?
                                             ~I1a91347d29cd64af8941a3e042228a52 + 1 :
                                             I1a91347d29cd64af8941a3e042228a52
                                             ;

            I138fb0c48f2d27e3315e237d9e61d653  <=  I1a91347d29cd64af8941a3e042228a52[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id1457221b58344b60070aa026436df2c     <=
                                             Ic6b16867c426103b3e53db94469de2cb[SGN_MAX_SUM_WDTH] ?
                                             ~Ic6b16867c426103b3e53db94469de2cb + 1 :
                                             Ic6b16867c426103b3e53db94469de2cb
                                             ;

            Id0b1c46fa4caa63a4c63a44ba3c5ef8a  <=  Ic6b16867c426103b3e53db94469de2cb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icc31966508e03d8869e81d8aeb243705     <=
                                             I7361a720882c68965c1c28c2d6ba1dff[SGN_MAX_SUM_WDTH] ?
                                             ~I7361a720882c68965c1c28c2d6ba1dff + 1 :
                                             I7361a720882c68965c1c28c2d6ba1dff
                                             ;

            I3566033cf5c9a06977c9182925750707  <=  I7361a720882c68965c1c28c2d6ba1dff[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9dcccf542ba434b6e0fde6f012f98f92     <=
                                             I668a239256c66a858129b4788b0001a5[SGN_MAX_SUM_WDTH] ?
                                             ~I668a239256c66a858129b4788b0001a5 + 1 :
                                             I668a239256c66a858129b4788b0001a5
                                             ;

            I02812a8a833bb69eb168a1004b6fafdf  <=  I668a239256c66a858129b4788b0001a5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I51ccbb824a5e1e340eefd173c4491728     <=
                                             I73a72fba51f575f80ded2357a6b71af0[SGN_MAX_SUM_WDTH] ?
                                             ~I73a72fba51f575f80ded2357a6b71af0 + 1 :
                                             I73a72fba51f575f80ded2357a6b71af0
                                             ;

            Ie886c5effc85f1fe0b6411db4a2cde77  <=  I73a72fba51f575f80ded2357a6b71af0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7ae1730dcd8bc708bbfcc6a9f97ac66     <=
                                             Ief9131d8e69f733c51e9f9167ad5fa4a[SGN_MAX_SUM_WDTH] ?
                                             ~Ief9131d8e69f733c51e9f9167ad5fa4a + 1 :
                                             Ief9131d8e69f733c51e9f9167ad5fa4a
                                             ;

            Ibab1d13cd6a4f7b0c79c9f845339e53f  <=  Ief9131d8e69f733c51e9f9167ad5fa4a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4714f5c91203fcfa552f0fcf71b87442     <=
                                             I1e6904544c93f0f4bf403793e50dbf99[SGN_MAX_SUM_WDTH] ?
                                             ~I1e6904544c93f0f4bf403793e50dbf99 + 1 :
                                             I1e6904544c93f0f4bf403793e50dbf99
                                             ;

            I7b813d83b13bb7bc13940cf5714c06ba  <=  I1e6904544c93f0f4bf403793e50dbf99[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3b6d1e84fdd1019249886fa5fe65895b     <=
                                             I74f9e6de534920d70eda17b59206a4af[SGN_MAX_SUM_WDTH] ?
                                             ~I74f9e6de534920d70eda17b59206a4af + 1 :
                                             I74f9e6de534920d70eda17b59206a4af
                                             ;

            I09031235f61238b0e32ff52641aab70e  <=  I74f9e6de534920d70eda17b59206a4af[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia8a7d4207dbabc7970bf36f3fe74f72d     <=
                                             Ied74515bab35cad5e94048a9f210b7a5[SGN_MAX_SUM_WDTH] ?
                                             ~Ied74515bab35cad5e94048a9f210b7a5 + 1 :
                                             Ied74515bab35cad5e94048a9f210b7a5
                                             ;

            I5402fd208dc7ca81dfd2920a9cfa2715  <=  Ied74515bab35cad5e94048a9f210b7a5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I84047457b43ef33874f4550c3b773460     <=
                                             If38f871a7b021ceb84cdb3010d08f667[SGN_MAX_SUM_WDTH] ?
                                             ~If38f871a7b021ceb84cdb3010d08f667 + 1 :
                                             If38f871a7b021ceb84cdb3010d08f667
                                             ;

            Ia01c82761aeb124cd92fb15ee367ee8b  <=  If38f871a7b021ceb84cdb3010d08f667[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5e51563c3e69beca0b463742e6e5f9ee     <=
                                             I12a578d51082c42fcc5a9e769535ac0a[SGN_MAX_SUM_WDTH] ?
                                             ~I12a578d51082c42fcc5a9e769535ac0a + 1 :
                                             I12a578d51082c42fcc5a9e769535ac0a
                                             ;

            Ib1a40247057324b0bd810c844bf11f51  <=  I12a578d51082c42fcc5a9e769535ac0a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6c8d14e31c80811ccab1b6ab09d28089     <=
                                             I404f31fea404e730a9c4e04bec369c1a[SGN_MAX_SUM_WDTH] ?
                                             ~I404f31fea404e730a9c4e04bec369c1a + 1 :
                                             I404f31fea404e730a9c4e04bec369c1a
                                             ;

            Ied8bd4b6fd0e4fbcced6d20eb7435f55  <=  I404f31fea404e730a9c4e04bec369c1a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I50b3b7490c9b65b6e662cc86b163a2df     <=
                                             I915d15cb464b6e78cf9939232618b14c[SGN_MAX_SUM_WDTH] ?
                                             ~I915d15cb464b6e78cf9939232618b14c + 1 :
                                             I915d15cb464b6e78cf9939232618b14c
                                             ;

            I4ee312036de8c08300c358edcff1e1e9  <=  I915d15cb464b6e78cf9939232618b14c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8351a2110a3d73ad8803cf17e3317017     <=
                                             Ia8531e691cc60dcc32225eef6d8e8a2b[SGN_MAX_SUM_WDTH] ?
                                             ~Ia8531e691cc60dcc32225eef6d8e8a2b + 1 :
                                             Ia8531e691cc60dcc32225eef6d8e8a2b
                                             ;

            I477a920e2326828bf026b0a6b6a18e2b  <=  Ia8531e691cc60dcc32225eef6d8e8a2b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1e6c696951688d581f21ab2302593335     <=
                                             I5f7cd38f8b6c42a3dcc52664ea7c08a5[SGN_MAX_SUM_WDTH] ?
                                             ~I5f7cd38f8b6c42a3dcc52664ea7c08a5 + 1 :
                                             I5f7cd38f8b6c42a3dcc52664ea7c08a5
                                             ;

            Ic11a6b77b84c44180eb99220a0c4c9f6  <=  I5f7cd38f8b6c42a3dcc52664ea7c08a5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie9840e28133eebdca0be313552195c7b     <=
                                             If3f0f6acad563083949c5116ad78ce20[SGN_MAX_SUM_WDTH] ?
                                             ~If3f0f6acad563083949c5116ad78ce20 + 1 :
                                             If3f0f6acad563083949c5116ad78ce20
                                             ;

            If0970d9f7b053fce3ced3521b4885588  <=  If3f0f6acad563083949c5116ad78ce20[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I82812258a8032e273cab7139266be1b6     <=
                                             I2b8c7ab8f53d7fbda984ab8760e05fd3[SGN_MAX_SUM_WDTH] ?
                                             ~I2b8c7ab8f53d7fbda984ab8760e05fd3 + 1 :
                                             I2b8c7ab8f53d7fbda984ab8760e05fd3
                                             ;

            Ic7ebdc317c978eb275eca41d5b9106a5  <=  I2b8c7ab8f53d7fbda984ab8760e05fd3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I27ab6fd9927518e29ed36d7a7a241498     <=
                                             I29d486911dcffddec336f69b981e1e50[SGN_MAX_SUM_WDTH] ?
                                             ~I29d486911dcffddec336f69b981e1e50 + 1 :
                                             I29d486911dcffddec336f69b981e1e50
                                             ;

            Ibe3d3e6bc58efc2e9d9eb1f96cdfe424  <=  I29d486911dcffddec336f69b981e1e50[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I05b0f33a3808ac53b29d8d8309447650     <=
                                             I893881a7874f85e519089559ac4604bf[SGN_MAX_SUM_WDTH] ?
                                             ~I893881a7874f85e519089559ac4604bf + 1 :
                                             I893881a7874f85e519089559ac4604bf
                                             ;

            I1dd4671765f8826c2fe20c592c5e32c8  <=  I893881a7874f85e519089559ac4604bf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If150ebf242231f0d22c996a71552f6eb     <=
                                             I0b730d0a75cf72482ffc5b0d0267fd83[SGN_MAX_SUM_WDTH] ?
                                             ~I0b730d0a75cf72482ffc5b0d0267fd83 + 1 :
                                             I0b730d0a75cf72482ffc5b0d0267fd83
                                             ;

            I6cde57127c5bd2732e71ecb7738fad6d  <=  I0b730d0a75cf72482ffc5b0d0267fd83[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If2d0a2b58510715e74787cb60719cb5b     <=
                                             I9beb581fcdf85cc7302da093363e3b02[SGN_MAX_SUM_WDTH] ?
                                             ~I9beb581fcdf85cc7302da093363e3b02 + 1 :
                                             I9beb581fcdf85cc7302da093363e3b02
                                             ;

            If6ce2fa9f0b8bc74442ed8262b5089cf  <=  I9beb581fcdf85cc7302da093363e3b02[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib6745a6d17034a29501e022bd846bf2f     <=
                                             I0e35fb521572c6f87dbd06a8ce213337[SGN_MAX_SUM_WDTH] ?
                                             ~I0e35fb521572c6f87dbd06a8ce213337 + 1 :
                                             I0e35fb521572c6f87dbd06a8ce213337
                                             ;

            Ib0001d7298ad1f3b1c7603173a70d8b5  <=  I0e35fb521572c6f87dbd06a8ce213337[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iae09c127dfe86c9f7bdbeff447c777f5     <=
                                             Ia01e93b03cf0ff22e2f002f2e84eb9d2[SGN_MAX_SUM_WDTH] ?
                                             ~Ia01e93b03cf0ff22e2f002f2e84eb9d2 + 1 :
                                             Ia01e93b03cf0ff22e2f002f2e84eb9d2
                                             ;

            I05e739fc87e962848f265e2c73338cac  <=  Ia01e93b03cf0ff22e2f002f2e84eb9d2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I742128de6b237ed48e3a7ccd3788f0d7     <=
                                             I98a2d427581a73c639cbc9f4bf4c8802[SGN_MAX_SUM_WDTH] ?
                                             ~I98a2d427581a73c639cbc9f4bf4c8802 + 1 :
                                             I98a2d427581a73c639cbc9f4bf4c8802
                                             ;

            Iaaaf373f7e6f55214915b93da9bd71d3  <=  I98a2d427581a73c639cbc9f4bf4c8802[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id5e8fda13ba8f6d95d694d0f30da75bb     <=
                                             Ie60ba6ee53f7a01764001bc74fb90d61[SGN_MAX_SUM_WDTH] ?
                                             ~Ie60ba6ee53f7a01764001bc74fb90d61 + 1 :
                                             Ie60ba6ee53f7a01764001bc74fb90d61
                                             ;

            I47b0847946b0e00961233ac0101fa2a7  <=  Ie60ba6ee53f7a01764001bc74fb90d61[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1aa5a04e40f9b1685c77e4d101c3ccf4     <=
                                             I508e632bacf8c083a8376f73cec11bc6[SGN_MAX_SUM_WDTH] ?
                                             ~I508e632bacf8c083a8376f73cec11bc6 + 1 :
                                             I508e632bacf8c083a8376f73cec11bc6
                                             ;

            I2f23d4cdb6f5f827513aa60266936e4f  <=  I508e632bacf8c083a8376f73cec11bc6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ife1adea26d13bc299bb2de241ad4a6ea     <=
                                             I47ac3c977bbfad06ee1782b8eac6d9ec[SGN_MAX_SUM_WDTH] ?
                                             ~I47ac3c977bbfad06ee1782b8eac6d9ec + 1 :
                                             I47ac3c977bbfad06ee1782b8eac6d9ec
                                             ;

            Ia67f9b902a21de0414eb8dda52171991  <=  I47ac3c977bbfad06ee1782b8eac6d9ec[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifcf6c761f0f253921710af87ab1d2247     <=
                                             If8537bb117e0bebd25ece101a23674c8[SGN_MAX_SUM_WDTH] ?
                                             ~If8537bb117e0bebd25ece101a23674c8 + 1 :
                                             If8537bb117e0bebd25ece101a23674c8
                                             ;

            I87b10521099179c18652c86d5887c908  <=  If8537bb117e0bebd25ece101a23674c8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1478e6a9113c124bdc4361908af6643f     <=
                                             Ica8f952cb456e825c608f2e73ec9abd7[SGN_MAX_SUM_WDTH] ?
                                             ~Ica8f952cb456e825c608f2e73ec9abd7 + 1 :
                                             Ica8f952cb456e825c608f2e73ec9abd7
                                             ;

            I84057a3b319ab3d6a2ed8f2310f970fc  <=  Ica8f952cb456e825c608f2e73ec9abd7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0afd42151925883835844cf5deef6156     <=
                                             I1a332ceae6f1a640e4577c82b2bf4511[SGN_MAX_SUM_WDTH] ?
                                             ~I1a332ceae6f1a640e4577c82b2bf4511 + 1 :
                                             I1a332ceae6f1a640e4577c82b2bf4511
                                             ;

            I67d57e38df8cb35ca686ac2eb44e233e  <=  I1a332ceae6f1a640e4577c82b2bf4511[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2b4ab0aadffb3a1bb86f45ebc8acf085     <=
                                             I82c5b5deaae0b927c14adfa3b477c8df[SGN_MAX_SUM_WDTH] ?
                                             ~I82c5b5deaae0b927c14adfa3b477c8df + 1 :
                                             I82c5b5deaae0b927c14adfa3b477c8df
                                             ;

            I23955b54e486f0f0d21a2809a9472b86  <=  I82c5b5deaae0b927c14adfa3b477c8df[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iffa867719ba9c31a8756cc5e6bf81147     <=
                                             I37b08ee3258fb8359ba4c1653101e03c[SGN_MAX_SUM_WDTH] ?
                                             ~I37b08ee3258fb8359ba4c1653101e03c + 1 :
                                             I37b08ee3258fb8359ba4c1653101e03c
                                             ;

            I1e11f0088959aa40b4ad1a047b59caf4  <=  I37b08ee3258fb8359ba4c1653101e03c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibb62b6cb003f0d5549c864075f23d19b     <=
                                             I58fa785303fe60b1f1c596420aab4b5e[SGN_MAX_SUM_WDTH] ?
                                             ~I58fa785303fe60b1f1c596420aab4b5e + 1 :
                                             I58fa785303fe60b1f1c596420aab4b5e
                                             ;

            I68c35d63dc95baff41b4dc27a86d2342  <=  I58fa785303fe60b1f1c596420aab4b5e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3690d101ae99f258cc58b4482cc378c8     <=
                                             I1ceca376c3f4cd24c22cf8672c9343ba[SGN_MAX_SUM_WDTH] ?
                                             ~I1ceca376c3f4cd24c22cf8672c9343ba + 1 :
                                             I1ceca376c3f4cd24c22cf8672c9343ba
                                             ;

            I837183265ee22d080e81fea468ab0887  <=  I1ceca376c3f4cd24c22cf8672c9343ba[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id597e95ce8a168ab67890085a26870d0     <=
                                             Ieca948a12a0806b9fd483ace71c8b98e[SGN_MAX_SUM_WDTH] ?
                                             ~Ieca948a12a0806b9fd483ace71c8b98e + 1 :
                                             Ieca948a12a0806b9fd483ace71c8b98e
                                             ;

            I413b1c1985a6c9c6f202e85ff901e3a8  <=  Ieca948a12a0806b9fd483ace71c8b98e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I98df60eb8f65641f9cccce4023be905c     <=
                                             Icd2579fee72faaa432876ec8fa124d40[SGN_MAX_SUM_WDTH] ?
                                             ~Icd2579fee72faaa432876ec8fa124d40 + 1 :
                                             Icd2579fee72faaa432876ec8fa124d40
                                             ;

            Ic32c6734132776c290155a80025fe366  <=  Icd2579fee72faaa432876ec8fa124d40[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibcb4fbdee372353b79c460cdeafdfe4e     <=
                                             Iec4164641d5b71630d9d5aefb1ed5676[SGN_MAX_SUM_WDTH] ?
                                             ~Iec4164641d5b71630d9d5aefb1ed5676 + 1 :
                                             Iec4164641d5b71630d9d5aefb1ed5676
                                             ;

            I624958486d181501c7a8ec2642cb503c  <=  Iec4164641d5b71630d9d5aefb1ed5676[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I74dbf75966d047a4a9e91c1bc793666f     <=
                                             Ie43841b2ee3b5369c3863417b60e5851[SGN_MAX_SUM_WDTH] ?
                                             ~Ie43841b2ee3b5369c3863417b60e5851 + 1 :
                                             Ie43841b2ee3b5369c3863417b60e5851
                                             ;

            I04864c28351edb33b61a103add6fb875  <=  Ie43841b2ee3b5369c3863417b60e5851[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I79b8d9f9447c4c1b551ec6c1e8903040     <=
                                             I1e7346a531973e40fb2582a68f96e383[SGN_MAX_SUM_WDTH] ?
                                             ~I1e7346a531973e40fb2582a68f96e383 + 1 :
                                             I1e7346a531973e40fb2582a68f96e383
                                             ;

            Ida3dd5e990ce3c237e9628a9a090901e  <=  I1e7346a531973e40fb2582a68f96e383[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib34b66548621fabe0753223712b1369f     <=
                                             I53b62438d1bb777cf10761bf95b22718[SGN_MAX_SUM_WDTH] ?
                                             ~I53b62438d1bb777cf10761bf95b22718 + 1 :
                                             I53b62438d1bb777cf10761bf95b22718
                                             ;

            Id182a776b03f48fb139c28194ae7ab6b  <=  I53b62438d1bb777cf10761bf95b22718[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie5b3eb4c00bedfaecc3215d43ff28362     <=
                                             I6b8a0d9d8fe6ac6fa08c495b0d0d5264[SGN_MAX_SUM_WDTH] ?
                                             ~I6b8a0d9d8fe6ac6fa08c495b0d0d5264 + 1 :
                                             I6b8a0d9d8fe6ac6fa08c495b0d0d5264
                                             ;

            I0c5539373b3868d0664a92157b4b4226  <=  I6b8a0d9d8fe6ac6fa08c495b0d0d5264[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icf3a1b0b6dbcf959b44379024f3c4169     <=
                                             Ibcec436bb431239047a99c495262bf87[SGN_MAX_SUM_WDTH] ?
                                             ~Ibcec436bb431239047a99c495262bf87 + 1 :
                                             Ibcec436bb431239047a99c495262bf87
                                             ;

            Ic0191941cb968bbd7644c21767423d2e  <=  Ibcec436bb431239047a99c495262bf87[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I918c2bbe7c71f8c6a07b0bad8811f4e7     <=
                                             Id9d1f164781aad87bbb332ef7c0b5113[SGN_MAX_SUM_WDTH] ?
                                             ~Id9d1f164781aad87bbb332ef7c0b5113 + 1 :
                                             Id9d1f164781aad87bbb332ef7c0b5113
                                             ;

            I163cf58b9a308e0439a8dc7c1526e6b5  <=  Id9d1f164781aad87bbb332ef7c0b5113[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iedd960a21b1c08b4a5293cff200218b3     <=
                                             I76a91ad2a7f0323b5874f857eb914d67[SGN_MAX_SUM_WDTH] ?
                                             ~I76a91ad2a7f0323b5874f857eb914d67 + 1 :
                                             I76a91ad2a7f0323b5874f857eb914d67
                                             ;

            Ie08ad9bd71329858c1742c8f571a1c36  <=  I76a91ad2a7f0323b5874f857eb914d67[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9722c28747df3a59b0ecf8200907e98     <=
                                             I9aab2781bbd57dbe4381c695f130d5b7[SGN_MAX_SUM_WDTH] ?
                                             ~I9aab2781bbd57dbe4381c695f130d5b7 + 1 :
                                             I9aab2781bbd57dbe4381c695f130d5b7
                                             ;

            I3c10d579f80bd0106506ad047d75f188  <=  I9aab2781bbd57dbe4381c695f130d5b7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib83df72c8b73a333d0699a8bbbec16be     <=
                                             I11c62ef31300f66f787bb7285596b995[SGN_MAX_SUM_WDTH] ?
                                             ~I11c62ef31300f66f787bb7285596b995 + 1 :
                                             I11c62ef31300f66f787bb7285596b995
                                             ;

            Ieca2767ac27170058499d83016447aa7  <=  I11c62ef31300f66f787bb7285596b995[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ide3798a77f709a9f694523338b081f70     <=
                                             I7e62705e1f1e7abb04ee4a94753183b4[SGN_MAX_SUM_WDTH] ?
                                             ~I7e62705e1f1e7abb04ee4a94753183b4 + 1 :
                                             I7e62705e1f1e7abb04ee4a94753183b4
                                             ;

            Ib9c194ec16f435a9357cb344cf25bdcc  <=  I7e62705e1f1e7abb04ee4a94753183b4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0a9722a805604433562f85c62b168b96     <=
                                             Ia4d8ab77dd8598d550c4b3c57f02b328[SGN_MAX_SUM_WDTH] ?
                                             ~Ia4d8ab77dd8598d550c4b3c57f02b328 + 1 :
                                             Ia4d8ab77dd8598d550c4b3c57f02b328
                                             ;

            Ic920452d5997a8477724fa78c86c0fba  <=  Ia4d8ab77dd8598d550c4b3c57f02b328[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9480ec13cd538ed03a43e56bd6264a6     <=
                                             I23c2886f2707bae85fe967379c105eb5[SGN_MAX_SUM_WDTH] ?
                                             ~I23c2886f2707bae85fe967379c105eb5 + 1 :
                                             I23c2886f2707bae85fe967379c105eb5
                                             ;

            I6eea5fde8e2517554ad6ba25018572dc  <=  I23c2886f2707bae85fe967379c105eb5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I433ecf86b7704c5552e5fb5cafe0d529     <=
                                             Idfb980ae7487145d65bdf83b97751e6f[SGN_MAX_SUM_WDTH] ?
                                             ~Idfb980ae7487145d65bdf83b97751e6f + 1 :
                                             Idfb980ae7487145d65bdf83b97751e6f
                                             ;

            I9ad2f6fd2d7f68011fc926ec9abd5c34  <=  Idfb980ae7487145d65bdf83b97751e6f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8326f0b2d25139609e2c5e466724f224     <=
                                             If7916cdab9aa2621009bc0671d985133[SGN_MAX_SUM_WDTH] ?
                                             ~If7916cdab9aa2621009bc0671d985133 + 1 :
                                             If7916cdab9aa2621009bc0671d985133
                                             ;

            Ied33f18cbb778d5ba744d249f91c950b  <=  If7916cdab9aa2621009bc0671d985133[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibbe211d9955cdf2810c9003d1fb78074     <=
                                             I1969f6d312f67452ec24690813fc07ae[SGN_MAX_SUM_WDTH] ?
                                             ~I1969f6d312f67452ec24690813fc07ae + 1 :
                                             I1969f6d312f67452ec24690813fc07ae
                                             ;

            Ibabf61085ca7af8dfc7927b3656a76f7  <=  I1969f6d312f67452ec24690813fc07ae[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If15e950b569a92b590127d0ca6f20a16     <=
                                             I6b3c96ebbba2bfe8c549caea4a266656[SGN_MAX_SUM_WDTH] ?
                                             ~I6b3c96ebbba2bfe8c549caea4a266656 + 1 :
                                             I6b3c96ebbba2bfe8c549caea4a266656
                                             ;

            Iddc5b5b4501f9f13bcaf22081e5a70f4  <=  I6b3c96ebbba2bfe8c549caea4a266656[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I03e0532841ba39eb1d4ae823c4de2f7d     <=
                                             I73172f8b4bcb0bdbe27a09cd7ec204e0[SGN_MAX_SUM_WDTH] ?
                                             ~I73172f8b4bcb0bdbe27a09cd7ec204e0 + 1 :
                                             I73172f8b4bcb0bdbe27a09cd7ec204e0
                                             ;

            I67f87fbb746dd937fffc534c596f36c4  <=  I73172f8b4bcb0bdbe27a09cd7ec204e0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1be81a7b73987ee023e396cec87312d1     <=
                                             I96acfb8f7e6c42f616a880b3657f42a9[SGN_MAX_SUM_WDTH] ?
                                             ~I96acfb8f7e6c42f616a880b3657f42a9 + 1 :
                                             I96acfb8f7e6c42f616a880b3657f42a9
                                             ;

            I45bdd0cfe107da0d57cad1333bf95e3b  <=  I96acfb8f7e6c42f616a880b3657f42a9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4ce1a767a78673590c4074f3f03bad8d     <=
                                             I5cdce64ba621df381f9efbb8b0c8e10a[SGN_MAX_SUM_WDTH] ?
                                             ~I5cdce64ba621df381f9efbb8b0c8e10a + 1 :
                                             I5cdce64ba621df381f9efbb8b0c8e10a
                                             ;

            I4d54dd2ee2f32909098d3cc2b6689220  <=  I5cdce64ba621df381f9efbb8b0c8e10a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I57806bb7da625881e68ae315543f70d6     <=
                                             I61389621065261b79f16e6dae7c7cdac[SGN_MAX_SUM_WDTH] ?
                                             ~I61389621065261b79f16e6dae7c7cdac + 1 :
                                             I61389621065261b79f16e6dae7c7cdac
                                             ;

            I7bfb4c5d9e22d1bd8811844d9c74dff8  <=  I61389621065261b79f16e6dae7c7cdac[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8b0ab476b4790150575abb06bcdce2b3     <=
                                             Ide44caca4eb1b6edc9b55c584239ff94[SGN_MAX_SUM_WDTH] ?
                                             ~Ide44caca4eb1b6edc9b55c584239ff94 + 1 :
                                             Ide44caca4eb1b6edc9b55c584239ff94
                                             ;

            Ib9d58222da98f29fa302b4896594fe26  <=  Ide44caca4eb1b6edc9b55c584239ff94[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8846a8961b7d557df4fc62dada679c33     <=
                                             I892e07e7e972dd521f273519694e4ee7[SGN_MAX_SUM_WDTH] ?
                                             ~I892e07e7e972dd521f273519694e4ee7 + 1 :
                                             I892e07e7e972dd521f273519694e4ee7
                                             ;

            Iea3e35ece9fdb3aff3b9ff5369e9a7e0  <=  I892e07e7e972dd521f273519694e4ee7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7909a0f96a92e93f95023cddc742a5eb     <=
                                             I43c8950bb200a93cec12c09af4a38dae[SGN_MAX_SUM_WDTH] ?
                                             ~I43c8950bb200a93cec12c09af4a38dae + 1 :
                                             I43c8950bb200a93cec12c09af4a38dae
                                             ;

            Ic44eab478be232721e7a43d14beca32f  <=  I43c8950bb200a93cec12c09af4a38dae[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I43ac4857544c0fb79d04e850435ef673     <=
                                             I591f0a636f176d5a398cb6ed6d67f627[SGN_MAX_SUM_WDTH] ?
                                             ~I591f0a636f176d5a398cb6ed6d67f627 + 1 :
                                             I591f0a636f176d5a398cb6ed6d67f627
                                             ;

            Ifab075b1437495268b6a3be4cb022e71  <=  I591f0a636f176d5a398cb6ed6d67f627[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia6dfa47c465325c1d9fb9b9c5ce08f01     <=
                                             I8be467496bf21fa2c46fc5db2442a339[SGN_MAX_SUM_WDTH] ?
                                             ~I8be467496bf21fa2c46fc5db2442a339 + 1 :
                                             I8be467496bf21fa2c46fc5db2442a339
                                             ;

            I2919272e9ae3996a3e1d602ff72ba86d  <=  I8be467496bf21fa2c46fc5db2442a339[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2e9eda5bea0cc3d88359ce8a7a82f21f     <=
                                             Ifa0294e878bf5a4f1c6c7cfa52c46e7d[SGN_MAX_SUM_WDTH] ?
                                             ~Ifa0294e878bf5a4f1c6c7cfa52c46e7d + 1 :
                                             Ifa0294e878bf5a4f1c6c7cfa52c46e7d
                                             ;

            Ib6fbe376477afa58bfcc17a8564f78b2  <=  Ifa0294e878bf5a4f1c6c7cfa52c46e7d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I53ec2486418e41b2ccfa8fd82777eaf0     <=
                                             I35a8b04ecb2c6d2d7bd52a64010038ff[SGN_MAX_SUM_WDTH] ?
                                             ~I35a8b04ecb2c6d2d7bd52a64010038ff + 1 :
                                             I35a8b04ecb2c6d2d7bd52a64010038ff
                                             ;

            I659322a9fd0d5eac514437b02e0491b3  <=  I35a8b04ecb2c6d2d7bd52a64010038ff[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I18387c05cef21970ecbc39c20a87aafb     <=
                                             I38629158c9fc8600b05a3e32589cbeda[SGN_MAX_SUM_WDTH] ?
                                             ~I38629158c9fc8600b05a3e32589cbeda + 1 :
                                             I38629158c9fc8600b05a3e32589cbeda
                                             ;

            Ic68f500938d80460ffdb33a0adc48298  <=  I38629158c9fc8600b05a3e32589cbeda[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2b23eae78cb925008ad59f45e80e165b     <=
                                             Ie20705331f5fabb4c9f720a5c6592c7d[SGN_MAX_SUM_WDTH] ?
                                             ~Ie20705331f5fabb4c9f720a5c6592c7d + 1 :
                                             Ie20705331f5fabb4c9f720a5c6592c7d
                                             ;

            If5ae6fbf843fdeee17945bc5ce81aec8  <=  Ie20705331f5fabb4c9f720a5c6592c7d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic69eb7677638a90b7a54389d47be46de     <=
                                             I425d66a6ead3859f364e20a797b0e4e2[SGN_MAX_SUM_WDTH] ?
                                             ~I425d66a6ead3859f364e20a797b0e4e2 + 1 :
                                             I425d66a6ead3859f364e20a797b0e4e2
                                             ;

            I94460b6ce7b776bcc5eca149eab80c26  <=  I425d66a6ead3859f364e20a797b0e4e2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8cb9a216f4da7c27f678386cb214c59d     <=
                                             I66a2577a791bae1f31c5b99b0c3f324d[SGN_MAX_SUM_WDTH] ?
                                             ~I66a2577a791bae1f31c5b99b0c3f324d + 1 :
                                             I66a2577a791bae1f31c5b99b0c3f324d
                                             ;

            I3347717ba9556e69de30ce7533d4f5a4  <=  I66a2577a791bae1f31c5b99b0c3f324d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I48cb720a6323697084ac3bbd8fcadfcb     <=
                                             I77350e171f060c2d49e50c636fab084f[SGN_MAX_SUM_WDTH] ?
                                             ~I77350e171f060c2d49e50c636fab084f + 1 :
                                             I77350e171f060c2d49e50c636fab084f
                                             ;

            I2db290170ddae8dc52ce07edaf48b365  <=  I77350e171f060c2d49e50c636fab084f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib8dc3c1885c92cdcce7fcb58d65d03e7     <=
                                             I2101d085d5e55ef5b8247de3898a80e7[SGN_MAX_SUM_WDTH] ?
                                             ~I2101d085d5e55ef5b8247de3898a80e7 + 1 :
                                             I2101d085d5e55ef5b8247de3898a80e7
                                             ;

            Idd775d9fe6fa8dbdbfb07d4071b9caa5  <=  I2101d085d5e55ef5b8247de3898a80e7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3aa51a5c758405fa6e2dbed707555b2     <=
                                             Id38879e0d52fba6818597bd60dfc2b2c[SGN_MAX_SUM_WDTH] ?
                                             ~Id38879e0d52fba6818597bd60dfc2b2c + 1 :
                                             Id38879e0d52fba6818597bd60dfc2b2c
                                             ;

            I6cbc06919b9c695d99621db6f8d768cb  <=  Id38879e0d52fba6818597bd60dfc2b2c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4d418179c859feb8bc7d750416bb1004     <=
                                             I68081efdf01e540fe5e07643a2bc3463[SGN_MAX_SUM_WDTH] ?
                                             ~I68081efdf01e540fe5e07643a2bc3463 + 1 :
                                             I68081efdf01e540fe5e07643a2bc3463
                                             ;

            I5b8a1e1a6b904b0f6822c224ee0486e3  <=  I68081efdf01e540fe5e07643a2bc3463[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If207b2adc6f668f85cb76bf54673fe18     <=
                                             I2d70e6f392396c2ee505687f5a950a6f[SGN_MAX_SUM_WDTH] ?
                                             ~I2d70e6f392396c2ee505687f5a950a6f + 1 :
                                             I2d70e6f392396c2ee505687f5a950a6f
                                             ;

            I3f5053e519a928640ae49cf4e5b39d1e  <=  I2d70e6f392396c2ee505687f5a950a6f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib08b8067ea75e210e83526ca4a37217e     <=
                                             I6e6eae8e8a955b80abb7cb722a940e27[SGN_MAX_SUM_WDTH] ?
                                             ~I6e6eae8e8a955b80abb7cb722a940e27 + 1 :
                                             I6e6eae8e8a955b80abb7cb722a940e27
                                             ;

            I7c965c047d862c973d09a81abe03a845  <=  I6e6eae8e8a955b80abb7cb722a940e27[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95b30f641cbf7bec1886643c4468017d     <=
                                             I54cfd5f12219687ba48be0c57a979add[SGN_MAX_SUM_WDTH] ?
                                             ~I54cfd5f12219687ba48be0c57a979add + 1 :
                                             I54cfd5f12219687ba48be0c57a979add
                                             ;

            I9b8023f4dced915cd52c91bc9d4ed78f  <=  I54cfd5f12219687ba48be0c57a979add[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1978531a6f8d1d25ee6d404025ec4753     <=
                                             Ifda70e49dbdc4b5511961649914ecc71[SGN_MAX_SUM_WDTH] ?
                                             ~Ifda70e49dbdc4b5511961649914ecc71 + 1 :
                                             Ifda70e49dbdc4b5511961649914ecc71
                                             ;

            Idc6b6357741c9887a9db1037ccc2d922  <=  Ifda70e49dbdc4b5511961649914ecc71[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6c9698ba88db16b8d22ccebd58cc541d     <=
                                             I0feba37f523d6c6371bd934796519c59[SGN_MAX_SUM_WDTH] ?
                                             ~I0feba37f523d6c6371bd934796519c59 + 1 :
                                             I0feba37f523d6c6371bd934796519c59
                                             ;

            Ibe97860165dc5d9a076ebd935385ae51  <=  I0feba37f523d6c6371bd934796519c59[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0d8ac5e09b200a55bf5ba6f834cc9174     <=
                                             Ibaf70dff036e0bc11df75e2a1fe4fb34[SGN_MAX_SUM_WDTH] ?
                                             ~Ibaf70dff036e0bc11df75e2a1fe4fb34 + 1 :
                                             Ibaf70dff036e0bc11df75e2a1fe4fb34
                                             ;

            I777ee54ff20d0544af18ad8a870d6915  <=  Ibaf70dff036e0bc11df75e2a1fe4fb34[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib58b7d3d77a54ff1a180c6fa5f1400e6     <=
                                             Ib00eb8856f044c3af325f0134d16a970[SGN_MAX_SUM_WDTH] ?
                                             ~Ib00eb8856f044c3af325f0134d16a970 + 1 :
                                             Ib00eb8856f044c3af325f0134d16a970
                                             ;

            Id18c5a1d4eaa73a94e699e5f9e3c3d35  <=  Ib00eb8856f044c3af325f0134d16a970[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icf6b990098b7ab91800bfcf1e643153c     <=
                                             I4e89f11e414b55e9574f5c3d79dc4506[SGN_MAX_SUM_WDTH] ?
                                             ~I4e89f11e414b55e9574f5c3d79dc4506 + 1 :
                                             I4e89f11e414b55e9574f5c3d79dc4506
                                             ;

            I72939e49bf2d9c6a84e404419fc644a1  <=  I4e89f11e414b55e9574f5c3d79dc4506[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie4308b9ac6fb6de9329ba02b1eeb0e8a     <=
                                             If25b7447f1f34072a597f70a4234a16e[SGN_MAX_SUM_WDTH] ?
                                             ~If25b7447f1f34072a597f70a4234a16e + 1 :
                                             If25b7447f1f34072a597f70a4234a16e
                                             ;

            I57b7b48f13436b19a8d6a47e014eb41f  <=  If25b7447f1f34072a597f70a4234a16e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I01d4f02a356c51d7e4e1993de0d8eebd     <=
                                             I76ae0b929aefad162304529ea04b725f[SGN_MAX_SUM_WDTH] ?
                                             ~I76ae0b929aefad162304529ea04b725f + 1 :
                                             I76ae0b929aefad162304529ea04b725f
                                             ;

            Ia3ef2f70c5abaa852586a33c505aee0d  <=  I76ae0b929aefad162304529ea04b725f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I36c351e3641b01cc43e1dd5de0a649e5     <=
                                             Idffaf5edec0ef7b25c24f3c5e636fb75[SGN_MAX_SUM_WDTH] ?
                                             ~Idffaf5edec0ef7b25c24f3c5e636fb75 + 1 :
                                             Idffaf5edec0ef7b25c24f3c5e636fb75
                                             ;

            I6d423a7d17e05a3c597ec6ef6c5a7cba  <=  Idffaf5edec0ef7b25c24f3c5e636fb75[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4fc983e94c5b8f7bafca61fb0d351c08     <=
                                             Id041de10db620915a3755358fc2d9a41[SGN_MAX_SUM_WDTH] ?
                                             ~Id041de10db620915a3755358fc2d9a41 + 1 :
                                             Id041de10db620915a3755358fc2d9a41
                                             ;

            I48e3309c61918c3991852b45d9c72ea5  <=  Id041de10db620915a3755358fc2d9a41[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1fcb82fdf96cda14a55fa6358cb62c1e     <=
                                             I92ddd31add3c914ce6b0271e77cb67a0[SGN_MAX_SUM_WDTH] ?
                                             ~I92ddd31add3c914ce6b0271e77cb67a0 + 1 :
                                             I92ddd31add3c914ce6b0271e77cb67a0
                                             ;

            I472352e7027b9df2fa957d9fd68443ff  <=  I92ddd31add3c914ce6b0271e77cb67a0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I665e54ea6bdca483149d3b7f3ee42a2b     <=
                                             If80ebbd3419cd9fd63a745412b7233b6[SGN_MAX_SUM_WDTH] ?
                                             ~If80ebbd3419cd9fd63a745412b7233b6 + 1 :
                                             If80ebbd3419cd9fd63a745412b7233b6
                                             ;

            Idbbf2ce4a30787c5f07c3b908a73da75  <=  If80ebbd3419cd9fd63a745412b7233b6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I925df2307b5af6d1b166e5435641d3bd     <=
                                             I0b67c1f8e03165404e0b76d1a05d88de[SGN_MAX_SUM_WDTH] ?
                                             ~I0b67c1f8e03165404e0b76d1a05d88de + 1 :
                                             I0b67c1f8e03165404e0b76d1a05d88de
                                             ;

            Ibc9a860879ccc58c815b9f6caa23320a  <=  I0b67c1f8e03165404e0b76d1a05d88de[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9b14f48aa357d09e460a445da86cdf89     <=
                                             If78c15d7c2dc19cef26743eccbb52e6c[SGN_MAX_SUM_WDTH] ?
                                             ~If78c15d7c2dc19cef26743eccbb52e6c + 1 :
                                             If78c15d7c2dc19cef26743eccbb52e6c
                                             ;

            Ia71cf07b645c58cffe33be1a9a960eb2  <=  If78c15d7c2dc19cef26743eccbb52e6c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I78e94ecb6c92fa8ee24edaff33b6f82d     <=
                                             I228c0b3c3919aaf70ea24874f314eaa5[SGN_MAX_SUM_WDTH] ?
                                             ~I228c0b3c3919aaf70ea24874f314eaa5 + 1 :
                                             I228c0b3c3919aaf70ea24874f314eaa5
                                             ;

            I0ceb14ac0187d804f9692e0c55b8e941  <=  I228c0b3c3919aaf70ea24874f314eaa5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5ebeb9ce5adee72a7c9527ea6d3a3028     <=
                                             I986ca3b0590709588c3d9d2274a1fd34[SGN_MAX_SUM_WDTH] ?
                                             ~I986ca3b0590709588c3d9d2274a1fd34 + 1 :
                                             I986ca3b0590709588c3d9d2274a1fd34
                                             ;

            Ief18a19d451f05f6051e3cc8de16d73c  <=  I986ca3b0590709588c3d9d2274a1fd34[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I90d7b28ec09142ca8086836fc0c5ea0d     <=
                                             I765867ea6452d51f31e96ec83f68f9df[SGN_MAX_SUM_WDTH] ?
                                             ~I765867ea6452d51f31e96ec83f68f9df + 1 :
                                             I765867ea6452d51f31e96ec83f68f9df
                                             ;

            I30be0b18e4415ca50f2d8149efaaafe6  <=  I765867ea6452d51f31e96ec83f68f9df[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I27d9985415e6d0b117e5a4c2863aa7f8     <=
                                             I6e970e7bafbfa1866203483ed18a7db7[SGN_MAX_SUM_WDTH] ?
                                             ~I6e970e7bafbfa1866203483ed18a7db7 + 1 :
                                             I6e970e7bafbfa1866203483ed18a7db7
                                             ;

            I7ec15b73b2811b44e1e50c74a9f921e9  <=  I6e970e7bafbfa1866203483ed18a7db7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idf9b563e5d10c2bdbcc07e81d74467eb     <=
                                             Ia31bbc3e099eb2180960917330d6b2e1[SGN_MAX_SUM_WDTH] ?
                                             ~Ia31bbc3e099eb2180960917330d6b2e1 + 1 :
                                             Ia31bbc3e099eb2180960917330d6b2e1
                                             ;

            I0fd2f706e374a4eb57ee26ab50201e15  <=  Ia31bbc3e099eb2180960917330d6b2e1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie351922194483938302ff6cafc477e4a     <=
                                             Ibc94d96e529274004dfed98c98915827[SGN_MAX_SUM_WDTH] ?
                                             ~Ibc94d96e529274004dfed98c98915827 + 1 :
                                             Ibc94d96e529274004dfed98c98915827
                                             ;

            I44f170d02bae7fe044456e125a98451d  <=  Ibc94d96e529274004dfed98c98915827[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifb2da5faf236ca8636677bc1dc35c4db     <=
                                             I60eb0a19c8d75780a4dae7d33ba46bd4[SGN_MAX_SUM_WDTH] ?
                                             ~I60eb0a19c8d75780a4dae7d33ba46bd4 + 1 :
                                             I60eb0a19c8d75780a4dae7d33ba46bd4
                                             ;

            I30c0fcd89e0cc7c5fa348df7b4fa2ccf  <=  I60eb0a19c8d75780a4dae7d33ba46bd4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie15825d216685ae241b528fa9c158ff3     <=
                                             I701ff10dac46e4482b3bcaa387c9a725[SGN_MAX_SUM_WDTH] ?
                                             ~I701ff10dac46e4482b3bcaa387c9a725 + 1 :
                                             I701ff10dac46e4482b3bcaa387c9a725
                                             ;

            I13a98f98c54b2e412cd88c96f016c41b  <=  I701ff10dac46e4482b3bcaa387c9a725[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id92c2d8bc61245c0c8e40bec2424c3c8     <=
                                             Ifd170f2b9fa5df9a7d0817307b5586a2[SGN_MAX_SUM_WDTH] ?
                                             ~Ifd170f2b9fa5df9a7d0817307b5586a2 + 1 :
                                             Ifd170f2b9fa5df9a7d0817307b5586a2
                                             ;

            I9890f7fc708c7b8cf460849b4a30025b  <=  Ifd170f2b9fa5df9a7d0817307b5586a2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icd9fd8d7114b6e894dbee493b6797df6     <=
                                             Ia5feb8ce451f12382cb66853e948047d[SGN_MAX_SUM_WDTH] ?
                                             ~Ia5feb8ce451f12382cb66853e948047d + 1 :
                                             Ia5feb8ce451f12382cb66853e948047d
                                             ;

            I5e69e930a318dcb0594a823b3129d650  <=  Ia5feb8ce451f12382cb66853e948047d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I29ff688c085f2b18e7a3af969f18af76     <=
                                             I3a971f30fe10de02e604402b55c181da[SGN_MAX_SUM_WDTH] ?
                                             ~I3a971f30fe10de02e604402b55c181da + 1 :
                                             I3a971f30fe10de02e604402b55c181da
                                             ;

            I403303228c0df825f67436f4a7e64061  <=  I3a971f30fe10de02e604402b55c181da[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6d56db9fcfe69dfcd747521a1ff62297     <=
                                             I3350d782125dfaa1c32d06e6ede68e0f[SGN_MAX_SUM_WDTH] ?
                                             ~I3350d782125dfaa1c32d06e6ede68e0f + 1 :
                                             I3350d782125dfaa1c32d06e6ede68e0f
                                             ;

            I946246be5b4745508b7d4b578f83aaa2  <=  I3350d782125dfaa1c32d06e6ede68e0f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2f17f7c79a0118b39a63894917c6affa     <=
                                             Ia07581cdc470c8ba833acbc8a58f7d0e[SGN_MAX_SUM_WDTH] ?
                                             ~Ia07581cdc470c8ba833acbc8a58f7d0e + 1 :
                                             Ia07581cdc470c8ba833acbc8a58f7d0e
                                             ;

            I95f0acd4f955058041c035789c3a4d99  <=  Ia07581cdc470c8ba833acbc8a58f7d0e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7350af5d5ee09ad28c459e3674a829ab     <=
                                             Id91d824405f52636dc30344bf8c088ec[SGN_MAX_SUM_WDTH] ?
                                             ~Id91d824405f52636dc30344bf8c088ec + 1 :
                                             Id91d824405f52636dc30344bf8c088ec
                                             ;

            I4082b3564c1949a19ed35bd5a88e1ef4  <=  Id91d824405f52636dc30344bf8c088ec[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I67b6415c5135e3d6a41d56d98d3f8315     <=
                                             I36beed9320665d5988556ea089ee26f8[SGN_MAX_SUM_WDTH] ?
                                             ~I36beed9320665d5988556ea089ee26f8 + 1 :
                                             I36beed9320665d5988556ea089ee26f8
                                             ;

            Ia7606050c683ecefc510ba92ac539a9c  <=  I36beed9320665d5988556ea089ee26f8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4a6fffd8bb7244599383f2aa3a1c8916     <=
                                             If05d018c797e7d4348fe5bd5423b23cb[SGN_MAX_SUM_WDTH] ?
                                             ~If05d018c797e7d4348fe5bd5423b23cb + 1 :
                                             If05d018c797e7d4348fe5bd5423b23cb
                                             ;

            I5446c1c323774715371c73bd1be66697  <=  If05d018c797e7d4348fe5bd5423b23cb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7dbcd21016231546b76aab175cac9f74     <=
                                             Ia78ed58e20602b99c01f2208cec79dfd[SGN_MAX_SUM_WDTH] ?
                                             ~Ia78ed58e20602b99c01f2208cec79dfd + 1 :
                                             Ia78ed58e20602b99c01f2208cec79dfd
                                             ;

            I3a8e9e7d2cd6751e8500a5567cef5acc  <=  Ia78ed58e20602b99c01f2208cec79dfd[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9aeff3dc44ed0d0f32518590a900dcc9     <=
                                             I229890d0e3576523fabea29f8594a853[SGN_MAX_SUM_WDTH] ?
                                             ~I229890d0e3576523fabea29f8594a853 + 1 :
                                             I229890d0e3576523fabea29f8594a853
                                             ;

            I621b20d29d3a9a9f41065bc3c3bbd2d8  <=  I229890d0e3576523fabea29f8594a853[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I988b7d5d56d22d2c77c5c8c125129a50     <=
                                             I3f0ac12bf9d4014f5418383146bcc1ab[SGN_MAX_SUM_WDTH] ?
                                             ~I3f0ac12bf9d4014f5418383146bcc1ab + 1 :
                                             I3f0ac12bf9d4014f5418383146bcc1ab
                                             ;

            I263aad78110a1136eb7012c6983b2a8d  <=  I3f0ac12bf9d4014f5418383146bcc1ab[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iff35cd97f2a6d37a7861b9cc1a655ef5     <=
                                             I38e35040b0a7e5476f308d265b7fbf67[SGN_MAX_SUM_WDTH] ?
                                             ~I38e35040b0a7e5476f308d265b7fbf67 + 1 :
                                             I38e35040b0a7e5476f308d265b7fbf67
                                             ;

            If4308ed204e33952c9931f8fe257aca4  <=  I38e35040b0a7e5476f308d265b7fbf67[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifb3f2a1bedfe41c73d198046a2a3f177     <=
                                             I90c35b33579355f50d23995dc25cc2af[SGN_MAX_SUM_WDTH] ?
                                             ~I90c35b33579355f50d23995dc25cc2af + 1 :
                                             I90c35b33579355f50d23995dc25cc2af
                                             ;

            Iddcfab4a7022e0f12fd20cb34e9b9d02  <=  I90c35b33579355f50d23995dc25cc2af[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I37ddc6ccbc188a3eb8c33a501de820be     <=
                                             I19a71e86490479795328e31521b6b842[SGN_MAX_SUM_WDTH] ?
                                             ~I19a71e86490479795328e31521b6b842 + 1 :
                                             I19a71e86490479795328e31521b6b842
                                             ;

            I759409e242eaeb144a53e630a8cfd514  <=  I19a71e86490479795328e31521b6b842[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica608f1136da397e2ab61bd4a5d83201     <=
                                             I5505d84d5ef89111fd375ce986e33c52[SGN_MAX_SUM_WDTH] ?
                                             ~I5505d84d5ef89111fd375ce986e33c52 + 1 :
                                             I5505d84d5ef89111fd375ce986e33c52
                                             ;

            I5f96a68d20e3ebc71dad4b43305baa20  <=  I5505d84d5ef89111fd375ce986e33c52[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I80636a3df4541bf29780bcb4d0ee48f9     <=
                                             Ie47404148e49f0bfa2775b3573dee999[SGN_MAX_SUM_WDTH] ?
                                             ~Ie47404148e49f0bfa2775b3573dee999 + 1 :
                                             Ie47404148e49f0bfa2775b3573dee999
                                             ;

            I5d92fdff96b9cd64f3af2b28b13e9956  <=  Ie47404148e49f0bfa2775b3573dee999[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ad99d544187db3cc7090b92c9933a31     <=
                                             Ibae1afc3891aaf6fa2751a693cbf5e1c[SGN_MAX_SUM_WDTH] ?
                                             ~Ibae1afc3891aaf6fa2751a693cbf5e1c + 1 :
                                             Ibae1afc3891aaf6fa2751a693cbf5e1c
                                             ;

            Iab2f643f81921ed8464e1bbd9fa8c68e  <=  Ibae1afc3891aaf6fa2751a693cbf5e1c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iaa8a2b6fcd469869efcf0b75ca38e68f     <=
                                             Icbc45a900f0692fde798caa8c1b9b223[SGN_MAX_SUM_WDTH] ?
                                             ~Icbc45a900f0692fde798caa8c1b9b223 + 1 :
                                             Icbc45a900f0692fde798caa8c1b9b223
                                             ;

            I17d7f36fdade16dbcf621fe302bd7e57  <=  Icbc45a900f0692fde798caa8c1b9b223[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9a171d2d8eee362a0073ab7b139d3037     <=
                                             Ib8aaa1d409ba2d09187c3cf4ad4a1fec[SGN_MAX_SUM_WDTH] ?
                                             ~Ib8aaa1d409ba2d09187c3cf4ad4a1fec + 1 :
                                             Ib8aaa1d409ba2d09187c3cf4ad4a1fec
                                             ;

            I23afd747ecece714e32fbb896b5c022a  <=  Ib8aaa1d409ba2d09187c3cf4ad4a1fec[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I84cdcba86bc5991feb391003cd7be40b     <=
                                             I6a97c95991e02e0e36ec0a1f7c006626[SGN_MAX_SUM_WDTH] ?
                                             ~I6a97c95991e02e0e36ec0a1f7c006626 + 1 :
                                             I6a97c95991e02e0e36ec0a1f7c006626
                                             ;

            I388528eaf83566cc56b23485a9c05962  <=  I6a97c95991e02e0e36ec0a1f7c006626[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9e5c3a848acce5daf570458f78f6aad     <=
                                             I30c34fb37caafa3e5870ae3ee43693c1[SGN_MAX_SUM_WDTH] ?
                                             ~I30c34fb37caafa3e5870ae3ee43693c1 + 1 :
                                             I30c34fb37caafa3e5870ae3ee43693c1
                                             ;

            Iea424dd9d8916c4951b8746408b8a521  <=  I30c34fb37caafa3e5870ae3ee43693c1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I73247d4348333f67a491fc607b15af0e     <=
                                             I8f23d2c62e919062678a00aa98eff7ea[SGN_MAX_SUM_WDTH] ?
                                             ~I8f23d2c62e919062678a00aa98eff7ea + 1 :
                                             I8f23d2c62e919062678a00aa98eff7ea
                                             ;

            I73bbf90b625d56f663ad10f9d21d8e76  <=  I8f23d2c62e919062678a00aa98eff7ea[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I021c745eee4b85a2cd91d9d8d2b18b2c     <=
                                             Iaddc9a87ebf5cfb7bbabe07260c592b1[SGN_MAX_SUM_WDTH] ?
                                             ~Iaddc9a87ebf5cfb7bbabe07260c592b1 + 1 :
                                             Iaddc9a87ebf5cfb7bbabe07260c592b1
                                             ;

            I41796b587316c600bf583edc62649bd8  <=  Iaddc9a87ebf5cfb7bbabe07260c592b1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1381c0a0bd28b1c5542992084635b355     <=
                                             I24abea8ce306ff137aabea504932da94[SGN_MAX_SUM_WDTH] ?
                                             ~I24abea8ce306ff137aabea504932da94 + 1 :
                                             I24abea8ce306ff137aabea504932da94
                                             ;

            I7009c18515dd43d8dd2e5d1ee6779641  <=  I24abea8ce306ff137aabea504932da94[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie74eeddc21428254a8fc4c3e293b5eb7     <=
                                             Ibee212f9caef9ff8a725aa08e2e955bf[SGN_MAX_SUM_WDTH] ?
                                             ~Ibee212f9caef9ff8a725aa08e2e955bf + 1 :
                                             Ibee212f9caef9ff8a725aa08e2e955bf
                                             ;

            I797c9cb725f88c07be28f017871d17f8  <=  Ibee212f9caef9ff8a725aa08e2e955bf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib1d0f94258b45de4bfe610086d8990c5     <=
                                             Ie62effeaea232e1a8a50ac3f744f3f3b[SGN_MAX_SUM_WDTH] ?
                                             ~Ie62effeaea232e1a8a50ac3f744f3f3b + 1 :
                                             Ie62effeaea232e1a8a50ac3f744f3f3b
                                             ;

            I06b48093d4c9b0327c3efc6fa4ca7daf  <=  Ie62effeaea232e1a8a50ac3f744f3f3b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I138d6d5d60df37870cdbb1d9c51a94af     <=
                                             I6712564d12398f5407fade724db8792c[SGN_MAX_SUM_WDTH] ?
                                             ~I6712564d12398f5407fade724db8792c + 1 :
                                             I6712564d12398f5407fade724db8792c
                                             ;

            I04c734eb876aa722e84d6b9edd297978  <=  I6712564d12398f5407fade724db8792c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I706378735e63e15c8d5395446ea41db8     <=
                                             I5a699ad31ee84bb49eff73572bcaf84a[SGN_MAX_SUM_WDTH] ?
                                             ~I5a699ad31ee84bb49eff73572bcaf84a + 1 :
                                             I5a699ad31ee84bb49eff73572bcaf84a
                                             ;

            Ifb89e7ad8ef661959d82b7c22f187243  <=  I5a699ad31ee84bb49eff73572bcaf84a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If8680a7fc4f5532a660006bf4ca6a66e     <=
                                             I63f0b04113e2c8b0cf0474f8aa4fc1cb[SGN_MAX_SUM_WDTH] ?
                                             ~I63f0b04113e2c8b0cf0474f8aa4fc1cb + 1 :
                                             I63f0b04113e2c8b0cf0474f8aa4fc1cb
                                             ;

            Id1dce2b9eafc35fa71df33ada4aac539  <=  I63f0b04113e2c8b0cf0474f8aa4fc1cb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic59d1ff3051a95166c3c2d5a2881221b     <=
                                             I0dd55598c5774df690bb002eefd62dae[SGN_MAX_SUM_WDTH] ?
                                             ~I0dd55598c5774df690bb002eefd62dae + 1 :
                                             I0dd55598c5774df690bb002eefd62dae
                                             ;

            Ied19cb51636bfb029ba8a2c390f97105  <=  I0dd55598c5774df690bb002eefd62dae[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I54a551af28c505601cdfaf8faaa94afb     <=
                                             I361cee04efb7ccdb28fbf44a7f9c3467[SGN_MAX_SUM_WDTH] ?
                                             ~I361cee04efb7ccdb28fbf44a7f9c3467 + 1 :
                                             I361cee04efb7ccdb28fbf44a7f9c3467
                                             ;

            Ie46b71f55aef4d00168202431d47dce0  <=  I361cee04efb7ccdb28fbf44a7f9c3467[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6a3124c03eb83d41c16704133bd1cfde     <=
                                             I26225a10fd6209094b91ed34531ca2b4[SGN_MAX_SUM_WDTH] ?
                                             ~I26225a10fd6209094b91ed34531ca2b4 + 1 :
                                             I26225a10fd6209094b91ed34531ca2b4
                                             ;

            I8c0c1a0a35f4f7a688f516c567242d39  <=  I26225a10fd6209094b91ed34531ca2b4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie9ee27b9761af611ab96f0010abd47a3     <=
                                             Ib269184699c52eafef7d54ca1fda31d7[SGN_MAX_SUM_WDTH] ?
                                             ~Ib269184699c52eafef7d54ca1fda31d7 + 1 :
                                             Ib269184699c52eafef7d54ca1fda31d7
                                             ;

            I53222c82827cab7c770e057ae91bc10e  <=  Ib269184699c52eafef7d54ca1fda31d7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I305436919f84066a22ab1417ebabd737     <=
                                             I586e24737da989e9591444e6d260cc9c[SGN_MAX_SUM_WDTH] ?
                                             ~I586e24737da989e9591444e6d260cc9c + 1 :
                                             I586e24737da989e9591444e6d260cc9c
                                             ;

            I8015717cd36aabbf2cf4aa3a5c234690  <=  I586e24737da989e9591444e6d260cc9c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I78e63717f436493b756efa32d66cdefd     <=
                                             I01fe0c5ce70d18bdced623e1bfeb55c4[SGN_MAX_SUM_WDTH] ?
                                             ~I01fe0c5ce70d18bdced623e1bfeb55c4 + 1 :
                                             I01fe0c5ce70d18bdced623e1bfeb55c4
                                             ;

            Ic0c13c9a929c8c46e8702cef74de8955  <=  I01fe0c5ce70d18bdced623e1bfeb55c4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic965ba971642db19ca773eb68dc0b9bf     <=
                                             I31e6b870600dcb417653fd673d0c1a55[SGN_MAX_SUM_WDTH] ?
                                             ~I31e6b870600dcb417653fd673d0c1a55 + 1 :
                                             I31e6b870600dcb417653fd673d0c1a55
                                             ;

            I71d7f72d83b7410de31e09ea96adb95c  <=  I31e6b870600dcb417653fd673d0c1a55[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I579480a66a5f6331fb46de13090ce888     <=
                                             Id79c1fa529c3b719ef4534d1c3abc975[SGN_MAX_SUM_WDTH] ?
                                             ~Id79c1fa529c3b719ef4534d1c3abc975 + 1 :
                                             Id79c1fa529c3b719ef4534d1c3abc975
                                             ;

            I1db4ea6916125702e7fb09d0f742e60a  <=  Id79c1fa529c3b719ef4534d1c3abc975[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I38d78b447217271a63f30f78b424e2ae     <=
                                             I496765810959107754d8f764be715da4[SGN_MAX_SUM_WDTH] ?
                                             ~I496765810959107754d8f764be715da4 + 1 :
                                             I496765810959107754d8f764be715da4
                                             ;

            Idc445d3f5b3b62562b0ac83e5f17e92a  <=  I496765810959107754d8f764be715da4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4c8d7e5474b19a7c63444d0cb6143728     <=
                                             If1b62fde8c7b6aa858dff5eba22d51a8[SGN_MAX_SUM_WDTH] ?
                                             ~If1b62fde8c7b6aa858dff5eba22d51a8 + 1 :
                                             If1b62fde8c7b6aa858dff5eba22d51a8
                                             ;

            Iee6e52d75c093a24eb4e5e0b45feb256  <=  If1b62fde8c7b6aa858dff5eba22d51a8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia4bc4b7414bf31305ec8f63e7eda61e7     <=
                                             I5a86b5c97d7b531c201169167a720d2b[SGN_MAX_SUM_WDTH] ?
                                             ~I5a86b5c97d7b531c201169167a720d2b + 1 :
                                             I5a86b5c97d7b531c201169167a720d2b
                                             ;

            Id48fe0672aa98f987162931527e9f9bc  <=  I5a86b5c97d7b531c201169167a720d2b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibbebe287d56c7d627f3ffcf706575e77     <=
                                             I8e0d580b0f875a9373a3d8fb5523183d[SGN_MAX_SUM_WDTH] ?
                                             ~I8e0d580b0f875a9373a3d8fb5523183d + 1 :
                                             I8e0d580b0f875a9373a3d8fb5523183d
                                             ;

            Idce46f6d03376bea1ba361e8c59f8bd1  <=  I8e0d580b0f875a9373a3d8fb5523183d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I83867e6ee369fff7e39ef5c8d5398fef     <=
                                             I0a35c9a4f7596b64d8a6e39878fbc83a[SGN_MAX_SUM_WDTH] ?
                                             ~I0a35c9a4f7596b64d8a6e39878fbc83a + 1 :
                                             I0a35c9a4f7596b64d8a6e39878fbc83a
                                             ;

            Ie79ce8adeef2c3c24a3386f054d0cf5b  <=  I0a35c9a4f7596b64d8a6e39878fbc83a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1d40df7dbf99674f987bd06db714a702     <=
                                             I9eed09a7c7b86123ee154b783cb7e720[SGN_MAX_SUM_WDTH] ?
                                             ~I9eed09a7c7b86123ee154b783cb7e720 + 1 :
                                             I9eed09a7c7b86123ee154b783cb7e720
                                             ;

            I0d41bef808860bde56d48792764612d5  <=  I9eed09a7c7b86123ee154b783cb7e720[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I92f42789cb81760ff2973e3a5fe915c3     <=
                                             I45efcc842b324efcbf828c6d68f19e84[SGN_MAX_SUM_WDTH] ?
                                             ~I45efcc842b324efcbf828c6d68f19e84 + 1 :
                                             I45efcc842b324efcbf828c6d68f19e84
                                             ;

            Ib6ae81df8db1dae269437861ee11ec0d  <=  I45efcc842b324efcbf828c6d68f19e84[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idbd5f2a25ab05808721cf9c403017565     <=
                                             I4922b2f4381eb54d365a270b32c944c0[SGN_MAX_SUM_WDTH] ?
                                             ~I4922b2f4381eb54d365a270b32c944c0 + 1 :
                                             I4922b2f4381eb54d365a270b32c944c0
                                             ;

            I33ddee677715877c11a1df45cbfb01ac  <=  I4922b2f4381eb54d365a270b32c944c0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7ca5f07d6d3c2a045dfd55ae5214dd65     <=
                                             Ica29fa9ccbb761ae142e6ae7186aa830[SGN_MAX_SUM_WDTH] ?
                                             ~Ica29fa9ccbb761ae142e6ae7186aa830 + 1 :
                                             Ica29fa9ccbb761ae142e6ae7186aa830
                                             ;

            I433dd5092cf1851cd196feade3cfa6d8  <=  Ica29fa9ccbb761ae142e6ae7186aa830[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7f4e1445c68abbadce23944b99d206f9     <=
                                             Ie1e5ff68116424c122e4763955e243ac[SGN_MAX_SUM_WDTH] ?
                                             ~Ie1e5ff68116424c122e4763955e243ac + 1 :
                                             Ie1e5ff68116424c122e4763955e243ac
                                             ;

            I71d3a999d88e591e102398409b3adebf  <=  Ie1e5ff68116424c122e4763955e243ac[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id9f28016678e5e2127d9f0aa93e0b534     <=
                                             I1c817dbc1d0d04ab8d417d31ef477daf[SGN_MAX_SUM_WDTH] ?
                                             ~I1c817dbc1d0d04ab8d417d31ef477daf + 1 :
                                             I1c817dbc1d0d04ab8d417d31ef477daf
                                             ;

            Iebecd2d19f9174d87deedc1a273e7baa  <=  I1c817dbc1d0d04ab8d417d31ef477daf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6b939c57a8b7c7c51ab43e1b1df12f6a     <=
                                             Id4bf2c50adae02e36a8c7a862a470efb[SGN_MAX_SUM_WDTH] ?
                                             ~Id4bf2c50adae02e36a8c7a862a470efb + 1 :
                                             Id4bf2c50adae02e36a8c7a862a470efb
                                             ;

            I168afc1863f909dbcb6a9230db9f3e00  <=  Id4bf2c50adae02e36a8c7a862a470efb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic5d0df586d56bf4cb322d4c3ad677385     <=
                                             I11f3867bc6c57b2f58b19c0ffbbc0827[SGN_MAX_SUM_WDTH] ?
                                             ~I11f3867bc6c57b2f58b19c0ffbbc0827 + 1 :
                                             I11f3867bc6c57b2f58b19c0ffbbc0827
                                             ;

            I1c4b29e48d0effac4839037ae5688334  <=  I11f3867bc6c57b2f58b19c0ffbbc0827[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2e287724873cf6761799eaf464ed6302     <=
                                             I630f6f37116aab84814e74017b6d3c4c[SGN_MAX_SUM_WDTH] ?
                                             ~I630f6f37116aab84814e74017b6d3c4c + 1 :
                                             I630f6f37116aab84814e74017b6d3c4c
                                             ;

            I431fc2e9533012c8571d8158d4777dea  <=  I630f6f37116aab84814e74017b6d3c4c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia7a10cffe31a53aafa1104b97543280b     <=
                                             I3b0edd5d01b89026be06cf00b6eca7c0[SGN_MAX_SUM_WDTH] ?
                                             ~I3b0edd5d01b89026be06cf00b6eca7c0 + 1 :
                                             I3b0edd5d01b89026be06cf00b6eca7c0
                                             ;

            Ief72606c77113ae37845e4aa4a2ae5e7  <=  I3b0edd5d01b89026be06cf00b6eca7c0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ieeb089c6a18791a2227c8571913d689a     <=
                                             Ifad4e44440835f78f56065a3aa29ad3f[SGN_MAX_SUM_WDTH] ?
                                             ~Ifad4e44440835f78f56065a3aa29ad3f + 1 :
                                             Ifad4e44440835f78f56065a3aa29ad3f
                                             ;

            I641539560711ff1824bd90baa0f21f96  <=  Ifad4e44440835f78f56065a3aa29ad3f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib29b00328971c3cd67209a5ea5b63b0a     <=
                                             I93a1ba64d41cef26b742ba06755d77a1[SGN_MAX_SUM_WDTH] ?
                                             ~I93a1ba64d41cef26b742ba06755d77a1 + 1 :
                                             I93a1ba64d41cef26b742ba06755d77a1
                                             ;

            I3ac0799861144b599995318bdade2114  <=  I93a1ba64d41cef26b742ba06755d77a1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I517e0868f2bb9a22c287a1f3eeaad2f3     <=
                                             Ib2531654b83ce43d8f11a08c36cca4f7[SGN_MAX_SUM_WDTH] ?
                                             ~Ib2531654b83ce43d8f11a08c36cca4f7 + 1 :
                                             Ib2531654b83ce43d8f11a08c36cca4f7
                                             ;

            Ie83fa8157a7cce44c2e25f46ce897dbb  <=  Ib2531654b83ce43d8f11a08c36cca4f7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2bc9f76469e2a3f9846560ad1975cf54     <=
                                             I984fc2e5cd03bcf452fd7eb62be1b5b6[SGN_MAX_SUM_WDTH] ?
                                             ~I984fc2e5cd03bcf452fd7eb62be1b5b6 + 1 :
                                             I984fc2e5cd03bcf452fd7eb62be1b5b6
                                             ;

            I8be4711146486fea913843e497065b50  <=  I984fc2e5cd03bcf452fd7eb62be1b5b6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9f089315e435cd69d2929fdd936a8a77     <=
                                             Ide09ff97f4d7b3049872064c78fd2b14[SGN_MAX_SUM_WDTH] ?
                                             ~Ide09ff97f4d7b3049872064c78fd2b14 + 1 :
                                             Ide09ff97f4d7b3049872064c78fd2b14
                                             ;

            I65171c9ee8449407484e5c82d13c6751  <=  Ide09ff97f4d7b3049872064c78fd2b14[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9b54c9fb4179423c731217286e329930     <=
                                             I99c143788bcb9dfcb14e29b1f9117770[SGN_MAX_SUM_WDTH] ?
                                             ~I99c143788bcb9dfcb14e29b1f9117770 + 1 :
                                             I99c143788bcb9dfcb14e29b1f9117770
                                             ;

            I7353ebf3a1cde89d2bb3fa667f7f5485  <=  I99c143788bcb9dfcb14e29b1f9117770[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I82fb41ab743146badfd2e82258afb310     <=
                                             I4c4a40069ce9f6b40b8a1ec7787cade1[SGN_MAX_SUM_WDTH] ?
                                             ~I4c4a40069ce9f6b40b8a1ec7787cade1 + 1 :
                                             I4c4a40069ce9f6b40b8a1ec7787cade1
                                             ;

            I669d34b955d2991ebbb31c149ad1b6f8  <=  I4c4a40069ce9f6b40b8a1ec7787cade1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5619b91de99eead78befdcba1c62411e     <=
                                             I5a345140c4181b5307ea3c5b79e62b11[SGN_MAX_SUM_WDTH] ?
                                             ~I5a345140c4181b5307ea3c5b79e62b11 + 1 :
                                             I5a345140c4181b5307ea3c5b79e62b11
                                             ;

            Iabb01dc9980b4879a7356712b51df0d6  <=  I5a345140c4181b5307ea3c5b79e62b11[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I83dd2047dece99cd841b2e7955819d57     <=
                                             Ib9e2a08275b9e2571238c39945aba5d2[SGN_MAX_SUM_WDTH] ?
                                             ~Ib9e2a08275b9e2571238c39945aba5d2 + 1 :
                                             Ib9e2a08275b9e2571238c39945aba5d2
                                             ;

            I373841aa2bcbad8232d54ac9035a3ef9  <=  Ib9e2a08275b9e2571238c39945aba5d2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8c927e66ccbf4d19f07af5ef9fbfe3fb     <=
                                             I203718fd22ec9e6e4ac7a9c1973d6837[SGN_MAX_SUM_WDTH] ?
                                             ~I203718fd22ec9e6e4ac7a9c1973d6837 + 1 :
                                             I203718fd22ec9e6e4ac7a9c1973d6837
                                             ;

            Ib6124faff821158c6a2c9a9c454ab68c  <=  I203718fd22ec9e6e4ac7a9c1973d6837[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0793fa8938acdf65486e5582d01b9e5a     <=
                                             I8fa60b209a1ac0d2738e58662612206f[SGN_MAX_SUM_WDTH] ?
                                             ~I8fa60b209a1ac0d2738e58662612206f + 1 :
                                             I8fa60b209a1ac0d2738e58662612206f
                                             ;

            I6f7a45fe64ffeda9ed120be3a4519aea  <=  I8fa60b209a1ac0d2738e58662612206f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ied68d7ba0ee9974eb33767e737760b4d     <=
                                             I579c31eb0b51668db2b1edb1f10a372f[SGN_MAX_SUM_WDTH] ?
                                             ~I579c31eb0b51668db2b1edb1f10a372f + 1 :
                                             I579c31eb0b51668db2b1edb1f10a372f
                                             ;

            Id1dafb7e45b860d506e0c2c91b28142e  <=  I579c31eb0b51668db2b1edb1f10a372f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I95ba37056659b29fd4318a68d85445e8     <=
                                             I425545d21b0a9447b41481b5874c6a26[SGN_MAX_SUM_WDTH] ?
                                             ~I425545d21b0a9447b41481b5874c6a26 + 1 :
                                             I425545d21b0a9447b41481b5874c6a26
                                             ;

            I5f1609647f1e71cef4ba2d605c6c8445  <=  I425545d21b0a9447b41481b5874c6a26[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I08d7051a18f358d08728f1c401c15c47     <=
                                             I2d1670c45bd1cc15172a12175f7fb906[SGN_MAX_SUM_WDTH] ?
                                             ~I2d1670c45bd1cc15172a12175f7fb906 + 1 :
                                             I2d1670c45bd1cc15172a12175f7fb906
                                             ;

            If17c0096ce34b88007247bf4c429d5c4  <=  I2d1670c45bd1cc15172a12175f7fb906[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I768b6f55827ac49eb6ac2655e9397be1     <=
                                             Ia4c9bac1a64e1a17f7964491d880660e[SGN_MAX_SUM_WDTH] ?
                                             ~Ia4c9bac1a64e1a17f7964491d880660e + 1 :
                                             Ia4c9bac1a64e1a17f7964491d880660e
                                             ;

            Ifc2963762403a00c4f3662b2863c991e  <=  Ia4c9bac1a64e1a17f7964491d880660e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic66f737fe60c55d4c10e5d72b307a061     <=
                                             Ibff15c9092ff0ab60ccfd9528d5477bf[SGN_MAX_SUM_WDTH] ?
                                             ~Ibff15c9092ff0ab60ccfd9528d5477bf + 1 :
                                             Ibff15c9092ff0ab60ccfd9528d5477bf
                                             ;

            I5fdd8e1550feaecd81b82069fe73ed7e  <=  Ibff15c9092ff0ab60ccfd9528d5477bf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5653779f15c6c9b0f3b26927c48d6234     <=
                                             Iac2e396e7f63a651c52c6aa372419808[SGN_MAX_SUM_WDTH] ?
                                             ~Iac2e396e7f63a651c52c6aa372419808 + 1 :
                                             Iac2e396e7f63a651c52c6aa372419808
                                             ;

            I85654bd3a07b4329aba17d8b27777f4e  <=  Iac2e396e7f63a651c52c6aa372419808[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iac550729fc437fd67151fab57134ec88     <=
                                             Ice856d92219493a98683a6e36f6a81f6[SGN_MAX_SUM_WDTH] ?
                                             ~Ice856d92219493a98683a6e36f6a81f6 + 1 :
                                             Ice856d92219493a98683a6e36f6a81f6
                                             ;

            Ibf2a253afde05c905d0b2404c5a808a0  <=  Ice856d92219493a98683a6e36f6a81f6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I853b03c5826eedc3c67a2fae7a640212     <=
                                             I5e784ab32ea84026fa63ce432c6f604f[SGN_MAX_SUM_WDTH] ?
                                             ~I5e784ab32ea84026fa63ce432c6f604f + 1 :
                                             I5e784ab32ea84026fa63ce432c6f604f
                                             ;

            I3ade5535a79ce83857481ac771cd8618  <=  I5e784ab32ea84026fa63ce432c6f604f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If46a6b47c1c52243cc0bc92d1edb594f     <=
                                             I32251a5b768526c3599f145a3eed1949[SGN_MAX_SUM_WDTH] ?
                                             ~I32251a5b768526c3599f145a3eed1949 + 1 :
                                             I32251a5b768526c3599f145a3eed1949
                                             ;

            I221524a69e18854f029cad30e8f94e8a  <=  I32251a5b768526c3599f145a3eed1949[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I75b36a9b429cd657afc8151b9613aca6     <=
                                             I6357b0d86d75dc1018fa50248f3e2deb[SGN_MAX_SUM_WDTH] ?
                                             ~I6357b0d86d75dc1018fa50248f3e2deb + 1 :
                                             I6357b0d86d75dc1018fa50248f3e2deb
                                             ;

            Ied764ee7730ad129b6f62837ef50774a  <=  I6357b0d86d75dc1018fa50248f3e2deb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ife682dd9f677da4d27294fb61b141948     <=
                                             I8a50948f1b1f5589972c137e91e4eee0[SGN_MAX_SUM_WDTH] ?
                                             ~I8a50948f1b1f5589972c137e91e4eee0 + 1 :
                                             I8a50948f1b1f5589972c137e91e4eee0
                                             ;

            Ic98f33c6a4613534bcc9b6bc4b4f2d17  <=  I8a50948f1b1f5589972c137e91e4eee0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2b6177a9c586b274b68b25584e6df2c     <=
                                             Icce2cc29f7ad95af1a9605954033fce0[SGN_MAX_SUM_WDTH] ?
                                             ~Icce2cc29f7ad95af1a9605954033fce0 + 1 :
                                             Icce2cc29f7ad95af1a9605954033fce0
                                             ;

            I92eb6f60c14ee9eecb01718b01ea980f  <=  Icce2cc29f7ad95af1a9605954033fce0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0d23011c4381496a19cced7bf7960546     <=
                                             I276997085c2cbcdac1c886e74bc2e530[SGN_MAX_SUM_WDTH] ?
                                             ~I276997085c2cbcdac1c886e74bc2e530 + 1 :
                                             I276997085c2cbcdac1c886e74bc2e530
                                             ;

            I97e82e5f6775d1e31537b891597223bd  <=  I276997085c2cbcdac1c886e74bc2e530[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic5992d5eaeafd5dded641a7d9801e763     <=
                                             I7299d046eb7c80908def7e3ec9665c88[SGN_MAX_SUM_WDTH] ?
                                             ~I7299d046eb7c80908def7e3ec9665c88 + 1 :
                                             I7299d046eb7c80908def7e3ec9665c88
                                             ;

            Iba1c0ebd9cefeb0dd7f690bdbbbfec58  <=  I7299d046eb7c80908def7e3ec9665c88[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic9e7fe68b9045c6c9eb86185b5f5872e     <=
                                             I8f993e6b8e7313dfb4323ebf4ccdb640[SGN_MAX_SUM_WDTH] ?
                                             ~I8f993e6b8e7313dfb4323ebf4ccdb640 + 1 :
                                             I8f993e6b8e7313dfb4323ebf4ccdb640
                                             ;

            I235c3a9fd3e8ea1cee762c10bc8e2c53  <=  I8f993e6b8e7313dfb4323ebf4ccdb640[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I51ad746720b5e6e09ab50f0283552f1a     <=
                                             I2b75fcd754488677526db195256ddc06[SGN_MAX_SUM_WDTH] ?
                                             ~I2b75fcd754488677526db195256ddc06 + 1 :
                                             I2b75fcd754488677526db195256ddc06
                                             ;

            Idd474d80b50992537d6f527faf279800  <=  I2b75fcd754488677526db195256ddc06[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0c8964888a1315507f5d71959dd24cf0     <=
                                             Ide04235316ff1098fd97e125d76797c2[SGN_MAX_SUM_WDTH] ?
                                             ~Ide04235316ff1098fd97e125d76797c2 + 1 :
                                             Ide04235316ff1098fd97e125d76797c2
                                             ;

            I88a89b2d938552458dab9bc34728959b  <=  Ide04235316ff1098fd97e125d76797c2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id4d4f814a0bb3418cbf70c306acf048f     <=
                                             I39755c95fddbe19ae343164be78b0fff[SGN_MAX_SUM_WDTH] ?
                                             ~I39755c95fddbe19ae343164be78b0fff + 1 :
                                             I39755c95fddbe19ae343164be78b0fff
                                             ;

            Ib105151d91678f81978495ff94b1e651  <=  I39755c95fddbe19ae343164be78b0fff[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic91bd7b4bd148e526ca21d4a5ba87be9     <=
                                             I37d4177c1ea3ac376d3906e49a4a3224[SGN_MAX_SUM_WDTH] ?
                                             ~I37d4177c1ea3ac376d3906e49a4a3224 + 1 :
                                             I37d4177c1ea3ac376d3906e49a4a3224
                                             ;

            I4edd64d1f1da865b1eb886e22726a033  <=  I37d4177c1ea3ac376d3906e49a4a3224[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7959dddc32f0f181b3ba39149afe1016     <=
                                             Ifd04130d9f32af7f7debe20de6b6fa57[SGN_MAX_SUM_WDTH] ?
                                             ~Ifd04130d9f32af7f7debe20de6b6fa57 + 1 :
                                             Ifd04130d9f32af7f7debe20de6b6fa57
                                             ;

            Ia7c9c24f8e993526e76c6915e56908c4  <=  Ifd04130d9f32af7f7debe20de6b6fa57[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I087263600b5f38be072a4f1db787aea7     <=
                                             I7ee40f0225ba9aad10df1dec7a0f25fd[SGN_MAX_SUM_WDTH] ?
                                             ~I7ee40f0225ba9aad10df1dec7a0f25fd + 1 :
                                             I7ee40f0225ba9aad10df1dec7a0f25fd
                                             ;

            Ib0dadebad37d9ea9d01350054872863c  <=  I7ee40f0225ba9aad10df1dec7a0f25fd[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I78d17a56de5cbe08191ef23b9731c485     <=
                                             Ic780d894a72f9111937594d50a9ce311[SGN_MAX_SUM_WDTH] ?
                                             ~Ic780d894a72f9111937594d50a9ce311 + 1 :
                                             Ic780d894a72f9111937594d50a9ce311
                                             ;

            I76fd9005abd511c3c5bf6c77de8bf2f3  <=  Ic780d894a72f9111937594d50a9ce311[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I82f713a43596df3b935d6da6f8041dc2     <=
                                             I36feeea802ed7e4122a43a71d976b7d2[SGN_MAX_SUM_WDTH] ?
                                             ~I36feeea802ed7e4122a43a71d976b7d2 + 1 :
                                             I36feeea802ed7e4122a43a71d976b7d2
                                             ;

            Ic124975d36a292816146a2fe61ab3ab9  <=  I36feeea802ed7e4122a43a71d976b7d2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I422987396853a6a39dabb6e7ddbf91fb     <=
                                             I698319d790c8eb982fb1b113437d93be[SGN_MAX_SUM_WDTH] ?
                                             ~I698319d790c8eb982fb1b113437d93be + 1 :
                                             I698319d790c8eb982fb1b113437d93be
                                             ;

            I70a4926e9e6a05fa9ee51a26988862fe  <=  I698319d790c8eb982fb1b113437d93be[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibb6556671e104141dd33188ea5fc024d     <=
                                             I69c4cabd4c61dd816fbc44ae02f3d8ab[SGN_MAX_SUM_WDTH] ?
                                             ~I69c4cabd4c61dd816fbc44ae02f3d8ab + 1 :
                                             I69c4cabd4c61dd816fbc44ae02f3d8ab
                                             ;

            Idc5e98f6958786ccf95d39b922b42ea9  <=  I69c4cabd4c61dd816fbc44ae02f3d8ab[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie42ce76076a2a5e887e0112086012da6     <=
                                             Id504dcc780b333a51585556c4b58c610[SGN_MAX_SUM_WDTH] ?
                                             ~Id504dcc780b333a51585556c4b58c610 + 1 :
                                             Id504dcc780b333a51585556c4b58c610
                                             ;

            I8879df010bbdf6e5fc9370e2fb3289b4  <=  Id504dcc780b333a51585556c4b58c610[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4aea430599b9c0702b3bebd5960b5c91     <=
                                             I0c8aff3de7ee8ede0d8755cb4aebe427[SGN_MAX_SUM_WDTH] ?
                                             ~I0c8aff3de7ee8ede0d8755cb4aebe427 + 1 :
                                             I0c8aff3de7ee8ede0d8755cb4aebe427
                                             ;

            I94a9de743d5bedbea3876de954f479bd  <=  I0c8aff3de7ee8ede0d8755cb4aebe427[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icbe11a3970136e485eee1bc5053e7273     <=
                                             I1898ec6433c0e994bf697eb3b7ae5eb3[SGN_MAX_SUM_WDTH] ?
                                             ~I1898ec6433c0e994bf697eb3b7ae5eb3 + 1 :
                                             I1898ec6433c0e994bf697eb3b7ae5eb3
                                             ;

            I17c9d8f658dd6b2916b645d103f4702a  <=  I1898ec6433c0e994bf697eb3b7ae5eb3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0a7f1ea1719c1f5ff104445a4130a5a8     <=
                                             I41b391dce086564a0de53aa3f82b510a[SGN_MAX_SUM_WDTH] ?
                                             ~I41b391dce086564a0de53aa3f82b510a + 1 :
                                             I41b391dce086564a0de53aa3f82b510a
                                             ;

            I384e50fa8daa639124f083dda56fac00  <=  I41b391dce086564a0de53aa3f82b510a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1802d759f26dd919bc315bfd4156238d     <=
                                             I90c35450751e2a9607e95ebe3115c51c[SGN_MAX_SUM_WDTH] ?
                                             ~I90c35450751e2a9607e95ebe3115c51c + 1 :
                                             I90c35450751e2a9607e95ebe3115c51c
                                             ;

            Ie165d0729542c81ca89f45d15e0afd3d  <=  I90c35450751e2a9607e95ebe3115c51c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2148493e253783fad70f4f2807b83008     <=
                                             I02be13e15f91f4957ba7086ee96c1ca7[SGN_MAX_SUM_WDTH] ?
                                             ~I02be13e15f91f4957ba7086ee96c1ca7 + 1 :
                                             I02be13e15f91f4957ba7086ee96c1ca7
                                             ;

            Ie8e29053f122a9247b0dec291c6ef4f3  <=  I02be13e15f91f4957ba7086ee96c1ca7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I39e7f78d33aa7f50264908d2efe23634     <=
                                             I02cc4624a6245c0c54b079dfe50420d4[SGN_MAX_SUM_WDTH] ?
                                             ~I02cc4624a6245c0c54b079dfe50420d4 + 1 :
                                             I02cc4624a6245c0c54b079dfe50420d4
                                             ;

            I453dd7d7c0a2f003f0b67e909630d641  <=  I02cc4624a6245c0c54b079dfe50420d4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I844be5874def16af98de935019f35fe8     <=
                                             Ib0942c283a523d31d5d11a51f01fa016[SGN_MAX_SUM_WDTH] ?
                                             ~Ib0942c283a523d31d5d11a51f01fa016 + 1 :
                                             Ib0942c283a523d31d5d11a51f01fa016
                                             ;

            I5707d30ca29842b6a96cfaeb44ac6668  <=  Ib0942c283a523d31d5d11a51f01fa016[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iee5172ba70a6e368b4903f9ff1d93471     <=
                                             I93ad63d6294ac100b7027b8190f15387[SGN_MAX_SUM_WDTH] ?
                                             ~I93ad63d6294ac100b7027b8190f15387 + 1 :
                                             I93ad63d6294ac100b7027b8190f15387
                                             ;

            I3fbd40faa4c3b78b547b8348c466fd1f  <=  I93ad63d6294ac100b7027b8190f15387[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1f34b473283291e0970879465c005e2f     <=
                                             I8b92187b5833150d05b4b09f74441a20[SGN_MAX_SUM_WDTH] ?
                                             ~I8b92187b5833150d05b4b09f74441a20 + 1 :
                                             I8b92187b5833150d05b4b09f74441a20
                                             ;

            I9a403c511fe2d44472ab319a9477199c  <=  I8b92187b5833150d05b4b09f74441a20[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie1e0b5120737a7f4bf845618ccd22239     <=
                                             I02846f27754a2fbc493cc1d0848b9090[SGN_MAX_SUM_WDTH] ?
                                             ~I02846f27754a2fbc493cc1d0848b9090 + 1 :
                                             I02846f27754a2fbc493cc1d0848b9090
                                             ;

            I9db50007841762c9a10f6b7e9d40f858  <=  I02846f27754a2fbc493cc1d0848b9090[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8abec3020ee5358f8768e5595e9992b4     <=
                                             Iea2573c99c098c5fe2ee97a9c1aae44d[SGN_MAX_SUM_WDTH] ?
                                             ~Iea2573c99c098c5fe2ee97a9c1aae44d + 1 :
                                             Iea2573c99c098c5fe2ee97a9c1aae44d
                                             ;

            I89c5af1a6176cefa1f77ee69996473cb  <=  Iea2573c99c098c5fe2ee97a9c1aae44d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6fe683073211a484cb6e3c416b365d9f     <=
                                             I8c250d6e46e2d8a7f2f77035526c1f8e[SGN_MAX_SUM_WDTH] ?
                                             ~I8c250d6e46e2d8a7f2f77035526c1f8e + 1 :
                                             I8c250d6e46e2d8a7f2f77035526c1f8e
                                             ;

            I5ede62333e0f7ddc5446b653ba9a2382  <=  I8c250d6e46e2d8a7f2f77035526c1f8e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id7d764da58ade36853e8a45b5ee19dc3     <=
                                             Ic968e5570985a076b609845c9968110c[SGN_MAX_SUM_WDTH] ?
                                             ~Ic968e5570985a076b609845c9968110c + 1 :
                                             Ic968e5570985a076b609845c9968110c
                                             ;

            I69d82ab774d52c219509e993e7cc4deb  <=  Ic968e5570985a076b609845c9968110c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3cee2fdf353643deac7d6bca20c8fb52     <=
                                             Iccd14e61a9147bf5aefe4a196485ef03[SGN_MAX_SUM_WDTH] ?
                                             ~Iccd14e61a9147bf5aefe4a196485ef03 + 1 :
                                             Iccd14e61a9147bf5aefe4a196485ef03
                                             ;

            I0eaa22f5eca8f33dd254fe241017a098  <=  Iccd14e61a9147bf5aefe4a196485ef03[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie9b8f8f0434fe3783c3d8f68fef30e50     <=
                                             I4e09b4d678ce7239bad645b57535df20[SGN_MAX_SUM_WDTH] ?
                                             ~I4e09b4d678ce7239bad645b57535df20 + 1 :
                                             I4e09b4d678ce7239bad645b57535df20
                                             ;

            I570c036d0237c53bb069c52d621e539e  <=  I4e09b4d678ce7239bad645b57535df20[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I68cba8ad7742cbb34d0b1fb16be4a58a     <=
                                             I6bdb1743d21a19cf2ce13b056271d1b0[SGN_MAX_SUM_WDTH] ?
                                             ~I6bdb1743d21a19cf2ce13b056271d1b0 + 1 :
                                             I6bdb1743d21a19cf2ce13b056271d1b0
                                             ;

            I9d7614d286377329eb3999213889b707  <=  I6bdb1743d21a19cf2ce13b056271d1b0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idcea56657d40e0fdf9a1c2d920938fd6     <=
                                             I6259bbd85d21c216632a71648eddae35[SGN_MAX_SUM_WDTH] ?
                                             ~I6259bbd85d21c216632a71648eddae35 + 1 :
                                             I6259bbd85d21c216632a71648eddae35
                                             ;

            I3eab1582cc42db0ac7739386cce2a712  <=  I6259bbd85d21c216632a71648eddae35[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic549ffab8f0ce161a177faa2ffd1326d     <=
                                             I8a654b2420f09bd4b14bc5f5faa7d40d[SGN_MAX_SUM_WDTH] ?
                                             ~I8a654b2420f09bd4b14bc5f5faa7d40d + 1 :
                                             I8a654b2420f09bd4b14bc5f5faa7d40d
                                             ;

            Ie4827dc0983c1a63053c08de6e36d375  <=  I8a654b2420f09bd4b14bc5f5faa7d40d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4d463d500f93f74b2724972ec1d62439     <=
                                             I50d163f8fe5bbb86e3843bea768f049e[SGN_MAX_SUM_WDTH] ?
                                             ~I50d163f8fe5bbb86e3843bea768f049e + 1 :
                                             I50d163f8fe5bbb86e3843bea768f049e
                                             ;

            I2eed3d32a27d51036e17c4a21382b4c1  <=  I50d163f8fe5bbb86e3843bea768f049e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iba2f362e263953331649c726afa9c481     <=
                                             Ic3e2b4869f7ac3d189713dcc40a1fb30[SGN_MAX_SUM_WDTH] ?
                                             ~Ic3e2b4869f7ac3d189713dcc40a1fb30 + 1 :
                                             Ic3e2b4869f7ac3d189713dcc40a1fb30
                                             ;

            Ie039ab562e9cf90289047b5425186123  <=  Ic3e2b4869f7ac3d189713dcc40a1fb30[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6a053d931fb030e03d4882856d3bda75     <=
                                             I3d8f79c5f5af5112dc5f7fdfaf0a2434[SGN_MAX_SUM_WDTH] ?
                                             ~I3d8f79c5f5af5112dc5f7fdfaf0a2434 + 1 :
                                             I3d8f79c5f5af5112dc5f7fdfaf0a2434
                                             ;

            Iefbdf686d9452a62cb99cf023a4d9fe7  <=  I3d8f79c5f5af5112dc5f7fdfaf0a2434[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I27ede93004e0c240efaa56cc8c570910     <=
                                             I0544d6bafecefee496a6227c698a4d1a[SGN_MAX_SUM_WDTH] ?
                                             ~I0544d6bafecefee496a6227c698a4d1a + 1 :
                                             I0544d6bafecefee496a6227c698a4d1a
                                             ;

            Idc5dd6caa4ed17a63746d30d381a944e  <=  I0544d6bafecefee496a6227c698a4d1a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I61a11c1711ca10eefea3438722b40bff     <=
                                             I6672e8613ad03882a4b7f4141a56d535[SGN_MAX_SUM_WDTH] ?
                                             ~I6672e8613ad03882a4b7f4141a56d535 + 1 :
                                             I6672e8613ad03882a4b7f4141a56d535
                                             ;

            I17086dc5193aa55e5c6f56ecd365cc00  <=  I6672e8613ad03882a4b7f4141a56d535[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia7924c88692cfddf24fb1eff66eacb7e     <=
                                             I1542f0db2447a8b733077daebe1d2321[SGN_MAX_SUM_WDTH] ?
                                             ~I1542f0db2447a8b733077daebe1d2321 + 1 :
                                             I1542f0db2447a8b733077daebe1d2321
                                             ;

            Ib2fe0f68044c11f879e512a200f8099e  <=  I1542f0db2447a8b733077daebe1d2321[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibcfd01e622f7f5a5156dd9b335b4e5e0     <=
                                             I3038115e5ee2b90df4a7ad7e25d5337d[SGN_MAX_SUM_WDTH] ?
                                             ~I3038115e5ee2b90df4a7ad7e25d5337d + 1 :
                                             I3038115e5ee2b90df4a7ad7e25d5337d
                                             ;

            I768720af835b02a8dab376ef23d17a15  <=  I3038115e5ee2b90df4a7ad7e25d5337d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7f6f418ea51b4298da8758bda3f6a21b     <=
                                             I758ce2910b56968ca8ebc74c19f2cb47[SGN_MAX_SUM_WDTH] ?
                                             ~I758ce2910b56968ca8ebc74c19f2cb47 + 1 :
                                             I758ce2910b56968ca8ebc74c19f2cb47
                                             ;

            I1d98943b01a6a2d8c4db18b98dd62f5c  <=  I758ce2910b56968ca8ebc74c19f2cb47[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7185da8937449e23abdd0f39a4b3ed7d     <=
                                             Ifd3191045c45b2f46fbbb63b1766e9fb[SGN_MAX_SUM_WDTH] ?
                                             ~Ifd3191045c45b2f46fbbb63b1766e9fb + 1 :
                                             Ifd3191045c45b2f46fbbb63b1766e9fb
                                             ;

            Id3b089fb6edd5bcfdbca142fddd5ff89  <=  Ifd3191045c45b2f46fbbb63b1766e9fb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idc3e3ffa31d9b76c7cf9358a5b2e65d7     <=
                                             I5a15f4c8b810f7234d421967f4d926c6[SGN_MAX_SUM_WDTH] ?
                                             ~I5a15f4c8b810f7234d421967f4d926c6 + 1 :
                                             I5a15f4c8b810f7234d421967f4d926c6
                                             ;

            I5196382b75d16892d550f17893de15ec  <=  I5a15f4c8b810f7234d421967f4d926c6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I31fe8c887c4aff7c69336676cd31aaa1     <=
                                             I6f82614fc25bf322e359b929caa86025[SGN_MAX_SUM_WDTH] ?
                                             ~I6f82614fc25bf322e359b929caa86025 + 1 :
                                             I6f82614fc25bf322e359b929caa86025
                                             ;

            I6387919f2426c283e2d70e471cda54a6  <=  I6f82614fc25bf322e359b929caa86025[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I59684d5fe6bbb4b54ac097bd25fceef5     <=
                                             I4dcffaa8c903a955a4c4b5197cd2d728[SGN_MAX_SUM_WDTH] ?
                                             ~I4dcffaa8c903a955a4c4b5197cd2d728 + 1 :
                                             I4dcffaa8c903a955a4c4b5197cd2d728
                                             ;

            I3b84dad6d0dd8730312b3e20c6d5a2a8  <=  I4dcffaa8c903a955a4c4b5197cd2d728[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I86a7cd69148f9590ce91d0aa270d6c54     <=
                                             I71dbc37567c4c703f28c39b97c44d1dc[SGN_MAX_SUM_WDTH] ?
                                             ~I71dbc37567c4c703f28c39b97c44d1dc + 1 :
                                             I71dbc37567c4c703f28c39b97c44d1dc
                                             ;

            I2a4bbedf880a9a7b4e1bf946f9f96c0e  <=  I71dbc37567c4c703f28c39b97c44d1dc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iabce1ccdd968980f622f0e137b159d11     <=
                                             I224678d6b3b2a1ed8f2368d7035134d4[SGN_MAX_SUM_WDTH] ?
                                             ~I224678d6b3b2a1ed8f2368d7035134d4 + 1 :
                                             I224678d6b3b2a1ed8f2368d7035134d4
                                             ;

            I49d35ec6369de10afb15be8e0cf135c3  <=  I224678d6b3b2a1ed8f2368d7035134d4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iff02977d7b4c733cca1794246f630931     <=
                                             I6942bdfb9c73af7b24e91f3cc2c40443[SGN_MAX_SUM_WDTH] ?
                                             ~I6942bdfb9c73af7b24e91f3cc2c40443 + 1 :
                                             I6942bdfb9c73af7b24e91f3cc2c40443
                                             ;

            Ic3ba4531855366e9a060cec1c7694844  <=  I6942bdfb9c73af7b24e91f3cc2c40443[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9026c904e5ead7ff2994c4f781d61466     <=
                                             I8eae50dae3f5eadae891e7875180bd47[SGN_MAX_SUM_WDTH] ?
                                             ~I8eae50dae3f5eadae891e7875180bd47 + 1 :
                                             I8eae50dae3f5eadae891e7875180bd47
                                             ;

            I4dbabfd592b74aef93b819163130ef5e  <=  I8eae50dae3f5eadae891e7875180bd47[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I99d7489ba87c629c6dd9702a9bbfd3c8     <=
                                             I5ab8c899cb9e33273d3e5758757dbdfd[SGN_MAX_SUM_WDTH] ?
                                             ~I5ab8c899cb9e33273d3e5758757dbdfd + 1 :
                                             I5ab8c899cb9e33273d3e5758757dbdfd
                                             ;

            I9ece87047aec25abc02a5eea72f0e647  <=  I5ab8c899cb9e33273d3e5758757dbdfd[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifaf191e0d00ba6da7019c2efcf08e1d9     <=
                                             I23890d77a1b1c3fea977146599cee178[SGN_MAX_SUM_WDTH] ?
                                             ~I23890d77a1b1c3fea977146599cee178 + 1 :
                                             I23890d77a1b1c3fea977146599cee178
                                             ;

            I3ed6426fbdba8aaf1c948cca7442b3a6  <=  I23890d77a1b1c3fea977146599cee178[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4c295991fb08c90862a2f3ba6489000a     <=
                                             Ib311a6a7fc40711d6920e3c43b31c5c2[SGN_MAX_SUM_WDTH] ?
                                             ~Ib311a6a7fc40711d6920e3c43b31c5c2 + 1 :
                                             Ib311a6a7fc40711d6920e3c43b31c5c2
                                             ;

            I24075f37c6bbd90c83370de1a2e58af2  <=  Ib311a6a7fc40711d6920e3c43b31c5c2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iee61d179da125934298400256788cbb8     <=
                                             Ifc3cc051690f3d687caa05e26dde6d93[SGN_MAX_SUM_WDTH] ?
                                             ~Ifc3cc051690f3d687caa05e26dde6d93 + 1 :
                                             Ifc3cc051690f3d687caa05e26dde6d93
                                             ;

            I3175159add7b814df637c2db8feb43f6  <=  Ifc3cc051690f3d687caa05e26dde6d93[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If87c84440426fb24070372dc1d4bf315     <=
                                             Ida60773a931859ee7e5e2db24b9bb72c[SGN_MAX_SUM_WDTH] ?
                                             ~Ida60773a931859ee7e5e2db24b9bb72c + 1 :
                                             Ida60773a931859ee7e5e2db24b9bb72c
                                             ;

            I0a569f6536789efb7ad2377c11842830  <=  Ida60773a931859ee7e5e2db24b9bb72c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib9259a807b31c1b7a528d336bfc403ee     <=
                                             Id5e39679bbe2407407a53366e77aed13[SGN_MAX_SUM_WDTH] ?
                                             ~Id5e39679bbe2407407a53366e77aed13 + 1 :
                                             Id5e39679bbe2407407a53366e77aed13
                                             ;

            Iae6ed7748692f2edf1aa9d73380075f0  <=  Id5e39679bbe2407407a53366e77aed13[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I411c4d909b2a571e685cd703245516d7     <=
                                             Ie3eab29a9004627e296a198708459545[SGN_MAX_SUM_WDTH] ?
                                             ~Ie3eab29a9004627e296a198708459545 + 1 :
                                             Ie3eab29a9004627e296a198708459545
                                             ;

            Ib4ae1cedd09d72c235765a6cd7e91366  <=  Ie3eab29a9004627e296a198708459545[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If8425453cca8fc8623cb85375c4b8a1d     <=
                                             I86c0872f8ce743bb3fa7b3fca2dea33b[SGN_MAX_SUM_WDTH] ?
                                             ~I86c0872f8ce743bb3fa7b3fca2dea33b + 1 :
                                             I86c0872f8ce743bb3fa7b3fca2dea33b
                                             ;

            Ie2d946edaddd3c87f328e861f3e72c0a  <=  I86c0872f8ce743bb3fa7b3fca2dea33b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I654b497f62df75fa283127b5de29b1ad     <=
                                             Id1aa022173e0fa45a3f26b4d31e113a3[SGN_MAX_SUM_WDTH] ?
                                             ~Id1aa022173e0fa45a3f26b4d31e113a3 + 1 :
                                             Id1aa022173e0fa45a3f26b4d31e113a3
                                             ;

            Id6b508145cd21ba088ab8fda34577c35  <=  Id1aa022173e0fa45a3f26b4d31e113a3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2768519342f7b8a1ee40c1d5ac502b66     <=
                                             I0bfd4314a81f9f0930e549a09ef4c68f[SGN_MAX_SUM_WDTH] ?
                                             ~I0bfd4314a81f9f0930e549a09ef4c68f + 1 :
                                             I0bfd4314a81f9f0930e549a09ef4c68f
                                             ;

            Ifa6e3541f5e12bf9677ffc51d0392749  <=  I0bfd4314a81f9f0930e549a09ef4c68f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8e354c1c5ba44fe5430887248ce0c43b     <=
                                             I2e90a66f2eedee35927bcb8c5ff26fbe[SGN_MAX_SUM_WDTH] ?
                                             ~I2e90a66f2eedee35927bcb8c5ff26fbe + 1 :
                                             I2e90a66f2eedee35927bcb8c5ff26fbe
                                             ;

            I21e72a7e5870151c3247d15121e5fb4f  <=  I2e90a66f2eedee35927bcb8c5ff26fbe[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8970d8a8aea29913e8696c14c153d16e     <=
                                             I9d6828434155b5672b44a1172ae9b6eb[SGN_MAX_SUM_WDTH] ?
                                             ~I9d6828434155b5672b44a1172ae9b6eb + 1 :
                                             I9d6828434155b5672b44a1172ae9b6eb
                                             ;

            Iba283e99a57d0a3b78ad2e309c316b65  <=  I9d6828434155b5672b44a1172ae9b6eb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3555c6e2fd480a6be11549bf95a9b0b1     <=
                                             I0483abcf888b35d85e8a62c901b6021b[SGN_MAX_SUM_WDTH] ?
                                             ~I0483abcf888b35d85e8a62c901b6021b + 1 :
                                             I0483abcf888b35d85e8a62c901b6021b
                                             ;

            Ifba3e46933049cb093d2c1809f3a8a3e  <=  I0483abcf888b35d85e8a62c901b6021b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8d5600a352e8ba4756f917f912fda6dd     <=
                                             I8f6514c2e33675cd94350a1e1b0b5f80[SGN_MAX_SUM_WDTH] ?
                                             ~I8f6514c2e33675cd94350a1e1b0b5f80 + 1 :
                                             I8f6514c2e33675cd94350a1e1b0b5f80
                                             ;

            I4af3e2bf2ebc913ac902b48da672c5b6  <=  I8f6514c2e33675cd94350a1e1b0b5f80[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7e99d73c95e7ae5c3fe07a3c60ef52eb     <=
                                             I23d3830f616b3be90cd63e45b606fc2e[SGN_MAX_SUM_WDTH] ?
                                             ~I23d3830f616b3be90cd63e45b606fc2e + 1 :
                                             I23d3830f616b3be90cd63e45b606fc2e
                                             ;

            Ifbadefd3a7ab50719a703400ddd742c6  <=  I23d3830f616b3be90cd63e45b606fc2e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I831633aebe5c6a52b98d630205376f3a     <=
                                             I106ef13f4b977bc5b978b5977cc06eb7[SGN_MAX_SUM_WDTH] ?
                                             ~I106ef13f4b977bc5b978b5977cc06eb7 + 1 :
                                             I106ef13f4b977bc5b978b5977cc06eb7
                                             ;

            If2042aede3390bd208a281f0380c95a4  <=  I106ef13f4b977bc5b978b5977cc06eb7[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I82e35482de74223be0d2558334ac2dfb     <=
                                             I3fdcbddec1b193cc85d20d4796aef72b[SGN_MAX_SUM_WDTH] ?
                                             ~I3fdcbddec1b193cc85d20d4796aef72b + 1 :
                                             I3fdcbddec1b193cc85d20d4796aef72b
                                             ;

            I19b73c5c93a71e90f620572f23f0e6d2  <=  I3fdcbddec1b193cc85d20d4796aef72b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iae2a6f9649ef1bb193e4f0ab5ecbc3e3     <=
                                             I3956ec3a4f9d8ea94a760b5c6388f2b0[SGN_MAX_SUM_WDTH] ?
                                             ~I3956ec3a4f9d8ea94a760b5c6388f2b0 + 1 :
                                             I3956ec3a4f9d8ea94a760b5c6388f2b0
                                             ;

            I4b99891bed4f5c149cd4a5b4f1dde0f0  <=  I3956ec3a4f9d8ea94a760b5c6388f2b0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie8eca65d791ad2f6e8f4ed244f22ae3d     <=
                                             I5541cea9c0da962da2b7d9154c66de98[SGN_MAX_SUM_WDTH] ?
                                             ~I5541cea9c0da962da2b7d9154c66de98 + 1 :
                                             I5541cea9c0da962da2b7d9154c66de98
                                             ;

            I3472ee8c06644490252e606b62bf9bd5  <=  I5541cea9c0da962da2b7d9154c66de98[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic24146b01094df9b9ccd455a791f239d     <=
                                             I0c1edbaa3c2f47d66034fccd799b5387[SGN_MAX_SUM_WDTH] ?
                                             ~I0c1edbaa3c2f47d66034fccd799b5387 + 1 :
                                             I0c1edbaa3c2f47d66034fccd799b5387
                                             ;

            Idb1efe99b5d7fd567a7f82cfd52f7eb8  <=  I0c1edbaa3c2f47d66034fccd799b5387[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1c9031fd54ff9417d44c9fb17dc1fc63     <=
                                             Ia6eb0c9c2e6c3a440defef2c3879de88[SGN_MAX_SUM_WDTH] ?
                                             ~Ia6eb0c9c2e6c3a440defef2c3879de88 + 1 :
                                             Ia6eb0c9c2e6c3a440defef2c3879de88
                                             ;

            I24f82a3f2c0e8df486fe495dd95cf8bc  <=  Ia6eb0c9c2e6c3a440defef2c3879de88[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idefa20487bc5ba6daff03e6b327d76c6     <=
                                             Ifcef7363a6ecbb3b3248cb65bb6b0d17[SGN_MAX_SUM_WDTH] ?
                                             ~Ifcef7363a6ecbb3b3248cb65bb6b0d17 + 1 :
                                             Ifcef7363a6ecbb3b3248cb65bb6b0d17
                                             ;

            I83ecf12f3b38fc14c3b75e47b71ecc09  <=  Ifcef7363a6ecbb3b3248cb65bb6b0d17[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6f984fd9ea27b40ab3afeac8afd29ade     <=
                                             I5e36ed7643bf47aef14bd47a835e1a01[SGN_MAX_SUM_WDTH] ?
                                             ~I5e36ed7643bf47aef14bd47a835e1a01 + 1 :
                                             I5e36ed7643bf47aef14bd47a835e1a01
                                             ;

            I74cbc0ec3bb682e0f927890eef8d7a58  <=  I5e36ed7643bf47aef14bd47a835e1a01[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0be92debced4961df5f461fe81e80bf1     <=
                                             Idc662c9332f4a6cafe820ad2bc0d16e1[SGN_MAX_SUM_WDTH] ?
                                             ~Idc662c9332f4a6cafe820ad2bc0d16e1 + 1 :
                                             Idc662c9332f4a6cafe820ad2bc0d16e1
                                             ;

            I989dda9add29306d7b3c0f376822763a  <=  Idc662c9332f4a6cafe820ad2bc0d16e1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia7bdaba4c6601b7146498aea6c9a3e07     <=
                                             Id51e465dc2adba5eedf6ad37d0a25aa3[SGN_MAX_SUM_WDTH] ?
                                             ~Id51e465dc2adba5eedf6ad37d0a25aa3 + 1 :
                                             Id51e465dc2adba5eedf6ad37d0a25aa3
                                             ;

            Ibc929201e2eeb3e61cc8f0acbade497a  <=  Id51e465dc2adba5eedf6ad37d0a25aa3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id450c0a1cabe087be051fbf4158e6016     <=
                                             If0d4550f2f3884c49d1cf5a40251cd58[SGN_MAX_SUM_WDTH] ?
                                             ~If0d4550f2f3884c49d1cf5a40251cd58 + 1 :
                                             If0d4550f2f3884c49d1cf5a40251cd58
                                             ;

            Ib0dfbbbca2d3d264065f73b4241caed5  <=  If0d4550f2f3884c49d1cf5a40251cd58[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I656d0d69f6e243746b87ad67764dbc3d     <=
                                             I3af1a3cc1733db0dc42ab6214351aa99[SGN_MAX_SUM_WDTH] ?
                                             ~I3af1a3cc1733db0dc42ab6214351aa99 + 1 :
                                             I3af1a3cc1733db0dc42ab6214351aa99
                                             ;

            I339786aa60d4c71d12c65db27ac420fe  <=  I3af1a3cc1733db0dc42ab6214351aa99[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iab9d870dc1ad159bbaecb20a9b72f005     <=
                                             I022b7b4693a7e7b654b8bd85a94f0d9c[SGN_MAX_SUM_WDTH] ?
                                             ~I022b7b4693a7e7b654b8bd85a94f0d9c + 1 :
                                             I022b7b4693a7e7b654b8bd85a94f0d9c
                                             ;

            I3ade020bbdf8f954821f737439513043  <=  I022b7b4693a7e7b654b8bd85a94f0d9c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id53b60854f19e095c38f2c255dc57f29     <=
                                             I5bd1d6563b4acb8dc10d348ec0a2346a[SGN_MAX_SUM_WDTH] ?
                                             ~I5bd1d6563b4acb8dc10d348ec0a2346a + 1 :
                                             I5bd1d6563b4acb8dc10d348ec0a2346a
                                             ;

            Ia50526cd3a3174bebc5a7a0889fda661  <=  I5bd1d6563b4acb8dc10d348ec0a2346a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9ba44a2e4a8f0b61692fc69ebeb82bd     <=
                                             I17bbbddc2ace71bcd660f93fdf5e32a4[SGN_MAX_SUM_WDTH] ?
                                             ~I17bbbddc2ace71bcd660f93fdf5e32a4 + 1 :
                                             I17bbbddc2ace71bcd660f93fdf5e32a4
                                             ;

            Ie9f37dba0791359bc426a73639ce33ad  <=  I17bbbddc2ace71bcd660f93fdf5e32a4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ief95e8620a1c8ddfd6df673a3a223bd8     <=
                                             I4eb0952c6dd9719774c57b76d3cbe87a[SGN_MAX_SUM_WDTH] ?
                                             ~I4eb0952c6dd9719774c57b76d3cbe87a + 1 :
                                             I4eb0952c6dd9719774c57b76d3cbe87a
                                             ;

            I9518532a8617fc8290eb6a5e981dea94  <=  I4eb0952c6dd9719774c57b76d3cbe87a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I61519bc0aa02ed461dbb91851d0ae19e     <=
                                             I6fb63afabfeb4cc43c164e04d35a6c76[SGN_MAX_SUM_WDTH] ?
                                             ~I6fb63afabfeb4cc43c164e04d35a6c76 + 1 :
                                             I6fb63afabfeb4cc43c164e04d35a6c76
                                             ;

            If66524125bfde5aa48ac70c4e448b38f  <=  I6fb63afabfeb4cc43c164e04d35a6c76[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie0c11d584811174a66ca221baf87c36b     <=
                                             I91ba6681ef5a1092784cd98b48dc420e[SGN_MAX_SUM_WDTH] ?
                                             ~I91ba6681ef5a1092784cd98b48dc420e + 1 :
                                             I91ba6681ef5a1092784cd98b48dc420e
                                             ;

            Ic3ec6375998b05a3e48f6c5fe7b3910b  <=  I91ba6681ef5a1092784cd98b48dc420e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If10f4f45ff0fd17541735934ad20f187     <=
                                             I6eda15abfd6c1f377d25d70e35373596[SGN_MAX_SUM_WDTH] ?
                                             ~I6eda15abfd6c1f377d25d70e35373596 + 1 :
                                             I6eda15abfd6c1f377d25d70e35373596
                                             ;

            I0ac421af6e311b6005c3e02e93ff94ce  <=  I6eda15abfd6c1f377d25d70e35373596[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I445919f07a6fa8654211301a9a6126bd     <=
                                             Idf9a54c3bd991a031e09982424a8054b[SGN_MAX_SUM_WDTH] ?
                                             ~Idf9a54c3bd991a031e09982424a8054b + 1 :
                                             Idf9a54c3bd991a031e09982424a8054b
                                             ;

            Ib9db80f43718305a8a8774d8d80c86c9  <=  Idf9a54c3bd991a031e09982424a8054b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I64102b82893352549abd2e2132b19476     <=
                                             I5d7b50b4839c16d1c7010ef2c8c535c2[SGN_MAX_SUM_WDTH] ?
                                             ~I5d7b50b4839c16d1c7010ef2c8c535c2 + 1 :
                                             I5d7b50b4839c16d1c7010ef2c8c535c2
                                             ;

            I3b775b06b5d78fcd7373c966a62f44ad  <=  I5d7b50b4839c16d1c7010ef2c8c535c2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1fc1933fe891ac26f35a42a1b242d919     <=
                                             I821836ca9d1bcb5e0d12c348bb323c9a[SGN_MAX_SUM_WDTH] ?
                                             ~I821836ca9d1bcb5e0d12c348bb323c9a + 1 :
                                             I821836ca9d1bcb5e0d12c348bb323c9a
                                             ;

            If2372a5956f21f97eeb9c76281b6675e  <=  I821836ca9d1bcb5e0d12c348bb323c9a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I84dfba8bcf8ad3b85f9472fd60d607b5     <=
                                             I31f94bb809811efebb378517c2138b7f[SGN_MAX_SUM_WDTH] ?
                                             ~I31f94bb809811efebb378517c2138b7f + 1 :
                                             I31f94bb809811efebb378517c2138b7f
                                             ;

            I7b32c2b108e24750e2a24785668af3ea  <=  I31f94bb809811efebb378517c2138b7f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4302fccefe5ee13161f9ad49f9ddf43c     <=
                                             I3f203b62c645fd01c54ed43399b390e5[SGN_MAX_SUM_WDTH] ?
                                             ~I3f203b62c645fd01c54ed43399b390e5 + 1 :
                                             I3f203b62c645fd01c54ed43399b390e5
                                             ;

            I8ec99197a7d823f5745d382c10161430  <=  I3f203b62c645fd01c54ed43399b390e5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I59d7153724d3b3805af799692fbe245a     <=
                                             Ic01c569fbe524a2fe3626e4d22414e62[SGN_MAX_SUM_WDTH] ?
                                             ~Ic01c569fbe524a2fe3626e4d22414e62 + 1 :
                                             Ic01c569fbe524a2fe3626e4d22414e62
                                             ;

            Ib895fec0b3756932b85962c1d129a03e  <=  Ic01c569fbe524a2fe3626e4d22414e62[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id1650d0e39be078027493f58e9bbcbdd     <=
                                             I5a30e151cf8a2259d8cde3fa76389e78[SGN_MAX_SUM_WDTH] ?
                                             ~I5a30e151cf8a2259d8cde3fa76389e78 + 1 :
                                             I5a30e151cf8a2259d8cde3fa76389e78
                                             ;

            I76aab345d13c6678fe37a4a7133cfd7d  <=  I5a30e151cf8a2259d8cde3fa76389e78[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If40ad4aca8dbb3bf7dde8c2ff2e5b8f2     <=
                                             Ic5340f7fa98175b85f475a03156a04a6[SGN_MAX_SUM_WDTH] ?
                                             ~Ic5340f7fa98175b85f475a03156a04a6 + 1 :
                                             Ic5340f7fa98175b85f475a03156a04a6
                                             ;

            Ib4f368fa3d3ec11d9ffb2ae9a2ae6310  <=  Ic5340f7fa98175b85f475a03156a04a6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie49f173549396caeab1d13da36e37c65     <=
                                             I0b25b22531e117125c9dc82b1fb69166[SGN_MAX_SUM_WDTH] ?
                                             ~I0b25b22531e117125c9dc82b1fb69166 + 1 :
                                             I0b25b22531e117125c9dc82b1fb69166
                                             ;

            Idd0f3cfc5599481c954a2bfe69f044e5  <=  I0b25b22531e117125c9dc82b1fb69166[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3002a0e0cdf8e79bc7186a876410d106     <=
                                             Ic0c22023bce6b4e011b52acb0ac89944[SGN_MAX_SUM_WDTH] ?
                                             ~Ic0c22023bce6b4e011b52acb0ac89944 + 1 :
                                             Ic0c22023bce6b4e011b52acb0ac89944
                                             ;

            Ie624c4dad5036a25ca314b94cf3c4b95  <=  Ic0c22023bce6b4e011b52acb0ac89944[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2b50fa03f584d10e9af3be085a02a12c     <=
                                             I7f474f465227aa0e2aaa3986574ed756[SGN_MAX_SUM_WDTH] ?
                                             ~I7f474f465227aa0e2aaa3986574ed756 + 1 :
                                             I7f474f465227aa0e2aaa3986574ed756
                                             ;

            Ibf4b3caa5655cfb6663f9b7e2383bbbf  <=  I7f474f465227aa0e2aaa3986574ed756[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If473d172a7bff5aeae99245bbb72978d     <=
                                             I8869bb7415e726932972a16630d4090a[SGN_MAX_SUM_WDTH] ?
                                             ~I8869bb7415e726932972a16630d4090a + 1 :
                                             I8869bb7415e726932972a16630d4090a
                                             ;

            I049d1c09c15def12ba7bae95fc1c3d55  <=  I8869bb7415e726932972a16630d4090a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib89f7b5625995290a64bcfb143d978ca     <=
                                             Ic1afbad56abd1a486de1d72dc835ea03[SGN_MAX_SUM_WDTH] ?
                                             ~Ic1afbad56abd1a486de1d72dc835ea03 + 1 :
                                             Ic1afbad56abd1a486de1d72dc835ea03
                                             ;

            Ide06ba186ddb179b489ba6e3e209e3e8  <=  Ic1afbad56abd1a486de1d72dc835ea03[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iebe0c9b4a87d58a1c55e2ee6b01603c4     <=
                                             I0cc174ebcf049214088dd4a7dad9ebf0[SGN_MAX_SUM_WDTH] ?
                                             ~I0cc174ebcf049214088dd4a7dad9ebf0 + 1 :
                                             I0cc174ebcf049214088dd4a7dad9ebf0
                                             ;

            I1b78785ebe2e7f77a3125a6334c4dc54  <=  I0cc174ebcf049214088dd4a7dad9ebf0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I104411bb641d2445c7e1385a809bb682     <=
                                             If9a4389e51bb56f222cf06e66dcefbbb[SGN_MAX_SUM_WDTH] ?
                                             ~If9a4389e51bb56f222cf06e66dcefbbb + 1 :
                                             If9a4389e51bb56f222cf06e66dcefbbb
                                             ;

            Ie79c93f1703121713fb9401617f349a8  <=  If9a4389e51bb56f222cf06e66dcefbbb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I47dd28b4ae4f7151aff5bb271e35b716     <=
                                             Iff6098f0561da4ad6ee64dbcbf7a8b94[SGN_MAX_SUM_WDTH] ?
                                             ~Iff6098f0561da4ad6ee64dbcbf7a8b94 + 1 :
                                             Iff6098f0561da4ad6ee64dbcbf7a8b94
                                             ;

            Icf25f076eec2bf81c899c66f6cfbebc0  <=  Iff6098f0561da4ad6ee64dbcbf7a8b94[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3a27d5573b748df459b90a5a347f9d09     <=
                                             I26a679e345a21470331cd4fb2512dea0[SGN_MAX_SUM_WDTH] ?
                                             ~I26a679e345a21470331cd4fb2512dea0 + 1 :
                                             I26a679e345a21470331cd4fb2512dea0
                                             ;

            Ic5c837a0556d1cb66edbf0294d08283a  <=  I26a679e345a21470331cd4fb2512dea0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2dbef85d2b2b95af39c3a98c4e143253     <=
                                             Iec11498f4ab0492570a3454760ed5679[SGN_MAX_SUM_WDTH] ?
                                             ~Iec11498f4ab0492570a3454760ed5679 + 1 :
                                             Iec11498f4ab0492570a3454760ed5679
                                             ;

            I51ff4bda38746682e3cd4c68118c3216  <=  Iec11498f4ab0492570a3454760ed5679[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I510d39830ae7b0a857ac11baa7c144d3     <=
                                             I78154c0ca0236b79bb58bc2942b0f51b[SGN_MAX_SUM_WDTH] ?
                                             ~I78154c0ca0236b79bb58bc2942b0f51b + 1 :
                                             I78154c0ca0236b79bb58bc2942b0f51b
                                             ;

            I1c074a53e6c0f2467bcdd7c952f51670  <=  I78154c0ca0236b79bb58bc2942b0f51b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2751a94a66ea4cb44c512df4c509937f     <=
                                             I3a2c3112d5ba223b037baab170e9da79[SGN_MAX_SUM_WDTH] ?
                                             ~I3a2c3112d5ba223b037baab170e9da79 + 1 :
                                             I3a2c3112d5ba223b037baab170e9da79
                                             ;

            I37c49c5a2af240496f5a5706b0d42ea6  <=  I3a2c3112d5ba223b037baab170e9da79[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic9a003bfb70ac2da6c229fcad09246d4     <=
                                             Ia56b6d58ede63ec2b56533f0804b16df[SGN_MAX_SUM_WDTH] ?
                                             ~Ia56b6d58ede63ec2b56533f0804b16df + 1 :
                                             Ia56b6d58ede63ec2b56533f0804b16df
                                             ;

            Ia94c439131e1df5c95fc8ad3cfdba473  <=  Ia56b6d58ede63ec2b56533f0804b16df[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I34ed986182a3311a8cb005b3dccc224b     <=
                                             If8bafc8e64df4d25c725f8c577e6db43[SGN_MAX_SUM_WDTH] ?
                                             ~If8bafc8e64df4d25c725f8c577e6db43 + 1 :
                                             If8bafc8e64df4d25c725f8c577e6db43
                                             ;

            I723a6fee3b2496f23c48b3584f8bf9ce  <=  If8bafc8e64df4d25c725f8c577e6db43[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic79281755397f6099ff30c5d07d7e6de     <=
                                             Ie7452b79bbda04bebf83147d7f2ddcec[SGN_MAX_SUM_WDTH] ?
                                             ~Ie7452b79bbda04bebf83147d7f2ddcec + 1 :
                                             Ie7452b79bbda04bebf83147d7f2ddcec
                                             ;

            I648b62fa0bc2185c1756ee531e8e34de  <=  Ie7452b79bbda04bebf83147d7f2ddcec[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8d6559ccc33cbc663584923a55b928b5     <=
                                             I29a84f35944a4e286c267c60d9899c62[SGN_MAX_SUM_WDTH] ?
                                             ~I29a84f35944a4e286c267c60d9899c62 + 1 :
                                             I29a84f35944a4e286c267c60d9899c62
                                             ;

            Ife631f9a3c4c64a3d92aa9586ae75f3c  <=  I29a84f35944a4e286c267c60d9899c62[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4f0a4c241844e390318f11899a0f2c5a     <=
                                             Iae0a8cc0afb8366a7c9df146c0d08eb0[SGN_MAX_SUM_WDTH] ?
                                             ~Iae0a8cc0afb8366a7c9df146c0d08eb0 + 1 :
                                             Iae0a8cc0afb8366a7c9df146c0d08eb0
                                             ;

            Iaac1d82f0846fce1bd88ebf8e60300ac  <=  Iae0a8cc0afb8366a7c9df146c0d08eb0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I45fffa266ce3838f82d755b59216a4d6     <=
                                             I39d0497d0550115c6a2c08676c451845[SGN_MAX_SUM_WDTH] ?
                                             ~I39d0497d0550115c6a2c08676c451845 + 1 :
                                             I39d0497d0550115c6a2c08676c451845
                                             ;

            I48cd09f035f668536cd288a23010b07b  <=  I39d0497d0550115c6a2c08676c451845[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8f0e65f5db47d5460d4ec2172807a3e1     <=
                                             Ia96a79462a86a7ed9e337df66d99bf92[SGN_MAX_SUM_WDTH] ?
                                             ~Ia96a79462a86a7ed9e337df66d99bf92 + 1 :
                                             Ia96a79462a86a7ed9e337df66d99bf92
                                             ;

            I119b2e5c2fea5338244c4019884af26f  <=  Ia96a79462a86a7ed9e337df66d99bf92[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I34127c0d1af2438e13b6f4709ece80ba     <=
                                             I8ef19b31ec6d7e52e78b0c673f23ce12[SGN_MAX_SUM_WDTH] ?
                                             ~I8ef19b31ec6d7e52e78b0c673f23ce12 + 1 :
                                             I8ef19b31ec6d7e52e78b0c673f23ce12
                                             ;

            I2bd34b2fd12f12bc301fd0d5d69c0fb6  <=  I8ef19b31ec6d7e52e78b0c673f23ce12[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3a67de0e76bbf29d8c77c21865abda2f     <=
                                             I8081b1486e6def0f6ae514513c7ef4de[SGN_MAX_SUM_WDTH] ?
                                             ~I8081b1486e6def0f6ae514513c7ef4de + 1 :
                                             I8081b1486e6def0f6ae514513c7ef4de
                                             ;

            Ib715b1e0061b84ce614a30d961a83e7e  <=  I8081b1486e6def0f6ae514513c7ef4de[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic64e64aeb754249b868e14311ea19759     <=
                                             Iee5a68c2d52ef1cdd3f19b0a912603cf[SGN_MAX_SUM_WDTH] ?
                                             ~Iee5a68c2d52ef1cdd3f19b0a912603cf + 1 :
                                             Iee5a68c2d52ef1cdd3f19b0a912603cf
                                             ;

            Ief8c2838abac83370fd7ec25c06d509b  <=  Iee5a68c2d52ef1cdd3f19b0a912603cf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic4aa0dc9014c8445f8d9a7723d7263f5     <=
                                             I4b5525780a9259b57497235bd0bc69a4[SGN_MAX_SUM_WDTH] ?
                                             ~I4b5525780a9259b57497235bd0bc69a4 + 1 :
                                             I4b5525780a9259b57497235bd0bc69a4
                                             ;

            I561d79eb079915c0b1732cbddb119c2d  <=  I4b5525780a9259b57497235bd0bc69a4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I47b988d017580bdfe8f443904b1f3aac     <=
                                             Ibd65f08dbbf43d438c3a985c7b17f2e3[SGN_MAX_SUM_WDTH] ?
                                             ~Ibd65f08dbbf43d438c3a985c7b17f2e3 + 1 :
                                             Ibd65f08dbbf43d438c3a985c7b17f2e3
                                             ;

            I8bb75bf828d5ef337fa6a965808e4638  <=  Ibd65f08dbbf43d438c3a985c7b17f2e3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ica9ff13e8c3850be6c70b0b06c1d9fbf     <=
                                             Ifaa5785a3e04cd1e3be505042347fe26[SGN_MAX_SUM_WDTH] ?
                                             ~Ifaa5785a3e04cd1e3be505042347fe26 + 1 :
                                             Ifaa5785a3e04cd1e3be505042347fe26
                                             ;

            I11ba339c8250d07b497c88a39a6df1ac  <=  Ifaa5785a3e04cd1e3be505042347fe26[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If2efeb489911f295dd7722cb22ea521d     <=
                                             If0cb8cd465ff1f65de99688abd92aef2[SGN_MAX_SUM_WDTH] ?
                                             ~If0cb8cd465ff1f65de99688abd92aef2 + 1 :
                                             If0cb8cd465ff1f65de99688abd92aef2
                                             ;

            I173aa69cf52114e223ac1410d90b4bfe  <=  If0cb8cd465ff1f65de99688abd92aef2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iaa16dffcc01e41e6ff17e92bdefe3df5     <=
                                             I10ff180c115b9372f9b4b12df313372f[SGN_MAX_SUM_WDTH] ?
                                             ~I10ff180c115b9372f9b4b12df313372f + 1 :
                                             I10ff180c115b9372f9b4b12df313372f
                                             ;

            Ia4e89e99acb95f4183474b94798ca35d  <=  I10ff180c115b9372f9b4b12df313372f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie8857b9841fbd795a4192976ef7ecc25     <=
                                             I64f177202fe847d13a8a12bd80a45946[SGN_MAX_SUM_WDTH] ?
                                             ~I64f177202fe847d13a8a12bd80a45946 + 1 :
                                             I64f177202fe847d13a8a12bd80a45946
                                             ;

            If4c36727ab1c29bf78f72e8acfc00d7c  <=  I64f177202fe847d13a8a12bd80a45946[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If12aef69eea28052aa3bdb6ac31af205     <=
                                             I5df97e26d5887da447669b8d932fbdd9[SGN_MAX_SUM_WDTH] ?
                                             ~I5df97e26d5887da447669b8d932fbdd9 + 1 :
                                             I5df97e26d5887da447669b8d932fbdd9
                                             ;

            I6426943b4ab66f17c2b7b399ccc7a6a9  <=  I5df97e26d5887da447669b8d932fbdd9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0b3c6162ae2b9221738a18a29489887f     <=
                                             Ibdc07eb6a0a66e1393cb2dbd9ac77c72[SGN_MAX_SUM_WDTH] ?
                                             ~Ibdc07eb6a0a66e1393cb2dbd9ac77c72 + 1 :
                                             Ibdc07eb6a0a66e1393cb2dbd9ac77c72
                                             ;

            Iddcffa815489773b3688fd68dba18bd8  <=  Ibdc07eb6a0a66e1393cb2dbd9ac77c72[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I08211bba29e87faf4079152bcc973e7d     <=
                                             I3d353247a021629a4dd38a784eba5c1e[SGN_MAX_SUM_WDTH] ?
                                             ~I3d353247a021629a4dd38a784eba5c1e + 1 :
                                             I3d353247a021629a4dd38a784eba5c1e
                                             ;

            Id00642563679fa9a6696f8e7bbdf6576  <=  I3d353247a021629a4dd38a784eba5c1e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibff3da265f1c3f21548f5b019e1a9dc1     <=
                                             I20d77ee5328ef46daa4a54c0ae98d31a[SGN_MAX_SUM_WDTH] ?
                                             ~I20d77ee5328ef46daa4a54c0ae98d31a + 1 :
                                             I20d77ee5328ef46daa4a54c0ae98d31a
                                             ;

            Ifda1c55899cd3506853cc82b450b3936  <=  I20d77ee5328ef46daa4a54c0ae98d31a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie9fa1762d7844b0d781afdfb0771cea9     <=
                                             I8284c3a4664f99934170474b8e0e73bd[SGN_MAX_SUM_WDTH] ?
                                             ~I8284c3a4664f99934170474b8e0e73bd + 1 :
                                             I8284c3a4664f99934170474b8e0e73bd
                                             ;

            Ib5d1a7cdbcba0b654c12063d4f1768e1  <=  I8284c3a4664f99934170474b8e0e73bd[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia677d504b9f7fc2698c0345f236428ba     <=
                                             Iaeb44f2b4b78055f103df8070110b5b3[SGN_MAX_SUM_WDTH] ?
                                             ~Iaeb44f2b4b78055f103df8070110b5b3 + 1 :
                                             Iaeb44f2b4b78055f103df8070110b5b3
                                             ;

            I5e8ed024e2f2548bb375a2ecf1918a5f  <=  Iaeb44f2b4b78055f103df8070110b5b3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idebce29121c0481df83d755b60ff632c     <=
                                             Ic8242c1f7d2f582c63c3cea63d929945[SGN_MAX_SUM_WDTH] ?
                                             ~Ic8242c1f7d2f582c63c3cea63d929945 + 1 :
                                             Ic8242c1f7d2f582c63c3cea63d929945
                                             ;

            Id25deba967318f049de8163e67262f4b  <=  Ic8242c1f7d2f582c63c3cea63d929945[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iad2c780a6386674d50cca54d8c4ebd86     <=
                                             Ib9dfa491b9914f9ac567ae8681a2cd6c[SGN_MAX_SUM_WDTH] ?
                                             ~Ib9dfa491b9914f9ac567ae8681a2cd6c + 1 :
                                             Ib9dfa491b9914f9ac567ae8681a2cd6c
                                             ;

            I925f6b549a25cdc8f85152eb21ea3b58  <=  Ib9dfa491b9914f9ac567ae8681a2cd6c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If1d7944e7c4828ddb91ffea28609cbc7     <=
                                             I029b75f94f58485022bf37590df82900[SGN_MAX_SUM_WDTH] ?
                                             ~I029b75f94f58485022bf37590df82900 + 1 :
                                             I029b75f94f58485022bf37590df82900
                                             ;

            I9b49e1acb81ef5b088b808d2e4ce9954  <=  I029b75f94f58485022bf37590df82900[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I843a68ceb0adab829091f31d0de56eb6     <=
                                             I1cc49a7f6f5c1ecd775d2734c3321364[SGN_MAX_SUM_WDTH] ?
                                             ~I1cc49a7f6f5c1ecd775d2734c3321364 + 1 :
                                             I1cc49a7f6f5c1ecd775d2734c3321364
                                             ;

            I6386a4dd26e7c36165dc265b3a2c93cf  <=  I1cc49a7f6f5c1ecd775d2734c3321364[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I59701b9eb54dda2744a79cebe7d73f3b     <=
                                             I596867e7be52dbcabd95cdd2600396a0[SGN_MAX_SUM_WDTH] ?
                                             ~I596867e7be52dbcabd95cdd2600396a0 + 1 :
                                             I596867e7be52dbcabd95cdd2600396a0
                                             ;

            Ia20709f08cfff3a51d4af1e81d640400  <=  I596867e7be52dbcabd95cdd2600396a0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If63cf5e8f47e4e51176401f0d954ea23     <=
                                             Iec0928bbbc2730b835fb20d75a988a7a[SGN_MAX_SUM_WDTH] ?
                                             ~Iec0928bbbc2730b835fb20d75a988a7a + 1 :
                                             Iec0928bbbc2730b835fb20d75a988a7a
                                             ;

            I1ff042bdb52aac5d69791e96e2f9706c  <=  Iec0928bbbc2730b835fb20d75a988a7a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id09454844b525697de3e3727d89551e4     <=
                                             Iabaf04fabdf2dc5fe29d1eae22b23f7e[SGN_MAX_SUM_WDTH] ?
                                             ~Iabaf04fabdf2dc5fe29d1eae22b23f7e + 1 :
                                             Iabaf04fabdf2dc5fe29d1eae22b23f7e
                                             ;

            Iaa2cbf59f6f61198b4fcf5a741cd5bc8  <=  Iabaf04fabdf2dc5fe29d1eae22b23f7e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6d1b2ce4368945b56eee7814638471cc     <=
                                             I678858a018330bbc4ddb8fe46ff09f49[SGN_MAX_SUM_WDTH] ?
                                             ~I678858a018330bbc4ddb8fe46ff09f49 + 1 :
                                             I678858a018330bbc4ddb8fe46ff09f49
                                             ;

            I01c94743a11042e75638ba6618356203  <=  I678858a018330bbc4ddb8fe46ff09f49[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6079945faa57335b1c902ccf7f960a70     <=
                                             I453a3e7067a9421392ad43b673f203e1[SGN_MAX_SUM_WDTH] ?
                                             ~I453a3e7067a9421392ad43b673f203e1 + 1 :
                                             I453a3e7067a9421392ad43b673f203e1
                                             ;

            I0a0340a0e52145f3597accfe4a4e8624  <=  I453a3e7067a9421392ad43b673f203e1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie7752906ac55cf51f3e96e8c0046f1aa     <=
                                             I1a3dcf633defa34860b0db5fed0d710d[SGN_MAX_SUM_WDTH] ?
                                             ~I1a3dcf633defa34860b0db5fed0d710d + 1 :
                                             I1a3dcf633defa34860b0db5fed0d710d
                                             ;

            I3bb4d24caaa0882a75125e466070f0b1  <=  I1a3dcf633defa34860b0db5fed0d710d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2d7d4135a94f5df949283c043228791f     <=
                                             Id4ba510039040276d71a221b3468977e[SGN_MAX_SUM_WDTH] ?
                                             ~Id4ba510039040276d71a221b3468977e + 1 :
                                             Id4ba510039040276d71a221b3468977e
                                             ;

            I44ead0ab5ccc53226fccc03024643771  <=  Id4ba510039040276d71a221b3468977e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I99c75e3d26c5d01f6ae9abcd05407d8c     <=
                                             I7b9204a45b89e3800944d49a811a930f[SGN_MAX_SUM_WDTH] ?
                                             ~I7b9204a45b89e3800944d49a811a930f + 1 :
                                             I7b9204a45b89e3800944d49a811a930f
                                             ;

            Iaded125f7fd5c833e7206dd7071069be  <=  I7b9204a45b89e3800944d49a811a930f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I81e6f97621dbfb2fed6fc236005a2b19     <=
                                             Ia9d671775a9c5d0c1c0886abc70c5100[SGN_MAX_SUM_WDTH] ?
                                             ~Ia9d671775a9c5d0c1c0886abc70c5100 + 1 :
                                             Ia9d671775a9c5d0c1c0886abc70c5100
                                             ;

            I373be7c3f9511a2906584e33e5048abf  <=  Ia9d671775a9c5d0c1c0886abc70c5100[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ieac60532dcfc916a65054e35cf31d6d2     <=
                                             Ief6f4ea0ada586ed46ce19d0761edf66[SGN_MAX_SUM_WDTH] ?
                                             ~Ief6f4ea0ada586ed46ce19d0761edf66 + 1 :
                                             Ief6f4ea0ada586ed46ce19d0761edf66
                                             ;

            Ie0b5f51835ebdb508a596eeebf0e4847  <=  Ief6f4ea0ada586ed46ce19d0761edf66[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ib7eb83ba73e0dc17f69c357b6ca555bf     <=
                                             I02e35fcbb30d8951f129525146af7f9d[SGN_MAX_SUM_WDTH] ?
                                             ~I02e35fcbb30d8951f129525146af7f9d + 1 :
                                             I02e35fcbb30d8951f129525146af7f9d
                                             ;

            Iddb75e0197b9a76b36a59ac2a7ccdf3a  <=  I02e35fcbb30d8951f129525146af7f9d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5139d8a7a099e3c619c60647c15b7420     <=
                                             Ia55f4e6ae1e56d5aee09414ba7617fc5[SGN_MAX_SUM_WDTH] ?
                                             ~Ia55f4e6ae1e56d5aee09414ba7617fc5 + 1 :
                                             Ia55f4e6ae1e56d5aee09414ba7617fc5
                                             ;

            I08c03198b9599b2f4590e3022e398f7c  <=  Ia55f4e6ae1e56d5aee09414ba7617fc5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6ccd2e11ebd5b2de80b120e20650a602     <=
                                             I4f077fadda92556acba301e0990a8d47[SGN_MAX_SUM_WDTH] ?
                                             ~I4f077fadda92556acba301e0990a8d47 + 1 :
                                             I4f077fadda92556acba301e0990a8d47
                                             ;

            Ia4f3cff223e24815ee1d86bf41756f06  <=  I4f077fadda92556acba301e0990a8d47[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie669cebe5fe39e1a841f8dd3c1f6bc57     <=
                                             I8fc930fd14a7605288eea0d3f7561930[SGN_MAX_SUM_WDTH] ?
                                             ~I8fc930fd14a7605288eea0d3f7561930 + 1 :
                                             I8fc930fd14a7605288eea0d3f7561930
                                             ;

            I56592e1452c4b559af19465b30230ec0  <=  I8fc930fd14a7605288eea0d3f7561930[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If32acb9fc212c4af34099acf6df2bc5a     <=
                                             I29eceabd1f5dfb4cc3028ec248645616[SGN_MAX_SUM_WDTH] ?
                                             ~I29eceabd1f5dfb4cc3028ec248645616 + 1 :
                                             I29eceabd1f5dfb4cc3028ec248645616
                                             ;

            I213ce488e5345fa405a9c5df297d6f74  <=  I29eceabd1f5dfb4cc3028ec248645616[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I075ce236a181bf925c8ccce91d9bc8cd     <=
                                             If55674824a5a3574ffb2f7da75e2f2d3[SGN_MAX_SUM_WDTH] ?
                                             ~If55674824a5a3574ffb2f7da75e2f2d3 + 1 :
                                             If55674824a5a3574ffb2f7da75e2f2d3
                                             ;

            Iefac1e428116a797c2c0803410ac5601  <=  If55674824a5a3574ffb2f7da75e2f2d3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I541d4e422b999a0dfca44d275178e1d9     <=
                                             I12b13bd78932e54099144478a82ae60d[SGN_MAX_SUM_WDTH] ?
                                             ~I12b13bd78932e54099144478a82ae60d + 1 :
                                             I12b13bd78932e54099144478a82ae60d
                                             ;

            I8b419d5827e5b1af9649d602401c189a  <=  I12b13bd78932e54099144478a82ae60d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I3e02657f3d9f79338cd083ed024bf96c     <=
                                             I09a98ded5754d5439ec3a384635d63c8[SGN_MAX_SUM_WDTH] ?
                                             ~I09a98ded5754d5439ec3a384635d63c8 + 1 :
                                             I09a98ded5754d5439ec3a384635d63c8
                                             ;

            Ie989550c9101de382056dd60d5da0e01  <=  I09a98ded5754d5439ec3a384635d63c8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia5e5537405ab8edcc7cd43c86837d43d     <=
                                             I802fd7e7eb9c1b2fd917b1eb657e71b9[SGN_MAX_SUM_WDTH] ?
                                             ~I802fd7e7eb9c1b2fd917b1eb657e71b9 + 1 :
                                             I802fd7e7eb9c1b2fd917b1eb657e71b9
                                             ;

            I259010e323e1e8dcd9dd719091131f6c  <=  I802fd7e7eb9c1b2fd917b1eb657e71b9[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I07ff388e3b6c7288f0f6c35a345023fe     <=
                                             I264cc4045cfc24b211d08488ad2eb105[SGN_MAX_SUM_WDTH] ?
                                             ~I264cc4045cfc24b211d08488ad2eb105 + 1 :
                                             I264cc4045cfc24b211d08488ad2eb105
                                             ;

            I389ac86954fd70464c9550e3fed4ed33  <=  I264cc4045cfc24b211d08488ad2eb105[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I56cb3b3e193ca5068734417fd0ec4e02     <=
                                             Iaa96c298cadeb650acccbd3e548cf281[SGN_MAX_SUM_WDTH] ?
                                             ~Iaa96c298cadeb650acccbd3e548cf281 + 1 :
                                             Iaa96c298cadeb650acccbd3e548cf281
                                             ;

            I77371f0e55b4684d1af196ed52d3d997  <=  Iaa96c298cadeb650acccbd3e548cf281[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I5bbf1765d8f81581d0cf31c0bc755fb3     <=
                                             I463f424b1cc557868a77721849b635a3[SGN_MAX_SUM_WDTH] ?
                                             ~I463f424b1cc557868a77721849b635a3 + 1 :
                                             I463f424b1cc557868a77721849b635a3
                                             ;

            I5a21996f5724a2a49fcf8e928c01b062  <=  I463f424b1cc557868a77721849b635a3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iaa1643095e518846cdede4d5a90dff84     <=
                                             I5fe371b91ca52980957e017a6dbd2308[SGN_MAX_SUM_WDTH] ?
                                             ~I5fe371b91ca52980957e017a6dbd2308 + 1 :
                                             I5fe371b91ca52980957e017a6dbd2308
                                             ;

            Id46108963921efa50aff64d4dd7d1701  <=  I5fe371b91ca52980957e017a6dbd2308[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iee6e12f4717a3279dd31b874eabae69e     <=
                                             Ia301618cac1f678b17595d3e87a85068[SGN_MAX_SUM_WDTH] ?
                                             ~Ia301618cac1f678b17595d3e87a85068 + 1 :
                                             Ia301618cac1f678b17595d3e87a85068
                                             ;

            I8da50e5093acefb6f809aed64564a53e  <=  Ia301618cac1f678b17595d3e87a85068[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic52a9edbbc5283844d2514ea142ca6e2     <=
                                             I0ce7b89ce37757be43c464793608e6da[SGN_MAX_SUM_WDTH] ?
                                             ~I0ce7b89ce37757be43c464793608e6da + 1 :
                                             I0ce7b89ce37757be43c464793608e6da
                                             ;

            I03b0694777d0160a83cbc82ac1397736  <=  I0ce7b89ce37757be43c464793608e6da[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ice3e978c8da2a7de5b28542a5589f0a2     <=
                                             I8abcaf2ec878673e81c94be11046e97e[SGN_MAX_SUM_WDTH] ?
                                             ~I8abcaf2ec878673e81c94be11046e97e + 1 :
                                             I8abcaf2ec878673e81c94be11046e97e
                                             ;

            I85c2bffb93569d9fe1b1bcb10b98bcac  <=  I8abcaf2ec878673e81c94be11046e97e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I336a425aed221c85ca80b9a97d21d6b1     <=
                                             Ie394af0713a3eb30d9d5c0cb38414b90[SGN_MAX_SUM_WDTH] ?
                                             ~Ie394af0713a3eb30d9d5c0cb38414b90 + 1 :
                                             Ie394af0713a3eb30d9d5c0cb38414b90
                                             ;

            Id00274c88b93867a80606343add1cdab  <=  Ie394af0713a3eb30d9d5c0cb38414b90[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie477c0f3b77bb299ba8b1a410d211ef7     <=
                                             Idc8ef4846c1f33c0510b0d4c1b027c81[SGN_MAX_SUM_WDTH] ?
                                             ~Idc8ef4846c1f33c0510b0d4c1b027c81 + 1 :
                                             Idc8ef4846c1f33c0510b0d4c1b027c81
                                             ;

            I61e829cbf7d6c0ef8ddc11677981e2cf  <=  Idc8ef4846c1f33c0510b0d4c1b027c81[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie62920d089ae762603cd33fbf97d92bb     <=
                                             Ib0e1198c7bb8c8bd611fd9afed1bf0ac[SGN_MAX_SUM_WDTH] ?
                                             ~Ib0e1198c7bb8c8bd611fd9afed1bf0ac + 1 :
                                             Ib0e1198c7bb8c8bd611fd9afed1bf0ac
                                             ;

            I9e8ae2aed048068b01b3bd46f30baae8  <=  Ib0e1198c7bb8c8bd611fd9afed1bf0ac[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2ca952e4e676537fd5a8fc71ecfa10e9     <=
                                             Ib2224de3f3f6f644c9e2278ca159eb90[SGN_MAX_SUM_WDTH] ?
                                             ~Ib2224de3f3f6f644c9e2278ca159eb90 + 1 :
                                             Ib2224de3f3f6f644c9e2278ca159eb90
                                             ;

            I7dab71adbe62687846fc027d2789451d  <=  Ib2224de3f3f6f644c9e2278ca159eb90[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iefd31e7ff3c829c88f60bc89d70afcf7     <=
                                             Iad987f88aaf1b32bee71e96904d0c51f[SGN_MAX_SUM_WDTH] ?
                                             ~Iad987f88aaf1b32bee71e96904d0c51f + 1 :
                                             Iad987f88aaf1b32bee71e96904d0c51f
                                             ;

            If1295608bd218ed60922a0b95bf1d098  <=  Iad987f88aaf1b32bee71e96904d0c51f[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iafa987a413fd8fcacfe872bc0f5bc2d6     <=
                                             I0831e757dd5e5868bb023dd9004fb68a[SGN_MAX_SUM_WDTH] ?
                                             ~I0831e757dd5e5868bb023dd9004fb68a + 1 :
                                             I0831e757dd5e5868bb023dd9004fb68a
                                             ;

            Idf04e08c120ed116af14a62659675b44  <=  I0831e757dd5e5868bb023dd9004fb68a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I305c1ea420d666f258e38c5a65847367     <=
                                             I64b4330df88134dffb32e0dfd8d4ab36[SGN_MAX_SUM_WDTH] ?
                                             ~I64b4330df88134dffb32e0dfd8d4ab36 + 1 :
                                             I64b4330df88134dffb32e0dfd8d4ab36
                                             ;

            Ieb7614ad1b1bfed3e2b0089a72fe214a  <=  I64b4330df88134dffb32e0dfd8d4ab36[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9f040c4088bfab72d74e5332e9710d1a     <=
                                             I5066c1fb5193c037de084c7463947151[SGN_MAX_SUM_WDTH] ?
                                             ~I5066c1fb5193c037de084c7463947151 + 1 :
                                             I5066c1fb5193c037de084c7463947151
                                             ;

            I589062eca318b25dfe5735da455b6fe1  <=  I5066c1fb5193c037de084c7463947151[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia2f41f9778324a06daeb185c736516a4     <=
                                             I76c57762b38b9546bc862bccfde73a81[SGN_MAX_SUM_WDTH] ?
                                             ~I76c57762b38b9546bc862bccfde73a81 + 1 :
                                             I76c57762b38b9546bc862bccfde73a81
                                             ;

            If3db87afb3ea184c9e4020c5e45cb161  <=  I76c57762b38b9546bc862bccfde73a81[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id9778ba5fbdbed4d33a092da6b68c414     <=
                                             I4720972ec687864e66b86780a4a03e47[SGN_MAX_SUM_WDTH] ?
                                             ~I4720972ec687864e66b86780a4a03e47 + 1 :
                                             I4720972ec687864e66b86780a4a03e47
                                             ;

            Ia14bc1fcd5bbdcb60b8e68298f7d716a  <=  I4720972ec687864e66b86780a4a03e47[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I27c2c79d0d719c71c8e28218d1174a13     <=
                                             Ib0da91fdb282ea40f13881671d9736b3[SGN_MAX_SUM_WDTH] ?
                                             ~Ib0da91fdb282ea40f13881671d9736b3 + 1 :
                                             Ib0da91fdb282ea40f13881671d9736b3
                                             ;

            I268b60cb371b3d46dc3f8b0009f541b1  <=  Ib0da91fdb282ea40f13881671d9736b3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2a9d6a774769b12ae20bc0cee0c36f5c     <=
                                             Ifac345df39972bcecf0cf454e30c0cea[SGN_MAX_SUM_WDTH] ?
                                             ~Ifac345df39972bcecf0cf454e30c0cea + 1 :
                                             Ifac345df39972bcecf0cf454e30c0cea
                                             ;

            If2cd93b57cd1c2b91ee7a73a97dd19f2  <=  Ifac345df39972bcecf0cf454e30c0cea[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I2c567b75f1399c069b95284f4c36b6d1     <=
                                             I47ee2c7239716a56029d9d7dd2efeec2[SGN_MAX_SUM_WDTH] ?
                                             ~I47ee2c7239716a56029d9d7dd2efeec2 + 1 :
                                             I47ee2c7239716a56029d9d7dd2efeec2
                                             ;

            Id81305359a07db527e49fda05cd2784f  <=  I47ee2c7239716a56029d9d7dd2efeec2[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If3d3eb609abfd6e315eec803d2e94490     <=
                                             I02398b40df5e80a6818d7f7c20896897[SGN_MAX_SUM_WDTH] ?
                                             ~I02398b40df5e80a6818d7f7c20896897 + 1 :
                                             I02398b40df5e80a6818d7f7c20896897
                                             ;

            Id8292eca087c1a17dc8b5a572a76f21f  <=  I02398b40df5e80a6818d7f7c20896897[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9c58aea7ce986b1d28f5808b347c015d     <=
                                             I5943d30c92a0938ea3933ba61819ce91[SGN_MAX_SUM_WDTH] ?
                                             ~I5943d30c92a0938ea3933ba61819ce91 + 1 :
                                             I5943d30c92a0938ea3933ba61819ce91
                                             ;

            Iddb19725b093506e5e521d8d68dcb8e1  <=  I5943d30c92a0938ea3933ba61819ce91[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Id139c7a783196941100003b6cb0cd1e7     <=
                                             Iab0a2d1699d14959918590a17d221dac[SGN_MAX_SUM_WDTH] ?
                                             ~Iab0a2d1699d14959918590a17d221dac + 1 :
                                             Iab0a2d1699d14959918590a17d221dac
                                             ;

            I0b573d3a86a3111451da661e46384876  <=  Iab0a2d1699d14959918590a17d221dac[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I524d7614b01460778da3ce98f6aaa3d9     <=
                                             If30544b94b0d43b30a8e4a1a6f67e461[SGN_MAX_SUM_WDTH] ?
                                             ~If30544b94b0d43b30a8e4a1a6f67e461 + 1 :
                                             If30544b94b0d43b30a8e4a1a6f67e461
                                             ;

            I0ff479e61d1a0cede88ebffb073c60be  <=  If30544b94b0d43b30a8e4a1a6f67e461[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8acda65f116d5c91cbe2662ac282aa31     <=
                                             I4d6cdcb3b63c51d9dd8b915eb0645255[SGN_MAX_SUM_WDTH] ?
                                             ~I4d6cdcb3b63c51d9dd8b915eb0645255 + 1 :
                                             I4d6cdcb3b63c51d9dd8b915eb0645255
                                             ;

            Icd6f8f5df6b4ca4c81855e974db76526  <=  I4d6cdcb3b63c51d9dd8b915eb0645255[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If67dbe22f8d22b3430215fb0deae8204     <=
                                             Id147fa768121368db44934717c87f635[SGN_MAX_SUM_WDTH] ?
                                             ~Id147fa768121368db44934717c87f635 + 1 :
                                             Id147fa768121368db44934717c87f635
                                             ;

            I7ce064a756dad56d37684d5d7d168047  <=  Id147fa768121368db44934717c87f635[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9a35cd7512787263abedd6d9913cf507     <=
                                             I7f67e05ed60a537f26feebbbe643a67c[SGN_MAX_SUM_WDTH] ?
                                             ~I7f67e05ed60a537f26feebbbe643a67c + 1 :
                                             I7f67e05ed60a537f26feebbbe643a67c
                                             ;

            Ied2ea62cfb21602645babc36e27b8218  <=  I7f67e05ed60a537f26feebbbe643a67c[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9cca23469c5e6001650f1f8b1360ae8     <=
                                             I376c401480a2d8e6131123a91e6fa1cc[SGN_MAX_SUM_WDTH] ?
                                             ~I376c401480a2d8e6131123a91e6fa1cc + 1 :
                                             I376c401480a2d8e6131123a91e6fa1cc
                                             ;

            I79b85da6e5ce0b02ebd1619115c98e24  <=  I376c401480a2d8e6131123a91e6fa1cc[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icc2606ae8f9a3b425225ae7339112b9d     <=
                                             Ic33856f32df0ab980accff5678cceebb[SGN_MAX_SUM_WDTH] ?
                                             ~Ic33856f32df0ab980accff5678cceebb + 1 :
                                             Ic33856f32df0ab980accff5678cceebb
                                             ;

            I8e1ddd7e4185c28caa71d30bc28138f3  <=  Ic33856f32df0ab980accff5678cceebb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I34aa1802d24e074ae54563898929abfa     <=
                                             I97e41b86305179e201cce4d69c2ffa21[SGN_MAX_SUM_WDTH] ?
                                             ~I97e41b86305179e201cce4d69c2ffa21 + 1 :
                                             I97e41b86305179e201cce4d69c2ffa21
                                             ;

            Iab0bff1633e2f3ea0bfbc291f3ab5d29  <=  I97e41b86305179e201cce4d69c2ffa21[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Icb85b3464dc40e8504c53c377e889c45     <=
                                             Iecaf532a526a0f689b65a6dd749d66cf[SGN_MAX_SUM_WDTH] ?
                                             ~Iecaf532a526a0f689b65a6dd749d66cf + 1 :
                                             Iecaf532a526a0f689b65a6dd749d66cf
                                             ;

            I5f0751fceaa008feba5c6867ced453dc  <=  Iecaf532a526a0f689b65a6dd749d66cf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie595a7d10b5ac84c0301fb55bebd3680     <=
                                             Ia54ab64aa44544f38180c57e0864e071[SGN_MAX_SUM_WDTH] ?
                                             ~Ia54ab64aa44544f38180c57e0864e071 + 1 :
                                             Ia54ab64aa44544f38180c57e0864e071
                                             ;

            I9f6751c15237c20b0cf2175575195ea7  <=  Ia54ab64aa44544f38180c57e0864e071[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9c217a672cabc05efbdff218637123ba     <=
                                             I8ed5770ee3c9a504d934506743f6b427[SGN_MAX_SUM_WDTH] ?
                                             ~I8ed5770ee3c9a504d934506743f6b427 + 1 :
                                             I8ed5770ee3c9a504d934506743f6b427
                                             ;

            I6ea50be10bc990a1206cdc9e28e0c4c2  <=  I8ed5770ee3c9a504d934506743f6b427[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If20f3780b4af857ffe8083056085517a     <=
                                             I7541c0e729546e0e13e98f4658b95a1d[SGN_MAX_SUM_WDTH] ?
                                             ~I7541c0e729546e0e13e98f4658b95a1d + 1 :
                                             I7541c0e729546e0e13e98f4658b95a1d
                                             ;

            I43c2fab87f70ea883321ab82de85f133  <=  I7541c0e729546e0e13e98f4658b95a1d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic2e275bfa8ab3d2002d2aa374ac9bfe2     <=
                                             Id861f8b6cc578cfb1d83d065ae78dedb[SGN_MAX_SUM_WDTH] ?
                                             ~Id861f8b6cc578cfb1d83d065ae78dedb + 1 :
                                             Id861f8b6cc578cfb1d83d065ae78dedb
                                             ;

            I1af02ed6cf00d4cb0704b5e44c83bfa3  <=  Id861f8b6cc578cfb1d83d065ae78dedb[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Iac5798fd9915b6778700da6a14f6a381     <=
                                             I6fd4a37bc3b6eb96e6b7e814b203ed21[SGN_MAX_SUM_WDTH] ?
                                             ~I6fd4a37bc3b6eb96e6b7e814b203ed21 + 1 :
                                             I6fd4a37bc3b6eb96e6b7e814b203ed21
                                             ;

            Ib71611afdd0381cc1884f5ddbbae1acc  <=  I6fd4a37bc3b6eb96e6b7e814b203ed21[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ide3204bf317fdfb993410d338085b174     <=
                                             Ie31fceaf1518af42616d21bd8247577a[SGN_MAX_SUM_WDTH] ?
                                             ~Ie31fceaf1518af42616d21bd8247577a + 1 :
                                             Ie31fceaf1518af42616d21bd8247577a
                                             ;

            I38fc49afce0298846ae8ed63ae715e81  <=  Ie31fceaf1518af42616d21bd8247577a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ic3a95140fc1029efa17a6557bc977719     <=
                                             I89ecfbed8d99ec79402dd5f3f1e64100[SGN_MAX_SUM_WDTH] ?
                                             ~I89ecfbed8d99ec79402dd5f3f1e64100 + 1 :
                                             I89ecfbed8d99ec79402dd5f3f1e64100
                                             ;

            Iddc3e44d83e8253e5129b6cbf5082df7  <=  I89ecfbed8d99ec79402dd5f3f1e64100[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I647d3a46bb2c7ed0f1ec08760b3858be     <=
                                             Iddde66a99ea9a0caa45b06e168194488[SGN_MAX_SUM_WDTH] ?
                                             ~Iddde66a99ea9a0caa45b06e168194488 + 1 :
                                             Iddde66a99ea9a0caa45b06e168194488
                                             ;

            I975a87bdda30c5b6be8d2f0e4b107450  <=  Iddde66a99ea9a0caa45b06e168194488[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4816747af9d9fc8dc85fd831336ec710     <=
                                             Ib645c9e05a543ca3e8ce0994e56aac70[SGN_MAX_SUM_WDTH] ?
                                             ~Ib645c9e05a543ca3e8ce0994e56aac70 + 1 :
                                             Ib645c9e05a543ca3e8ce0994e56aac70
                                             ;

            I582bd96afa764ded148202f738b7a1df  <=  Ib645c9e05a543ca3e8ce0994e56aac70[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1f66c026a5437320bd1f4df2ff71663d     <=
                                             I29fedc646a3ba823d0dcbb3ecb9b9ad6[SGN_MAX_SUM_WDTH] ?
                                             ~I29fedc646a3ba823d0dcbb3ecb9b9ad6 + 1 :
                                             I29fedc646a3ba823d0dcbb3ecb9b9ad6
                                             ;

            I6fb88d97bc9ed37a06b729020a1df140  <=  I29fedc646a3ba823d0dcbb3ecb9b9ad6[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If347c58c328193f420286ea27a4afa20     <=
                                             Ie89f6128d6d68c146ffcecb551618321[SGN_MAX_SUM_WDTH] ?
                                             ~Ie89f6128d6d68c146ffcecb551618321 + 1 :
                                             Ie89f6128d6d68c146ffcecb551618321
                                             ;

            I1500943c4a550e78fc169437b0a663b7  <=  Ie89f6128d6d68c146ffcecb551618321[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I7a126c8304be920f2a920315dc61ba7f     <=
                                             I3388d6fa5159183888944f2951de9361[SGN_MAX_SUM_WDTH] ?
                                             ~I3388d6fa5159183888944f2951de9361 + 1 :
                                             I3388d6fa5159183888944f2951de9361
                                             ;

            I0b83f4ef8ba9badb27e81b32765ec5b6  <=  I3388d6fa5159183888944f2951de9361[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I237327d6a74df1fb05537dc3691ebf11     <=
                                             I3575e2d60ee8b0b71c67d53b496e2775[SGN_MAX_SUM_WDTH] ?
                                             ~I3575e2d60ee8b0b71c67d53b496e2775 + 1 :
                                             I3575e2d60ee8b0b71c67d53b496e2775
                                             ;

            I2c420acf428e44cdd9ca9998e276f258  <=  I3575e2d60ee8b0b71c67d53b496e2775[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I64a3e8bb4c87b066806d33a5306a2c53     <=
                                             I52cf4fceee16d75ea59dbb574ea7c7b0[SGN_MAX_SUM_WDTH] ?
                                             ~I52cf4fceee16d75ea59dbb574ea7c7b0 + 1 :
                                             I52cf4fceee16d75ea59dbb574ea7c7b0
                                             ;

            Ic7b6dae3017b55dd3cd27423d5f1b0ec  <=  I52cf4fceee16d75ea59dbb574ea7c7b0[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ibbca6ec39234473fb517447a8beacafc     <=
                                             I59cfcae849791453127d60b213ff7355[SGN_MAX_SUM_WDTH] ?
                                             ~I59cfcae849791453127d60b213ff7355 + 1 :
                                             I59cfcae849791453127d60b213ff7355
                                             ;

            I4a91a7c9b2a0f3552b8f2ef4e2398be2  <=  I59cfcae849791453127d60b213ff7355[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I78327356176a16fc996188b83b058cbc     <=
                                             Ic218ffc97e5e89851d44554326aa5bae[SGN_MAX_SUM_WDTH] ?
                                             ~Ic218ffc97e5e89851d44554326aa5bae + 1 :
                                             Ic218ffc97e5e89851d44554326aa5bae
                                             ;

            I99ff29c7ba68b5d0819f1e1bead51287  <=  Ic218ffc97e5e89851d44554326aa5bae[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifec496c87a7a2474855067305ac8cba3     <=
                                             I6886b93a81c52c7f93b506404b6a4252[SGN_MAX_SUM_WDTH] ?
                                             ~I6886b93a81c52c7f93b506404b6a4252 + 1 :
                                             I6886b93a81c52c7f93b506404b6a4252
                                             ;

            If06b00be0356a2be5074d958ddcdb2f9  <=  I6886b93a81c52c7f93b506404b6a4252[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I41584165a62caaa37ddebbf79bb8b617     <=
                                             Id9c9ac52a48ef3207581bd31c0593b22[SGN_MAX_SUM_WDTH] ?
                                             ~Id9c9ac52a48ef3207581bd31c0593b22 + 1 :
                                             Id9c9ac52a48ef3207581bd31c0593b22
                                             ;

            I604283449f13c7b225ea03f99f2e296a  <=  Id9c9ac52a48ef3207581bd31c0593b22[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Idf0916d6b025aad6eccb98ada5ba3aca     <=
                                             Ib3c08e618350ef723607b4ee58bb4dd1[SGN_MAX_SUM_WDTH] ?
                                             ~Ib3c08e618350ef723607b4ee58bb4dd1 + 1 :
                                             Ib3c08e618350ef723607b4ee58bb4dd1
                                             ;

            I2b600e5f5c146ee97c4044c08e1f5ad5  <=  Ib3c08e618350ef723607b4ee58bb4dd1[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I00ef133d5a53f8f99f35b50327e5272b     <=
                                             I2481f5b76264c857df96942bdaa941ca[SGN_MAX_SUM_WDTH] ?
                                             ~I2481f5b76264c857df96942bdaa941ca + 1 :
                                             I2481f5b76264c857df96942bdaa941ca
                                             ;

            I9fe16403fc21bb1159a5e0305fd1ef69  <=  I2481f5b76264c857df96942bdaa941ca[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I6f0e302d38d75982d0761e306ce9f146     <=
                                             I3a5aa34be4c3adccf4aad2772c38e972[SGN_MAX_SUM_WDTH] ?
                                             ~I3a5aa34be4c3adccf4aad2772c38e972 + 1 :
                                             I3a5aa34be4c3adccf4aad2772c38e972
                                             ;

            Iabdb9374e5caee281c25b003624b2c4e  <=  I3a5aa34be4c3adccf4aad2772c38e972[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I127eed5de00e10a020717e796de76c7d     <=
                                             I95b6796cf442383290a32bad614664e8[SGN_MAX_SUM_WDTH] ?
                                             ~I95b6796cf442383290a32bad614664e8 + 1 :
                                             I95b6796cf442383290a32bad614664e8
                                             ;

            Ibd12036702fe60b57354b3aac921559d  <=  I95b6796cf442383290a32bad614664e8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If9aad73aefb1b225f35e8c813b85fe87     <=
                                             Ie45ac55c4add6c3390924c54d2e8d65e[SGN_MAX_SUM_WDTH] ?
                                             ~Ie45ac55c4add6c3390924c54d2e8d65e + 1 :
                                             Ie45ac55c4add6c3390924c54d2e8d65e
                                             ;

            Ib1639811de6eb1c38257800c201fb704  <=  Ie45ac55c4add6c3390924c54d2e8d65e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I00a89ac37676521a081a21b1ec1a0798     <=
                                             I0935498f4dd90c1fed52d2246ebe326b[SGN_MAX_SUM_WDTH] ?
                                             ~I0935498f4dd90c1fed52d2246ebe326b + 1 :
                                             I0935498f4dd90c1fed52d2246ebe326b
                                             ;

            If926d98f659e8fe4bbf36ad2c5c852c5  <=  I0935498f4dd90c1fed52d2246ebe326b[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I06f3a34f2b1770ef82ddc2a732b3d4fb     <=
                                             Iac314ba0cecbd52f3992323dbce81856[SGN_MAX_SUM_WDTH] ?
                                             ~Iac314ba0cecbd52f3992323dbce81856 + 1 :
                                             Iac314ba0cecbd52f3992323dbce81856
                                             ;

            I211f8d7f97ebb8eb3e50313513abfb1b  <=  Iac314ba0cecbd52f3992323dbce81856[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I4744d64a746f16004e3bedaaa41465f1     <=
                                             I2f8a71c2c9078e2581087c7662c961f4[SGN_MAX_SUM_WDTH] ?
                                             ~I2f8a71c2c9078e2581087c7662c961f4 + 1 :
                                             I2f8a71c2c9078e2581087c7662c961f4
                                             ;

            I304ac9f96945546cdf1b6f1fa7136731  <=  I2f8a71c2c9078e2581087c7662c961f4[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ifae0cc6cc1c65d24bbe84c4ba938e2ea     <=
                                             I38c53b94ea9a59a52cdcfe6681491da8[SGN_MAX_SUM_WDTH] ?
                                             ~I38c53b94ea9a59a52cdcfe6681491da8 + 1 :
                                             I38c53b94ea9a59a52cdcfe6681491da8
                                             ;

            I7a9800418bd5c195fc47a72370680b56  <=  I38c53b94ea9a59a52cdcfe6681491da8[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1223c21129382d41e4f38ef4bbe60c2f     <=
                                             I5c2c6a0ca07e820e699062299b7064e3[SGN_MAX_SUM_WDTH] ?
                                             ~I5c2c6a0ca07e820e699062299b7064e3 + 1 :
                                             I5c2c6a0ca07e820e699062299b7064e3
                                             ;

            I5f6a61c9f0c67510e148e596f553a4d6  <=  I5c2c6a0ca07e820e699062299b7064e3[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I14e36e16df00adcd7dc1973d3852d2d9     <=
                                             Ia962052eea10222a1c16ce5800e1c063[SGN_MAX_SUM_WDTH] ?
                                             ~Ia962052eea10222a1c16ce5800e1c063 + 1 :
                                             Ia962052eea10222a1c16ce5800e1c063
                                             ;

            I8e313ceb21359bcc44114ab217b1c394  <=  Ia962052eea10222a1c16ce5800e1c063[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0d05ae27b53fb6939e4c2f862a8d20b2     <=
                                             I33ecd2de3fc7f48821e40313b5dc2093[SGN_MAX_SUM_WDTH] ?
                                             ~I33ecd2de3fc7f48821e40313b5dc2093 + 1 :
                                             I33ecd2de3fc7f48821e40313b5dc2093
                                             ;

            I4c9518755c33d725221ad79ee6badba9  <=  I33ecd2de3fc7f48821e40313b5dc2093[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I97a6fcc08929c3b7d15e36d7706ed13d     <=
                                             Ie4d5fc4a5bf560bf75561f7f6baa761e[SGN_MAX_SUM_WDTH] ?
                                             ~Ie4d5fc4a5bf560bf75561f7f6baa761e + 1 :
                                             Ie4d5fc4a5bf560bf75561f7f6baa761e
                                             ;

            I3c3cffec9f47c9979cb9503f222f370c  <=  Ie4d5fc4a5bf560bf75561f7f6baa761e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I1f04e86bf27596718836d0a09adbe120     <=
                                             I57de351c4dcc2f9c6bacdf1f39961723[SGN_MAX_SUM_WDTH] ?
                                             ~I57de351c4dcc2f9c6bacdf1f39961723 + 1 :
                                             I57de351c4dcc2f9c6bacdf1f39961723
                                             ;

            I68d6769541fdc3df321e192f645c667f  <=  I57de351c4dcc2f9c6bacdf1f39961723[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie40873cfd6d10a61a94a761becf588a8     <=
                                             Ibf1a5a90d4a7922c4bd6273c9a3f1701[SGN_MAX_SUM_WDTH] ?
                                             ~Ibf1a5a90d4a7922c4bd6273c9a3f1701 + 1 :
                                             Ibf1a5a90d4a7922c4bd6273c9a3f1701
                                             ;

            Ided55428cbb77f454c2607ac783d7548  <=  Ibf1a5a90d4a7922c4bd6273c9a3f1701[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I61960ed74fee948cc12bd1fd8384559a     <=
                                             I8a9e51ef30c6434e44fe23412d20425a[SGN_MAX_SUM_WDTH] ?
                                             ~I8a9e51ef30c6434e44fe23412d20425a + 1 :
                                             I8a9e51ef30c6434e44fe23412d20425a
                                             ;

            Ifd3d4f3e2a388b3c70e7704d6351e0ba  <=  I8a9e51ef30c6434e44fe23412d20425a[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I8533a3ec4be4c49166184c94761eaebc     <=
                                             I796d4045b29e6c1100dfed4a78dbb912[SGN_MAX_SUM_WDTH] ?
                                             ~I796d4045b29e6c1100dfed4a78dbb912 + 1 :
                                             I796d4045b29e6c1100dfed4a78dbb912
                                             ;

            I17d32f292758416fe02527dfd938fa0d  <=  I796d4045b29e6c1100dfed4a78dbb912[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I00be319b5bdb85ffaf3bb0eca0b348b6     <=
                                             I32551e388a1ee2ecc7d7da3a4646177e[SGN_MAX_SUM_WDTH] ?
                                             ~I32551e388a1ee2ecc7d7da3a4646177e + 1 :
                                             I32551e388a1ee2ecc7d7da3a4646177e
                                             ;

            I9ce3942aba354c1fd7d6b9a39c994d7b  <=  I32551e388a1ee2ecc7d7da3a4646177e[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ie889c916b5af185b52ff5e2e3cc23045     <=
                                             I6c266cffd4d2836af16d4d81bbd11250[SGN_MAX_SUM_WDTH] ?
                                             ~I6c266cffd4d2836af16d4d81bbd11250 + 1 :
                                             I6c266cffd4d2836af16d4d81bbd11250
                                             ;

            I2c6c6041c9c69c84f4d64af6458955f5  <=  I6c266cffd4d2836af16d4d81bbd11250[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I89697be6dcb2e7f972db498c1b1dea71     <=
                                             I9feff48bffd8e1f9eee0a587b4b026d5[SGN_MAX_SUM_WDTH] ?
                                             ~I9feff48bffd8e1f9eee0a587b4b026d5 + 1 :
                                             I9feff48bffd8e1f9eee0a587b4b026d5
                                             ;

            I830a4fffe1244e071eb82c28ddc4a308  <=  I9feff48bffd8e1f9eee0a587b4b026d5[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If13dfbfff7cd8e197bb44006a3db73bf     <=
                                             I6c540a2cc92ae1fc269a3a395504a08d[SGN_MAX_SUM_WDTH] ?
                                             ~I6c540a2cc92ae1fc269a3a395504a08d + 1 :
                                             I6c540a2cc92ae1fc269a3a395504a08d
                                             ;

            Ifad8e46fc3844bbfaf434a14f6b5869d  <=  I6c540a2cc92ae1fc269a3a395504a08d[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I87ed6c3e172c7a06bf6aefe7bf718d70     <=
                                             I683c93eb9205a2272d286e4ad0e998fe[SGN_MAX_SUM_WDTH] ?
                                             ~I683c93eb9205a2272d286e4ad0e998fe + 1 :
                                             I683c93eb9205a2272d286e4ad0e998fe
                                             ;

            I10a6c6a8fdb0003de1f360c148777d0f  <=  I683c93eb9205a2272d286e4ad0e998fe[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I0db87adc849839fab3a4c9884d5a4882     <=
                                             Ic92cbaba339661a83c8bbd3f8377c105[SGN_MAX_SUM_WDTH] ?
                                             ~Ic92cbaba339661a83c8bbd3f8377c105 + 1 :
                                             Ic92cbaba339661a83c8bbd3f8377c105
                                             ;

            I4cde586fc28f8d03fc9934d56f7ff7b8  <=  Ic92cbaba339661a83c8bbd3f8377c105[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I535e01a6c35fd7b455e4b79b1d4bb414     <=
                                             I81850f6963cf07be478907b167cf9206[SGN_MAX_SUM_WDTH] ?
                                             ~I81850f6963cf07be478907b167cf9206 + 1 :
                                             I81850f6963cf07be478907b167cf9206
                                             ;

            Ib83a067fb08e118dcf794902beef9405  <=  I81850f6963cf07be478907b167cf9206[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            Ia2d1c752cc4b405adb97a815e90a7b96     <=
                                             I6d94790ac6714bb8c62a82bb06960fbf[SGN_MAX_SUM_WDTH] ?
                                             ~I6d94790ac6714bb8c62a82bb06960fbf + 1 :
                                             I6d94790ac6714bb8c62a82bb06960fbf
                                             ;

            I358cf9609272a4562423a85f9b2f56bf  <=  I6d94790ac6714bb8c62a82bb06960fbf[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            I9ac12eb3878f6fc7dc428fe5e7f35d97     <=
                                             Ie19542cb6dc9324368b1ea75a5d5c274[SGN_MAX_SUM_WDTH] ?
                                             ~Ie19542cb6dc9324368b1ea75a5d5c274 + 1 :
                                             Ie19542cb6dc9324368b1ea75a5d5c274
                                             ;

            Ic1e9d9113150ad57954c0e369259dc62  <=  Ie19542cb6dc9324368b1ea75a5d5c274[SGN_MAX_SUM_WDTH] ;

           end
           if (I3c62d5bd891bd3750b7bd1d32612f589) begin
            If46fa11dfadb0691eaaa0a40836e08d8     <=
                                             I6c96e6686c458cee66b9d93d6d71f350[SGN_MAX_SUM_WDTH] ?
                                             ~I6c96e6686c458cee66b9d93d6d71f350 + 1 :
                                             I6c96e6686c458cee66b9d93d6d71f350
                                             ;

            If7fe3f5ccbb5b279e41fd183c8ff3974  <=  I6c96e6686c458cee66b9d93d6d71f350[SGN_MAX_SUM_WDTH] ;

           end
       end

   end

assign Ic05b492587d8d5083e8570900995293a      = I748f85f6680918a2e992df339b4b6558 +  ~Iea07d1adf9016a29cffd61d183e268d0 +1;
assign Ibee9ba58404f1adb9e4e8e6f822a38c1      = I748f85f6680918a2e992df339b4b6558 +  ~If92db65b39a83e1c699e4cc6d7f9e57b +1;
assign Ifab38317b76e52f9d9d64bed976e2cc5      = I748f85f6680918a2e992df339b4b6558 +  ~I8f2986bc015fcc64ac5e5395ac6dd851 +1;
assign I86195d9a1da88ffc163298c54401039e      = I748f85f6680918a2e992df339b4b6558 +  ~I355725a804e0df68b4acf96ca98f2448 +1;
assign I27c02895bfd59c762d5c7a725aa5cefd      = I748f85f6680918a2e992df339b4b6558 +  ~I78212ae965ab2dcb2eed0b060d6b253f +1;
assign I60de515e03218ac363566ce7b92f5034      = I748f85f6680918a2e992df339b4b6558 +  ~I0b56aa7a1b7549c91dddd3a06ecbaacf +1;
assign I9b75e7451fbf27c3645bebbdba234996      = I748f85f6680918a2e992df339b4b6558 +  ~I71412803cc5229025487255aec62ec4f +1;
assign I056c79002bbba10ddee2448e36dc7478      = I748f85f6680918a2e992df339b4b6558 +  ~I32fcb28a27356bc6f403528836ea4c1f +1;
assign Ia5db5f66b7fb04e2344abff9b4f75404      = I748f85f6680918a2e992df339b4b6558 +  ~Iad354d876cb9fc72fc0143e6f7da9357 +1;
assign I250898de23a8793f0c21eb333d61af53      = I748f85f6680918a2e992df339b4b6558 +  ~If6e745bb85abba7282dae1f6f701225e +1;
assign I1320273c298c7953b3227b58439b54c4      = I748f85f6680918a2e992df339b4b6558 +  ~I93bb43c1b89d4c70a57bdc019d64fd22 +1;
assign I49a036af196fb318309a43c150540a2c      = I748f85f6680918a2e992df339b4b6558 +  ~I7a2e554d07bbea291f2cfc18694fca3a +1;
assign If115c3e5f121363c2b8a6c14905aebe7      = I748f85f6680918a2e992df339b4b6558 +  ~I3e59b2419c7dd1553b792d536208514e +1;
assign I5fcd95690fb291f9b95996e687de022c      = I748f85f6680918a2e992df339b4b6558 +  ~I46894c6526983bf1ce4b503159131b41 +1;
assign I5f6f8a4c5c5ab4cf1f9c496795c41ce8      = I748f85f6680918a2e992df339b4b6558 +  ~I6404d0df952b5bf8292c753e4c6f35d8 +1;
assign I775180b845280ec240e4adf20605b8fe      = I748f85f6680918a2e992df339b4b6558 +  ~I8522c402e654d007abffcb0e904af5e6 +1;
assign I642fe2c7978d7229d660431061a6f781      = I748f85f6680918a2e992df339b4b6558 +  ~I5ed85845c39337c37791f16e718069b4 +1;
assign I3ce66aa6048542c81a89c28e80412e70      = I748f85f6680918a2e992df339b4b6558 +  ~I89013d61c1ea8da8b1c6071cc21c316f +1;
assign I436fc89b03a41f35b8d2ab89464d07c0      = I748f85f6680918a2e992df339b4b6558 +  ~I4102100fa5f1dd299af0190862efcc42 +1;
assign I67861da88ed0edc52bb876287fc60261      = I748f85f6680918a2e992df339b4b6558 +  ~I4939f69abb1eac56d5021e06406a93b5 +1;
assign If51bec96c3139419947f0442b0ad7281      = I748f85f6680918a2e992df339b4b6558 +  ~Iadbd245bf842aebb456417579a3e6296 +1;
assign I5e126994711cd1782fcbd2fb3eec3cdc      = I748f85f6680918a2e992df339b4b6558 +  ~Ifc8ece44a4e68c3117eda9e65f3084d2 +1;
assign I44d2fe323e921ba0fd66c82a792302e1      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I91679dfab57a372eddc7f9b94a231edb +1;
assign I875b53feb16dc1ac263e9d1c2552dd38      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I2213c1a2b831f421707a261f5a58b1b1 +1;
assign I651f168318d2ce4746ade3230e052ace      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ic53b875b2ddcba11406eb2ca39354757 +1;
assign I00a65dc6a94fa280ec3aac7b04fd4aba      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I634484f00590216c0f74f975c9c83400 +1;
assign I38f5eb8d994476d2edb5fd71b7636452      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ib3b1db2d8b669988c887ed780e439b26 +1;
assign If0d9102fbff225bd3ef4f4e1aab2811b      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I735db8b0ee0ec98e4cce0030b11508da +1;
assign I09734a3840b1b01a467b075c65608f3e      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~If1607e907e626902ee26d15020a64c21 +1;
assign Icec563470fe1bec10dfa8d36561f6ed7      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I081b38dbb37d4c14a6a9fd3fefa13daa +1;
assign Iaa82bbd78ea7acbc1949f7db44d339eb      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ibac5e7b6d4bf5cd6926358318f0c418f +1;
assign I1bf879a8671257cec876577804bd6ffb      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Iadfc60386481092ae85cc148a2c40abb +1;
assign Ifdb571f08bb8fc78631b0af95d6f5b68      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ie0ee5445c56a5f9b41640b57422206de +1;
assign I06117d4a9cec69582f336796f82af871      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ie5f8620371236cb11c9e88c16b509ee8 +1;
assign I23178a40d717727916e4c44fb8ea7de9      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I8d7c1fe2e33bbd45379b0325a3c5e989 +1;
assign Idd1454bc7f85ca3c184a20fd0864c666      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I4fbdc4ee57a3be42b62d9bd43078d6ef +1;
assign Iee01a4b6a910ede0b61e2465d7d5d696      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I5510b88bfd65811b3200adf4ef975b48 +1;
assign I383d6b1028ae1e4e2ea40cfa22043d72      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~Ib57ef2f577cca54713c16717cbbd1ce9 +1;
assign Ifde4b0c41d42daf9b134ee6c05db336a      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I15943aa74e9fbbaebdc0d54eb6a3bffa +1;
assign I9f0b1952f54a14726de1d31a2302a95f      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I6ac24c46319a787daa5c545de8c6eeea +1;
assign I3991c8d4f24af7dfb52a65f70c3ab2d5      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I52403a0454e5fa002e79eaab7ea497bd +1;
assign Ie928ef6ba83900dca8b150428d713448      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I634f0ce28934600a1a31ab0d8e59b4a9 +1;
assign Ic085f1faeb81e3027f909a7bd890d359      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I7103aa739616a39c03e675ea0efb0335 +1;
assign I159df37fedc1447f6766308aa58ff70c      = Ib0f57837099e3fdf1b908d78bcda4a43 +  ~I0296d01fd3f9a269a617efd4beea9b8b +1;
assign I53491740a9877fcff56e6a3d8ac61643      = If75e99660e3997f53f7b903bc366f47f +  ~I065a81ba25962785215583e7ece27661 +1;
assign If9eba70be918197cc0bb2974f04c0687      = If75e99660e3997f53f7b903bc366f47f +  ~I631a3300cb6685f47da7781940ec5d27 +1;
assign I2a30d44d2006f17582bb431e397d3874      = If75e99660e3997f53f7b903bc366f47f +  ~I8bbe1a2ace8f51aa22cca5d9fc66f136 +1;
assign I4b64bd561b279a17da4758a188a2f395      = If75e99660e3997f53f7b903bc366f47f +  ~I38c3e3e136acb79c8a0ff850bcc55f16 +1;
assign I93d5297fada8dfdcffed4b7b56ef9c43      = If75e99660e3997f53f7b903bc366f47f +  ~I35b2c7e9cdc53a98913e1c16a3a47b37 +1;
assign Ic6e5118343e784f89cd1d3ba03309f20      = If75e99660e3997f53f7b903bc366f47f +  ~Ib1a2b31d49ae476e2f1fb9acba2d5af0 +1;
assign Ic5d76ee2f693c012e26dc17acb0086e2      = If75e99660e3997f53f7b903bc366f47f +  ~Ic72f41f9bbf470aee3c9b9b8787b31c3 +1;
assign Id4ad545c42b5e4c8d5383568ad1e2013      = If75e99660e3997f53f7b903bc366f47f +  ~I3ea4c33a9419820ed54460eb64134dff +1;
assign I3a6030885679b87e44a54cdac13681ad      = If75e99660e3997f53f7b903bc366f47f +  ~Ia0d940e16c8cbd4f7544f5a5cd7d83b2 +1;
assign I0791083d118ca9bf64108ec397af3d04      = If75e99660e3997f53f7b903bc366f47f +  ~I4a8abfa0896ce414d9b98093ef84455f +1;
assign Ic683598c8ec40f18eed02cb89e8a8270      = If75e99660e3997f53f7b903bc366f47f +  ~I680be647bf2a62e0ee9b5d379dc87b4f +1;
assign I1fc9bb5cc8d38dd67592141a4dbf2532      = If75e99660e3997f53f7b903bc366f47f +  ~If4d75f83299a21802b6fbe136913489f +1;
assign I7ec34dc5c899abcd284ccd637fccf4ba      = If75e99660e3997f53f7b903bc366f47f +  ~Ibddfda6413e3dd2f483c3174ea836b6a +1;
assign I2d43f4939c3509b6e7e540d3da880c35      = If75e99660e3997f53f7b903bc366f47f +  ~I33bddb0adcc2af7b12a83bf843036385 +1;
assign I385df2a645f7269a298cbadc418a54b9      = If75e99660e3997f53f7b903bc366f47f +  ~I529f92b82248efe2cf64f7da0ec8283c +1;
assign I5f90162de7034f414b502958f5ec9b3a      = If75e99660e3997f53f7b903bc366f47f +  ~I2f34af0036985cd94ade9cc905bec065 +1;
assign I74353ed1bcc55b22f5d1f406b5069eaa      = If75e99660e3997f53f7b903bc366f47f +  ~Ia1a0d8d7dfd6e877f15cce773f85f5b7 +1;
assign I6c28ab1bc42131e4ff3fa98c97990c37      = If75e99660e3997f53f7b903bc366f47f +  ~I5dd29fd1a73df5662d2b636e7285bad9 +1;
assign Ia7c2ca9384d0415bbfe92f719a8a4a2f      = If75e99660e3997f53f7b903bc366f47f +  ~Ide530e6f4622c8a7b101b6dce9650e42 +1;
assign Ice3a20a00f8742bbf47a043b84964ee3      = If75e99660e3997f53f7b903bc366f47f +  ~Ibaf00a6780325882067a79f0c4d693d2 +1;
assign I22bdaa7e1b37f335d3fb2232df587cfd      = If75e99660e3997f53f7b903bc366f47f +  ~I16e3559c63ebfed83d6698fc9a9cd93a +1;
assign I1c41347158d76f8b81dfa334e99d07ed      = If75e99660e3997f53f7b903bc366f47f +  ~I9747a02384abb1c2dd1f52b3a5a999cc +1;
assign I3464039cbf8ed089ae1894998c1e156b      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Iceb7a1d4c23806b8f5824016779ad129 +1;
assign Ie7409851212f99a429d94460669686b8      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I40ef50004a60ae58aedc49eb5e6797c9 +1;
assign Ia575bcac8f127884a151a3a323763614      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I753f92da60980736440aba814a156f1e +1;
assign I2a193624be6cb259f18ece3546c7ad21      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I4ac79b67a8904b95f7912d24af420585 +1;
assign If40ad1197633c486c3aadfa277f9ab51      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Iad44c932cfa5c249c5e59f8c706173a8 +1;
assign I629ddfee3e7d36b93b743e69b4c817d6      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I10f14b6433498e3b9e9bf021b60115e8 +1;
assign I3469ef81705fd1534d6e5eb194f1e4b4      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I96008f47b9f134c9c4274cfcfb28e550 +1;
assign I832d0a2832b2c665f1261b07ac6f9f2f      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Id0344146d1a53d418add6d2b185377dd +1;
assign I3c2aa289ff967b044d6a37f75f048ec8      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I1eede74f12d37331b399eb7136bc621f +1;
assign Id2ea09c8febd9e18d231a5b069beb3cf      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I3e4754acc31d99bc71525789bdee0c1a +1;
assign I7b80623d743adcc50430ab9c8591ff29      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I11c1fc94a3bd6dffa17e1571cc6ae97c +1;
assign I05750cd7c98f3c9726b8bbf5cdc76844      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I5395ee57418c31e11cf847f0f514ec19 +1;
assign I389c717754a30812dc8ae3c8dffa20fb      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Iff125392fa39afebae1637a19c4e23ec +1;
assign I8f151f04b124fa5023d7be59c9a43519      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Ia6308e16fae5428f4ab6560f5b21479a +1;
assign I29a6f7a5b1c0bcc988363bee48b6cdc9      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I5ea02b5349cd4d99ccbcb6b26f0cfdd7 +1;
assign If35ed918a1a2b59c5e0ba5f3e0a1a6f0      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I21de4f6194dec9e3c401934db92c25e7 +1;
assign I0816b1444f89b9c61ccfee1d16a72c1a      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I57d0920119f8901bd4dea2d5f8fb5d90 +1;
assign I4a292e7bcef3cdaa716ceb101685471e      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I89537301987d6da0dbe6cff3caab3ff4 +1;
assign I1d6b3fdfa7d64dc0761ebcb6ad076bff      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Iaf0bbbe791bb71d0f557dc71caa5fb87 +1;
assign I3ce8fb414e9fa103854658db43291eb0      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Ic7ff9cde71054c1ee9eef81eabdd7061 +1;
assign I01d190427900b3cef55d978630d6e035      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~I88c10c47ae424fbdcb852fbf1e94127c +1;
assign I59a613f178a100a88f479d85e5f01cbf      = I3253481bee7dbfc0f3eac94c3252ee4e +  ~Icd2e75e47cab1d539ba9ff1b6e1d7155 +1;
assign Ife0377dc8109d89213ab27df5304e1e0      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I37e6bc7aff363ed0ed1f84b23c5f3e34 +1;
assign Idb55c5acb92ff1b590670da114d3c668      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I733605337bf6972630c089d32fd7f98f +1;
assign Iefdc7b1d3aea42c3ddf9645510803a98      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Idcb1d8bbdeaed6768c2a418c3048e6ee +1;
assign Ieae82f715fb1dc2d6d173f82b1547c35      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ia89da2f1890524ad3519ab403dd0686c +1;
assign I18a9e19a2c41be29621e5da6a2b08e3e      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ie33a780b0221084898c9fc5b237b244a +1;
assign If4bfa23dd5ba282c7c9445769eb865f2      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Iabbd1668e0014df518ede5216232834c +1;
assign Id9717e06ce4a9b03b8430559671918d7      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ibd89458312687610aa166a9538968851 +1;
assign Ie54acd665004eec584ab9ff50df3961c      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Icbaf92a8e9875bcb19a1d074779a9ea5 +1;
assign I16c418af5cc92780b28cd56e8baa825a      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I80f3c8559da8e97bc5397bb8b621a0bd +1;
assign Iddb359180e3925dcf7081ba0560c27da      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I7a0eada108891aba06cecab5071232c9 +1;
assign I354ac9e0f361928cf5cc7aaf22fd9622      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ie21a2c9b22e7bf8425fb5c0f33e5f4f7 +1;
assign Ibf2b259738d54319e3af570db254a79f      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Iaa5b2807e5cc2403c5787eeb3d10ca6b +1;
assign I07150b2eb1a5818fe98aa210cb6e8221      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I6da2b3a481ee71b85f3087b36b399288 +1;
assign I5dea5fdbd4e09be8fd264360ae399b32      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I11094e852295755925c3c61f1df81643 +1;
assign I9c52550c142c131371199bbf8bc08c01      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I9c633aa620cca127b0ff8cf882178e76 +1;
assign I72d86068a1d9bdfe04f6ebe9afcf980f      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I694d471fd353eb54aae08a2afa7b645a +1;
assign I412dfb474dbd41f407bbd57b0dd75a4e      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I816704585ad393f685731104ad3ec64f +1;
assign Ie759523643b0c4becb96025e66635b3b      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I85d95015a9ce27a18ccbf73bbbcdbd70 +1;
assign I1ef0aa04ba8b896c7ca95c10513b0ecf      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I992e7c551b4aa818606c3465d33eb798 +1;
assign I880964445bdadb87455b7f8a865fa0e8      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I2ead0e9941e2280309ab53535b1e1ac1 +1;
assign I145bec82b2f3234d2299ea32c9cd32ef      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~I56873feb8418005b5661c7382f2dbeec +1;
assign Ib045b4ad82a55c17dd36f29467d49f36      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Ib6ea4a822da2ea32e0abf6cf8a33d295 +1;
assign I7a195d3fb06596483191024720bfae2c      = Ia80693da8182ee2c3708b6ec21d397d2 +  ~Id1659ccdeaea3e59eb2d3f65a65ebd05 +1;
assign Ib84c4b8d94ce1e35ab220224ffedf4e5      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ic2171967791a0329f3e39fc19d0a6bc8 +1;
assign Idd54eedf955c30f097484bd789eaa3d1      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I7d5041a6796c00188f74936d283defe6 +1;
assign I123677fa899ce173a83101d91990014a      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Iba7608ee0a01af103e022bcaf564bf6b +1;
assign I26617d3c93a1f4069ee6fb732264d935      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Iedbe9d0e48bd36064f59faea51afddb9 +1;
assign I00410cf0d9a85b1fa2f70212bed15642      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ic3871325d57b310c95ca02fcaca529eb +1;
assign I28f355e643584a4ab8d55777aa26fa78      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I42f9b1f8ef24ad56c10086852678b456 +1;
assign Id21bc865cd2de83bced952fb9c25f11a      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I3ed5d0fca86f35b3d4b4a89c6147d0cd +1;
assign Ib6fbb4e2ef502ae86dc697dccfe035a8      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ib0126fb335e32793c400a97c5a4a337c +1;
assign I2b0c304769c917cc6acc0855ada30c54      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I20590d8fb97ec0b2164ffe17826136a7 +1;
assign Iba61bc5c2e1230784d619375b7c756b4      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I3c128efc9f80c9b8334bf7b61de71b43 +1;
assign I613acad8a236e9deeb6967de9c067a48      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ic7147944f8835e26b9838fdbdc18ca41 +1;
assign I427eb014c821ba5108aaa6ebbd8bc23c      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I698b1dbc9d8664d1c86c7a763d97b3b7 +1;
assign I9b3fc0250b26e6faa2b7b44e863ff3f0      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I508bbade361787127e1a2e8687ec884c +1;
assign I79c12183f8bb94f4a3ce466570eadb80      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I2afeb2a7b199c0c6738938f156ae4274 +1;
assign Id4ba2f12931de7439cd52eb15b0241eb      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I86255756ddd1f88b74e070b19f8c3bfa +1;
assign I430558329b5398ffd51855414df8ba17      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I7d4924388dc5373ad7936dca76797473 +1;
assign I4eacf5b6fddf6cb1dad592392eeef166      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Ie317e5ea2ca4ba2060d0f491290af96f +1;
assign I64921a58b87a14a3d6d02647f5c4a496      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I56ea52c50a188ec47e48740839a031c9 +1;
assign I9a93abf3585f9f937118adfdacdd8736      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~Id9b9a8fe43992ec0793845715dd2226c +1;
assign Ib368c9afabdccf356ff389540397e3e9      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I93b69bfb228db4b569a6772179d603be +1;
assign I939d31990dc2265d78b3d5b9a031f0df      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I71afab29cdb962e1f1ca21b61dfb50c6 +1;
assign I3ded8a67a0163feb95cafacb2c539412      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I9905e2686b350e8a6e7f790563a91294 +1;
assign I20c10afd04ed128ce31162ca3c1a89fa      = I7fa3f2648baacebf9e4b59c179601fa6 +  ~I524e78ae6a4204e17ba4532dba047d4b +1;
assign I71db9043fb2adee1e96818330469e51d      = Id7699f8f89380c315303644fdebacb32 +  ~I71228fe4188ab1d9796081184a422094 +1;
assign I64112bb2686f6348b7caaf3e0cf6a4aa      = Id7699f8f89380c315303644fdebacb32 +  ~Ie19b39200436b0bfca13502ad36c21b9 +1;
assign Ib4d8b49de697e1a70b07e76e836872b5      = Id7699f8f89380c315303644fdebacb32 +  ~If6657f90c84ca5e2ba08ec705f34be03 +1;
assign I67dd716c2039d45a57fe94847cf2eef5      = Id7699f8f89380c315303644fdebacb32 +  ~I60ec7459bbe99fce295406bee1f2af46 +1;
assign I60558c2a8261a6c4a06491a95c40dfec      = Id7699f8f89380c315303644fdebacb32 +  ~I29ab844f80c105d247c5c15faa35863c +1;
assign I37e4ed1440968cf86567341f4febf6a7      = Id7699f8f89380c315303644fdebacb32 +  ~I856fa68463aa5ef1ae53442699d38b33 +1;
assign I369a541788e6ec2dbf5a29a93b8e9379      = Id7699f8f89380c315303644fdebacb32 +  ~Ic3d00a27f15f8983a120395082854d6b +1;
assign I7fcf3847a6884d9e2cb216ac22cc6eea      = Id7699f8f89380c315303644fdebacb32 +  ~I6b1d01c3cb8fb51e43cdb788b89816be +1;
assign Ifc34e5240f1440c3a0415cc944241208      = Id7699f8f89380c315303644fdebacb32 +  ~Ib74a56900c1f8b159ad381f61acee801 +1;
assign I7e7a9c6ba8c0e7b945fc5cbc7def9c6b      = Id7699f8f89380c315303644fdebacb32 +  ~Ia5eba52d169755c507b9e0094e467fab +1;
assign I8ea9c190206ea186295c33528d45551c      = Id7699f8f89380c315303644fdebacb32 +  ~I0899e8fec1a7209cd94757c0b2f87c9a +1;
assign I70f9d851136c9e8fb264fb43d6ebeb61      = Id7699f8f89380c315303644fdebacb32 +  ~I08ece7cd684e593e02321612b7a88cee +1;
assign Iea50b0ab0e00bfce47e6fdb129ea4cae      = Id7699f8f89380c315303644fdebacb32 +  ~I691c84d81c60a462e28e2b2bae3ea845 +1;
assign Ie74b8877e9a7df32f3f5674aab1300af      = Id7699f8f89380c315303644fdebacb32 +  ~I58dc9cce6384160c0a85c6efb3319cdb +1;
assign Iaa3d8acf714f23e5059aa21cc1c36dd4      = Id7699f8f89380c315303644fdebacb32 +  ~I56bf74b5890ec67090f499afdc0a9c88 +1;
assign Ic98698807ac6942eaa491de5a2a523c0      = Id7699f8f89380c315303644fdebacb32 +  ~Ibaf2f1f8bda2f6b932dc30f8369c0e1f +1;
assign I3579622172c0ccdf3eeb3bd490b2e6db      = Id7699f8f89380c315303644fdebacb32 +  ~Id9364a29fd79b52d0442e18dc0227854 +1;
assign I1369d79bd170cc9b7ed0352e0701261b      = Id7699f8f89380c315303644fdebacb32 +  ~Ica3a41ace27f7d94377981079952f4f7 +1;
assign I16196f7cfe21843797e1f3ef19b09048      = Id7699f8f89380c315303644fdebacb32 +  ~Ib57795a63d642a73456324bab41384b6 +1;
assign I20e403ad09d5eeb59020f7fe3b683432      = Id7699f8f89380c315303644fdebacb32 +  ~Iabf572c97b48c6a7dcc19e56676e3a82 +1;
assign I8d6ef29e41c3ef0fe66820e77c486591      = Id7699f8f89380c315303644fdebacb32 +  ~Iefd370d0df1a93639af482f78a1e8706 +1;
assign I77fcee77b0cb1c65ca313526461231e4      = Id7699f8f89380c315303644fdebacb32 +  ~I995d2809ffaf0ecda6a004d01cb9c8c4 +1;
assign I40c64a3c54b15800ed725dfce5144f17      = Id7699f8f89380c315303644fdebacb32 +  ~I4e8ebc46bc068c3f9889d970db131112 +1;
assign I57bddc5d3b9daf16fa9c2eaa3a148a03      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I7b561638da1b4a45ff59be81243e4471 +1;
assign I5d3dc544f4e02f31e8dbc2b399afa89e      = Ibf3e1ead3776901898d4b154aeb61267 +  ~If0a3b88a66a816b25f17ced5d0e8f775 +1;
assign I0bc53eebdddc25c9c1423068bbe7a2a1      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I0374ada4fe50717f2158468b7ad205d4 +1;
assign I23429a89ac40e62e5b13ec75e348e432      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I357137b41bb91e0659b1ac6ead9b5c12 +1;
assign I417ae67e3ed05fb6ac8b24bcba692a83      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I5d70bc64cf7b3d3ef4180e082e533237 +1;
assign I5edf732eb5451f0f84087b8ccccab387      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I7d9ad929660cd212387d893266b681da +1;
assign I26833c93cc1b8be86febb45560ae4707      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I34be4b353cf75603301372840c2f91c2 +1;
assign Iab7fe9d9176e8ceb00b7d04116dc0236      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I14834fc8e6489775359bcecf5a37ff4d +1;
assign Ie66e4f53df7e0bb44442a3c74883ab30      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I633a74e4dfa841c9fd13dbb6564c8493 +1;
assign I591dd226d239200c681a1aac16849d31      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I157bd468200e63385583b9045758d81e +1;
assign Ic572d19feb1b9d45cb81aa0aeee01340      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I918c46173eebc5b2a95e041cfd91d958 +1;
assign I31306ed55c012f4e3f3da72bc404d6ba      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I4f8792c18bd07b23e82bbc44b4ca947f +1;
assign I374c888e91b747a2a6b58649c4a1969b      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I8d0a1ae4c47edf1f2b99d1175aaa7197 +1;
assign Ic71fea427a788b416d088a44f2600c51      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I734e601f5f9d568a44a48834559e04db +1;
assign Ib6fec22f8466773bb13224a90a4e3c2d      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ie421da1dc5aaea57c50d0c7d9c5a2717 +1;
assign Id30dc8c00fd07e9ad68a8fc3c740557f      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ief5cbddfbfb98fce4812a676849b9a98 +1;
assign I85777d4d61b8e6fc99706bbe7fbfad8c      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Id113cab2dd1949d32e3c1c15273185c8 +1;
assign I707e0745e78aef8c802c0fd5a7b58ae5      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Icfe1a689e33b2b9aa9dba692d6d610b9 +1;
assign I513c23daa981e69789b074975a589954      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ia4b671f3360f3ce55db0dc0e4d78ddbe +1;
assign I3b0ea0ad1bf5f5820e582b0c1f97d949      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I60cbd4369e7ba9b6532f279e5c59084c +1;
assign I857759675a04284a230c6e09e993db26      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ifb6c65a00d9a2c31d8b1119b949828d8 +1;
assign I943326eaa918c39cb3fe412c77d8b131      = Ibf3e1ead3776901898d4b154aeb61267 +  ~I4a777f0dd62b19dd340ad31517c4e789 +1;
assign I9dcf55a3343d214ab70cbde50a34da4d      = Ibf3e1ead3776901898d4b154aeb61267 +  ~Ib75747cb32130d44b338ed8c8af8ca11 +1;
assign I1fe6a30dcbcbdcfc0b3d6bbe38e9c3bc      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ic7e35cf8d5cd230b94c40714f16e2418 +1;
assign I39216b818931b9d2fb6a93e5eda743aa      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ic51bb9184dfd103703cd0c6ad6edff4b +1;
assign I24238e5bba0bf63288ad44c5dd3545f3      = Ie486617fc1d6354c7f347692cdbd894d +  ~I103f1449c78c47396d6a54dc1c810934 +1;
assign Ic0a34c6b56cc30ddec7e5b755e18a27d      = Ie486617fc1d6354c7f347692cdbd894d +  ~I56b3a97dc3037f0bb2eed93a9482c813 +1;
assign I45e63318c784a30395ca1bbc692d1402      = Ie486617fc1d6354c7f347692cdbd894d +  ~I51e98035b35a35fdc52f5bab8f19c152 +1;
assign Iae0e9a6d88b4fba34944cd2f0dd5c9ed      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ia6a7f9beaceb08d81012f0e72171252f +1;
assign I91d8bc9088850978c17bfa5f0bf93b26      = Ie486617fc1d6354c7f347692cdbd894d +  ~I21b062856ced09cb9131c01b5e166f32 +1;
assign I014cecda30cbc4e25a1265a65ed0f0d4      = Ie486617fc1d6354c7f347692cdbd894d +  ~I4f1221ce7880729fe584b42ef3afe6b2 +1;
assign I845250d1ee6395d022a0a20698eea330      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ie7f3f1d6cee7f02ae1b17740ed54c049 +1;
assign I5d36a24496d96371aba3f0407c21e34d      = Ie486617fc1d6354c7f347692cdbd894d +  ~Ib196f5bcf9152703dc32c5101076600a +1;
assign If2f7a871f45dc098b3ebe056153235c7      = I7ba403c6745e7d026282ad704e065702 +  ~Ide9ef5a16d8fe32353c2c2a30e8ee3b0 +1;
assign Ib49df5d97f0ba140b6ec5f80aae719d6      = I7ba403c6745e7d026282ad704e065702 +  ~Iee6f2484a381bd42e441ff072ec582e4 +1;
assign Ib25900518732253ccc4800716f3d772d      = I7ba403c6745e7d026282ad704e065702 +  ~I53121a39de0bcba91a4d0438be2ae958 +1;
assign I9d9b410818773fca2bc21ed678683369      = I7ba403c6745e7d026282ad704e065702 +  ~Iff7950f24f0a6b0073942c37fff49d37 +1;
assign Ia003b700205a0b2faf1cefa2c85c4df0      = I7ba403c6745e7d026282ad704e065702 +  ~Ide86f019e9573706c25bd8b4552396a8 +1;
assign I3b98b4efc159ac3eb3c7ea322459b666      = I7ba403c6745e7d026282ad704e065702 +  ~I2370042234b0e93bb66e44b97fca3e43 +1;
assign Ibfe30b79869ff3125c248f623c494d09      = I7ba403c6745e7d026282ad704e065702 +  ~If9efe7a1c359ec03014a52870ac13aec +1;
assign Ice88c3ab21612bbd46676c650d9f4dbc      = I7ba403c6745e7d026282ad704e065702 +  ~I6a6eb62960b616043415406ebfc21346 +1;
assign Ideadf767ef2ab66a1495ead1806ffe47      = I7ba403c6745e7d026282ad704e065702 +  ~I06c7728ef64be8311f48d10d766d0c44 +1;
assign I28749b0f4f83f99b9082f7004e72aa70      = I7ba403c6745e7d026282ad704e065702 +  ~I9fe11f6c8147391aa4a5afd1a4e4f731 +1;
assign I71ef3d84207d8995c13e88c16a0bacf8      = I93cb3974b8594665b2e7ce5593fde69b +  ~Id50edc56fce48130247fdbc42eeff9ea +1;
assign I630979d7924b3c17fe0aeaa04507ed03      = I93cb3974b8594665b2e7ce5593fde69b +  ~If3e5161254eb9056914c46263b865c10 +1;
assign I50a84fa93d73bfe0287f3297707b1901      = I93cb3974b8594665b2e7ce5593fde69b +  ~I58703e8b6d04f8c69ac38f5fcfdc4efc +1;
assign I19d6383f6319e9ed4b4f16fdf7a40cef      = I93cb3974b8594665b2e7ce5593fde69b +  ~Ie1f41720e296ced1b74cb325b666d88f +1;
assign I3515fa4f304e4b1537c612ca0212b4bc      = I93cb3974b8594665b2e7ce5593fde69b +  ~I5d5701435c96f1078e741921b56e3c65 +1;
assign Ia154b83a5a01bf0ea74fcc873e45d980      = I93cb3974b8594665b2e7ce5593fde69b +  ~Id96e744d9b10dcddd1ae0115ea57a76a +1;
assign If021572d95ea7fcbae1454447dbbe212      = I93cb3974b8594665b2e7ce5593fde69b +  ~I0c0060fe260afa3cdc72f35ffb6938ff +1;
assign Ib6c860f3146839d2c0e925007ac02d67      = I93cb3974b8594665b2e7ce5593fde69b +  ~Iaec1f186cb4a65da21d41e637fc628f7 +1;
assign I21ae48e98044dcc69386800f72cc5fb7      = I93cb3974b8594665b2e7ce5593fde69b +  ~I9c15a6a5c0db11ede80ff6d04c9a56d8 +1;
assign I4f436764c02c61027d89854865770734      = I93cb3974b8594665b2e7ce5593fde69b +  ~I8922487573e02d684a3d71448c3828f5 +1;
assign If213a0715834eb56c9c8862dcd643f36      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I47f17afcd5871fc3ac378316fd3d7ae9 +1;
assign If1eced44ede97a4e0ec55c26df8d6935      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~Ia9642d79bb50567348083b4435c7d66d +1;
assign Ibe579be01c1b2925be397ab7d202c200      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I2b2bd845428c49346ef8e94e95b618f8 +1;
assign I675731b8fceb36c9a103803dea3700bc      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~Ib730fdb59198f23d1e590f6d6039e96a +1;
assign I01374171f18d419d149433d7c789f1ef      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I644e83f0a7d432fba38ffb2d99088eca +1;
assign I9f66291cd8f80896cf27fa0b8382f465      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I97f2b15ce0a74e68d5a4438111adcb0a +1;
assign I73341b7d2d30f5fe7ce2d8659331de3b      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I84c88b631bed5311cb6e99e58941149e +1;
assign Ieb9c6cc947f6e0429770118119be79e1      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I45c5e6710240685bf54b73b0d7a64271 +1;
assign I2c58e39ab3b79963fa0eddc7180070dc      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I5827bc87b5db1801b7db16e1e61515db +1;
assign I789b342281d9ed8dbc03af5c0c508062      = Id6a9ab06d58c3a01e1fe04fcf61406fd +  ~I1c85c8f73ef80a6808c6aec0c8eca8ab +1;
assign I95b62a2fcb0af75048d095dde733ddbc      = I261bd53528b82128acabd405389c8d60 +  ~Id13c99b7f7500c8195b54627efbc4232 +1;
assign I1e9d61b53dd7ce47230b341cc1b4e8b4      = I261bd53528b82128acabd405389c8d60 +  ~I4636821315d702a677dc93113872e647 +1;
assign If5d6db7c002ad813677ca165380839b0      = I261bd53528b82128acabd405389c8d60 +  ~I9c981b0614a29386ca5e8ebc06a17f15 +1;
assign I0f7ceff0b6160697dbd097293de15156      = I261bd53528b82128acabd405389c8d60 +  ~I4df3d4dac24877b14e6d361bafc1a800 +1;
assign I2e142efe8de226e1a283576d1ae9ced9      = I261bd53528b82128acabd405389c8d60 +  ~I913d818403024510c55b65b56a38dd89 +1;
assign I88e4b172c1b5c2733bf050fa442964ce      = If7fa833bf1b1438e7a5bc783ee745252 +  ~I57015930f5b09a6c6b030ed01dad2177 +1;
assign Ie1f997dc210ff90c7ff78737d1240c30      = If7fa833bf1b1438e7a5bc783ee745252 +  ~Ib54d55a70605119e37e9898b940ff636 +1;
assign I31307a02f9909905fd672eeaf54422a6      = If7fa833bf1b1438e7a5bc783ee745252 +  ~If7e146da4f3bd255b8457fd6902005f6 +1;
assign I1e2dbb3cd67d96f046b39fd52947ff4e      = If7fa833bf1b1438e7a5bc783ee745252 +  ~Ied00d87af99ae55144fdde41ebfc1357 +1;
assign Icad3b8650e3c4b3a425e1a1c7da14c1a      = If7fa833bf1b1438e7a5bc783ee745252 +  ~I7774313f1ae5a2de98855aad572b3676 +1;
assign I40acfb6473e56562b5bc1e7bfdeed8a6      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~I679baea452c3c6d04c53baa88edd8eb3 +1;
assign I06a6d7c6a5be68cb75d83b2d8a1d3217      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~If4132b39ddb92aa02d8d0346fb0e6691 +1;
assign I3d3ebea1cf84cec93ff60459177fdd18      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~Iba70e737d52e6812a67c159520e5192f +1;
assign I59868ed1411b6439564cc73edf55297d      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~Ib9ceb8315f0cd848f861bab677c2c694 +1;
assign I97ae3d6c75edf1fd87347a8fd50fd27d      = Ibb103853fc21f8f3d466ca16557ccd3e +  ~I7846bc2cc11e08d05f7c853c4920d555 +1;
assign If98ad7df6cb49466733052834b458bb1      = I37446eb66ccfd268cb418655b8160fe1 +  ~I0865623d3350645e63fa6e6c9b78ac57 +1;
assign I2ea63dcc06519b46da5b70cf36b68c76      = I37446eb66ccfd268cb418655b8160fe1 +  ~I0262b30a4efa9f1cfb11d1c3940de9e7 +1;
assign I979c3adad47ed2b8488aa7beaab7a565      = I37446eb66ccfd268cb418655b8160fe1 +  ~I7a2e79d42779ad235bca6ce3757cf588 +1;
assign Idc93f47a3946c69fc0c956ec3e4d4c28      = I37446eb66ccfd268cb418655b8160fe1 +  ~I09e9a3cd4c12d204f760758e873a177b +1;
assign I3d57c80540bbdb043ce47c688950fd18      = I37446eb66ccfd268cb418655b8160fe1 +  ~I30b0b1d54912c1a41a02a25ab238bb54 +1;
assign Id2083cbcf2aaa813c72071314c13ae6f      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~I49fb0909ddf66fc0073e6400f1a07844 +1;
assign Iea95f61532bffc857f39331b244188d0      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~I9938397dc94002481984f5b560fadc58 +1;
assign I42dd514d52d448707c7dcc5c799ee7f1      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~I4378d139db4b710e3587aa72df22b70d +1;
assign Ib6ee76ae9fed974530f73fb401405e27      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~Ifa43d74fa91b7b9884969f575ef9ca8e +1;
assign I3aea3d7d9965e4cde24ba83120af804e      = Id17f6250f8c7f1d7f75fd27f92698da3 +  ~I7c19a79f441ecbb73685db5a505e7479 +1;
assign I3b1550f5b3e421d44005a01b0075bf33      = I9957b02e8d0d888e6950eb553d9084d7 +  ~If2af8106efc1f7dd02c074af68278b3d +1;
assign I00bc9cf3ab66e198dd7bf2cc930aa2c5      = I9957b02e8d0d888e6950eb553d9084d7 +  ~I89a3f8d5f760d1a650f85814cbfdc017 +1;
assign I79d4eac1731095e588b7003d1c83aba7      = I9957b02e8d0d888e6950eb553d9084d7 +  ~Ifae345c79662c3df3dff0fe68ad68746 +1;
assign I6512194d646b949c1f8037e3911a8720      = I9957b02e8d0d888e6950eb553d9084d7 +  ~I88a61cf72347d695489909d0819332ab +1;
assign Ief2dcb1d14d5065729e66207068d0519      = I9957b02e8d0d888e6950eb553d9084d7 +  ~I9aaa036a6158d11c235bdc8406d79f4c +1;
assign Ib343818dd2f04189d56a6fc40c8da197      = Ic71258b745437bc8463fb4f847c55e27 +  ~Ie8df350430970b5f1229cda772440f85 +1;
assign Ie38501f8b5cd9e64ed80bed953adbb48      = Ic71258b745437bc8463fb4f847c55e27 +  ~I7d77ac9b64b2e8cae21c6e36947e3ca2 +1;
assign Id50a8c0b1739857f19228131b51f7937      = Ic71258b745437bc8463fb4f847c55e27 +  ~Ic1faed76fca5a9ceb7db26c2f43623d9 +1;
assign I8946d670fb58546b8854b34dad0e8430      = Ic71258b745437bc8463fb4f847c55e27 +  ~I3ca2b9b77ed8d78a10aff42a07a53b07 +1;
assign I122129edde3336f22ba613499bfabfc0      = Ic71258b745437bc8463fb4f847c55e27 +  ~I1f00849ea055a7893df386aed162a7b6 +1;
assign I2ce23daae62346911511cfea5bed788f      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~Iaf8a19fde3de660c3fa925593bebbe0c +1;
assign I5496ff29bde6957c01c5d7e5f2d8cbac      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~Icd1da43a4d95230e79dbd35a7ae41066 +1;
assign I66fe45afee3cd240ed3ef77262387f40      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~Ice9079fb6e08d629f8c0c9ce332c8f11 +1;
assign Id08a0b67ee6d6e08628238b1e5ac0dc8      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~I15fafe2baba4d2f28037023a81ce0a81 +1;
assign I2b94a5c3e2ee6f13fae5ec588be73ba0      = I24bb5c315eacf0f4e8c86f6582389e39 +  ~If4d5b48882e9e628cf51ad2ac2f38c22 +1;
assign I8b6ce93d2c7b309d4d043e938ef6cb12      = I607f203694ff76930cfee4103cb73c30 +  ~Id0eef1adba01447c14a6f005782dd9a2 +1;
assign I46d88449ca1db5f462e0442932bc5f53      = I607f203694ff76930cfee4103cb73c30 +  ~I1d1a7c5928982c278d068ebd262254da +1;
assign I402417fdf22d1b9e08e905e3206a6edc      = I607f203694ff76930cfee4103cb73c30 +  ~I6354a0e638340378124e4df7f3d145b8 +1;
assign I287e3042873300b74530542044f57277      = I607f203694ff76930cfee4103cb73c30 +  ~I0236c912c6d684bf4862b725be9d5951 +1;
assign I4c6118afff7012ebdec7b6168f1ba067      = I607f203694ff76930cfee4103cb73c30 +  ~I6f3be51d69b2b64a04e55b8946d5dd56 +1;
assign I444e2151e66af9ec6c1e984ad706b7a0      = I607f203694ff76930cfee4103cb73c30 +  ~Icde3e6dbcf985682041f30903ad95572 +1;
assign I3c800d94a189c70fb956298deb686700      = I607f203694ff76930cfee4103cb73c30 +  ~I46ee30b46020d91707689f3468f00e26 +1;
assign I0b3393ffccd4b2a9b42a68f185b074f8      = I607f203694ff76930cfee4103cb73c30 +  ~I2605f078c1a9006c93855a9a2b0cf6b9 +1;
assign Ie1996578a600cbb605703974fcd3494a      = I607f203694ff76930cfee4103cb73c30 +  ~I4d226dd2f0bfcdbea6a2e6a6613c1b64 +1;
assign Ib912bf53b3fc6753b228a488d9d25520      = I607f203694ff76930cfee4103cb73c30 +  ~I5c942076b173cf527e1be2ddb8560e84 +1;
assign I77f81eeb736f7ad4abcd88fa9b952bc0      = I607f203694ff76930cfee4103cb73c30 +  ~Ic95191bccb18e26c10e56be395ca6b1a +1;
assign Ic09db56c2b021b09e0cf4fe501f2a5ec      = I607f203694ff76930cfee4103cb73c30 +  ~Ia284f974dd8a526f31eb81ed71a06e94 +1;
assign I576cf92938eb1c168e0f9ee1b6bf0be7      = I607f203694ff76930cfee4103cb73c30 +  ~Icc93450a007cee4c0a42717ed7600528 +1;
assign Ia1d7ca394ee29ff9cc463c525fbf7947      = I607f203694ff76930cfee4103cb73c30 +  ~I9ec9f389d0489908d497487e44c6edcd +1;
assign I7fff588b55c99166b13cd816d6a5c166      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~If8a527cc7f06a9963a80a880d225d34c +1;
assign I755d06b657ce02dabc6dbb6d44e619e6      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I39ff4663007dbc89b403f3b08a69bb6c +1;
assign If86871aa91ead2d985e915f4d58408f3      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I9590eb28a81c730b83b92ef7653e71a1 +1;
assign Ie53d1075a122b58f8ee4282b91322ccc      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I2ba1acca919bddcc22a41a28d43a4e3e +1;
assign I54acee9cb56584f9876867492fabe469      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I62d8efd4227cb3dc88aa08b6585fafc8 +1;
assign Ia4e992a0d0c4f89e3bbaba81b6be3c41      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I749e987266a20840bb8a4b1a2a2fc5b0 +1;
assign I8c215a65ea37a535fc9230a0141d209f      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I7607af5d98e8070e3d15cee23cdf877e +1;
assign I564374188b8065f6a46972355d27b0a9      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I2e11a697d7f17ac30302eadb500de72d +1;
assign Ide9ea9ced1a2398876700b19dd25a080      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~Ia0886ce792e062e22d0c224158cdfb7d +1;
assign I999b0d3276b81801b5a6a5af4d98e6fc      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I6b3cd79aa87235ff174c0299b855dd3d +1;
assign I94b6767c45b74142ab2d457b5fe3b64e      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~Ie4ae993ddb776bdffec843db0def2f5c +1;
assign I2062510b4d8249d8a9b75377d4513266      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~I3ed2da9b53daac0852a06ad1acfad21b +1;
assign Iba97ce79b40d24270208680c74b41799      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~Idefa29d4d4e2a6e9147f84893520096f +1;
assign I35b405f29c891a3ccaf0b64443d114e9      = Ica8e4c56ebb37e189ca8e6b3daafdb80 +  ~Id1fbbe0594dae272856566522633bb3d +1;
assign Ib44c2f3a3916b3eaa7452f0126f934ab      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I8070a3b7d8b1a7ae90c1a2d27aed09aa +1;
assign I2f0d79178e118fb89f9504e5f75fd612      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ie88285ce2b9c71de02ebd62e8f44ca72 +1;
assign I1e5f655fd8601930d7c9307aab545391      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ica1997c6c569c1d1f45224fbaa4e6b59 +1;
assign I77691bc302dff581968daeeeaf44e9a9      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Iaf08bcaaeb15bb0c971432f7f8b16d0a +1;
assign Ic0f0982cdd813ef3da99d8534e23c9e7      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Idcb37cfc357cc088c775409fb9225b51 +1;
assign I449f136e29d92eedd2273b58bd34431c      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ic419255414995e7168afb97b051fa64f +1;
assign I0906f557008adaf488966d5aa989e6ae      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Iee6da3120d73373627b25ab7c0dedd28 +1;
assign Ic0b69b2b6f55b4613bac3aad8e864c9f      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I56fc99a22960232b305d6e683c66fcc7 +1;
assign I6ccadd50ca8d59878cf089a35319b6c0      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I0a9a09b0ab43d2a0f1d1d01e13f0333c +1;
assign Ia5aabf0fe6a5d3731b363c80a7238a14      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ibc73d07e0c97a6fcae791e04106cb082 +1;
assign I217dc03c6c19195b3c2f478b2b8b0bb8      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I224bbdf94ac86c5c376d1db4f4d4e060 +1;
assign I70c592140d0fd63e2b9b8ab9b619df9a      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I43f2b69c6b427de3095c44d4166b77cd +1;
assign I4d9ac478c0c0b7191a0ffeb3c6d7c521      = I7089386c94261e0febf3b4f7dc1aec30 +  ~I1e50c90010a3df1a8ce1cff811cc7a0c +1;
assign I8bb214c6ec5a16858101699241a1b4bb      = I7089386c94261e0febf3b4f7dc1aec30 +  ~Ie1817cbf3a80dae435a5571dfbd2f5ad +1;
assign Iff81d398838ac6181e09d95903bf57a9      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I0052d562fb3182890c8828e52d437b11 +1;
assign I710eb104c64c7eb72a55cbfc11bff827      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I1eedecb1d8ff505c75be7787199afada +1;
assign I9f2d9117540a1d6902b1a7ec3e9d5ab4      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I7ef544597a185b1de63b4ffc4a1d44c2 +1;
assign Ie3204e2e502d2c192994f3c74f1ea38f      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~Iadeedf3870f0b1eae98d0f7dbbeff04a +1;
assign I97f03a2baec02107032233e68c0b146b      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I70ae07db9b44d530be220f06401d3d3d +1;
assign I860ccc9f56a3376ea0e8137a045fe650      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I7992ea31927b4f0e268462a3b0f18c5d +1;
assign I7b00537ae91be6f2ad8be0776e29da79      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~Iadf927d18644a232ad1f1eba7db82934 +1;
assign I68413adceb35fe859824c32bb76d9906      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I2a9c673cdd7ded79e09ada38c0f47e6f +1;
assign Ib61183063f591e5845ca8ce70f598c79      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~Ia86740e870d8063f0266b68ad6d7481d +1;
assign Ia7a97e75655c4eaa8652f43c27d5ae50      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I6627bcdbaa8afb115123777abd45435b +1;
assign I0402af748fe9d48a514d23691a2cb6b8      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I96fe3eb633eff6958ac575b997460bb9 +1;
assign I5e9d62da7f6aeaa717f5a394e2531210      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~Iefdcb71f2903b11f5cb0b8857f7a1727 +1;
assign Idb3666a01522d57729513cd3f18c9798      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I2eb90278aaa54b9c8212b3b4af7c3617 +1;
assign Ifb6e917336ab665d9bfea6dcfe21bc8c      = Ia1e4f20f32f7371cb0078d6e80fe8b7e +  ~I43493f70f0336453d77caf7f27503daa +1;
assign I0adf84fd4ea2e882b59a42dad6683707      = I790cbca796af58b1726d0a4680cc164f +  ~I26a7fe395eb583258c1ac58aaaa3234a +1;
assign I1d0e0cb3903cece98c3a65f920e5ab21      = I790cbca796af58b1726d0a4680cc164f +  ~I21668ff77cf75570cae97f575cbcf644 +1;
assign I8b12d3b1f65fad05577cf25e8d7950a5      = I790cbca796af58b1726d0a4680cc164f +  ~Ie48be9e6b6fd63baa104d0a6a4561a1a +1;
assign Ifb24658924186dba2d1a85ee28fc0313      = I790cbca796af58b1726d0a4680cc164f +  ~I05370777439b01811fe7f750d2f724f4 +1;
assign I067250d29597d7c71da50f8cf557eb61      = I790cbca796af58b1726d0a4680cc164f +  ~Icdcd83341f6b5c404f91ec7e97d0550c +1;
assign Ic86c9a00eacc20772706da9399aab4ba      = I790cbca796af58b1726d0a4680cc164f +  ~Ibba4e82d1510ddc16eb4ef64893cec02 +1;
assign I8271913876a2729269e844dc4809a25f      = I790cbca796af58b1726d0a4680cc164f +  ~Ifb00ae47340bc99669c71da34cccc59e +1;
assign I3af8e500702e46e7330796cb23979266      = I0a93f095f9efb1542116a295c0db9c8b +  ~I75a4cf2948bebc58e12bb039ed273ff2 +1;
assign Ice852e353c55faedcde1922d0179b30a      = I0a93f095f9efb1542116a295c0db9c8b +  ~I5a9fdec7d7ff99fe33ad6cd8afd9e059 +1;
assign Ibb9864cd5bcd1ef1fc7bfd822db3150b      = I0a93f095f9efb1542116a295c0db9c8b +  ~I47b1695a74e4d27389b97543415dcc67 +1;
assign I13f58835ab9e6362ffddf06976c97207      = I0a93f095f9efb1542116a295c0db9c8b +  ~Ieb38fa62119a5a77c060d6634e051298 +1;
assign I35bfac2d8d88c61e93a27db564f9ecef      = I0a93f095f9efb1542116a295c0db9c8b +  ~I3459d98131faef5a5040a03847890b55 +1;
assign I7ecdf9f7726df27510f35fe6c1b5b4be      = I0a93f095f9efb1542116a295c0db9c8b +  ~Ie9b9221b2122087cd5f309570b6d31ca +1;
assign I7327385650ea109a8bb07f1c92252d28      = I0a93f095f9efb1542116a295c0db9c8b +  ~Id4451722e8e2393d627dcd0175dc9903 +1;
assign Ib5d66de65bb7bc9e1f7b3f05e4bd703b      = I989ba39f188a44475a83e65a4960d2af +  ~Ic10356f9069e3651b9c045c906e63512 +1;
assign Ifca73a480a501ea2636c47e487987167      = I989ba39f188a44475a83e65a4960d2af +  ~Ic3a431f39c678b7175ed30fde1fa6424 +1;
assign I75a3f16cb4ddc4b0478fb1c07c10aba8      = I989ba39f188a44475a83e65a4960d2af +  ~Ib01cfd833a63500e03333f263805db3d +1;
assign I5603979fb76ebb2bab9a8764c4833b52      = I989ba39f188a44475a83e65a4960d2af +  ~I0b7b4c0a8503c751229edfe0237cc903 +1;
assign I939430bcba9f8bb28f5782040a4c76e7      = I989ba39f188a44475a83e65a4960d2af +  ~Iace01234164c8a9f7c98eeb83268745b +1;
assign I71ed74fcff44b1a6ec1ddf7b18cf8a31      = I989ba39f188a44475a83e65a4960d2af +  ~Iace8b3b3a4c16763132b5aaa6b24212d +1;
assign Icc204071ef0dd850f42840be901a1c8c      = I989ba39f188a44475a83e65a4960d2af +  ~I80a89644e278e96b1cd1c4b7f764dc34 +1;
assign Ie8187be889aa7f205231e2e60cb827e3      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~Ia92d2276a8a23521ad1b88df7c27bc2e +1;
assign I18c57ba0c68acdec8308c2ba40482668      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~I39bbec42c442d1e8c818f46ad9c096a8 +1;
assign If45f0a6203e1a6ef6e0d86ccccab3920      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~I88f1b5c12759a5efb2d2ded8483c9ed2 +1;
assign I834626bbcdd99143f36052aa6e77de49      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~Iaf4ae293c576af16f5f43a8b86c1aa3d +1;
assign I58860aa281debf67db1369b2e22b9f5b      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~I68b575fcbc5321d4d26a22bcdbb506f6 +1;
assign I885d19716778193c3288c8322cfd32ae      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~Idf600b93ee1018ecf969ed7944b6bc7b +1;
assign I19a6d51c460b600130966b5be281d23e      = I9bcc1d9b3dd258fa7b6042f0185d48cb +  ~I1cd93172cf5996bc870063aa642188a2 +1;
assign I7a4326b2355162700b8647861c80f43f      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I4af080cb4e5cc525db95e5f401019e8c +1;
assign I40ce63d36b1aa901d29c0ecc3ad20a66      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I6fc8044eb226a14ff1a786ddc96d2414 +1;
assign I32230b8893dd9fd1da4ce1f2553b5550      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I27fd0073dbcdee599fbe85cf48806efc +1;
assign If7fb4fa70b6803a7e4c64a834669dbfa      = I9ba14715d9f33ef45681ad52f5be9593 +  ~Iaee6d725a8b2653eeac6d5acb91f8f36 +1;
assign Iaf1e5c8b7267eca64468227734dcfbdb      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I4afdeba4fc2a12a6cbe3567a519367fc +1;
assign I5ab38b4a054c50fced80e9323f4a9ddf      = I9ba14715d9f33ef45681ad52f5be9593 +  ~Ib42816335dd8475dcc78662c4c0786c1 +1;
assign I779f57a085e170d2ab7e7b5f046e42e6      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I343c9efe71164c01e9c7d599e032864a +1;
assign I120e630331e23d75054584a44aafaf63      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I108c269ceec4adcff9afeda01101b838 +1;
assign I3f690a6c75649328d7cccf08cc6ca81b      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I761983331fb6e3c6c437b3f1660f0b6b +1;
assign I2105fce588dc6840254a1eaf02b549c9      = I9ba14715d9f33ef45681ad52f5be9593 +  ~I70d32affde22f9dcb2d77430fca39069 +1;
assign Ic0b28cd43f561513b63ff20e31038f37      = I9ba14715d9f33ef45681ad52f5be9593 +  ~Ic08e85346f61da036a15345a13ac12f0 +1;
assign Ib4e0926a64eaefff0e36fdde4783e923      = I9ba14715d9f33ef45681ad52f5be9593 +  ~If5dfdadb3868ed5a495007362f7db648 +1;
assign Ieb485d7a868decbc901fad618f56412a      = I9ba14715d9f33ef45681ad52f5be9593 +  ~Ia1ee5579358b564de06c08ca418a9bf4 +1;
assign I71853033c5b7e4e98414209075b4d708      = I396a897f79b519f4fa02af39d0274f64 +  ~I9bb81dda8102b829441be46460eb8900 +1;
assign I37621b4bc9c88a42a47d3123465fa4d5      = I396a897f79b519f4fa02af39d0274f64 +  ~I8eef6ca0a61a21882ea28b3d63735228 +1;
assign Ied0d483617ee30ac0539009fba84a684      = I396a897f79b519f4fa02af39d0274f64 +  ~I438522d92cce6f7010246424746ca255 +1;
assign I574d31b300f16225a707bbae0918c445      = I396a897f79b519f4fa02af39d0274f64 +  ~I92496f68b44a94565af28a2c28d6fbae +1;
assign I9fef812393d8a5f87abc46add3371777      = I396a897f79b519f4fa02af39d0274f64 +  ~I66528f43f614f0edb715564eba3c77c1 +1;
assign I64a11eacbd9a28d7e65c56c38127876b      = I396a897f79b519f4fa02af39d0274f64 +  ~I8cab9fba615b94fd4bb6934325be8ab8 +1;
assign Id11f93a74e2de2ea1e27e9d2858a472f      = I396a897f79b519f4fa02af39d0274f64 +  ~I92d9fec22d36b1baac8bd78abfc1bbd5 +1;
assign Ibd0708af1cccb49fded84694d6ffd6f7      = I396a897f79b519f4fa02af39d0274f64 +  ~I4eadce87f47df6d8f0e4acd057de5a09 +1;
assign I18edce191243df3a622232f681b7e3f9      = I396a897f79b519f4fa02af39d0274f64 +  ~I73203143fe37933c16fff873c1abf512 +1;
assign Ib68ae994fc94acf008e424d8f8c8eb4b      = I396a897f79b519f4fa02af39d0274f64 +  ~Ibed2a63af723a7abf96dacf1951e5266 +1;
assign Icb6bc0221ed78051fa10967f5cce4a7f      = I396a897f79b519f4fa02af39d0274f64 +  ~Id667c80003b5541de9f84d3b8709c828 +1;
assign I3abb9a64f85be533ac16eafaf85c5ad1      = I396a897f79b519f4fa02af39d0274f64 +  ~I02cbb4255db2b21ea32140f9e9ddb36b +1;
assign If6badde34faca49e04b3dde9b11c0556      = I396a897f79b519f4fa02af39d0274f64 +  ~I65354f2069de0c25bbe7cd50fbe892aa +1;
assign I09d6aa4053f5e1280d70556ad1cc89a4      = I197c0cd576e16ee2197a28c86397f801 +  ~Ic279867ebf3055980f3d813d5dc8dec6 +1;
assign I9d1f949ca74fcf76431906a3a95d4866      = I197c0cd576e16ee2197a28c86397f801 +  ~I5c05da8a222ad5effb9815cbf3ec25f3 +1;
assign I10221054a7689d49c97a1e908e2fb44b      = I197c0cd576e16ee2197a28c86397f801 +  ~Ib8bf21f32c0e8b9cfa42a53807bfe3a3 +1;
assign I4ec67f577ac5c95d8a93f21935a4fb7f      = I197c0cd576e16ee2197a28c86397f801 +  ~I7208256bb198bfce1be71390b01bc028 +1;
assign I069f6a3e5c61b47031648ed6e7ab0330      = I197c0cd576e16ee2197a28c86397f801 +  ~I49f2a06ceb3a59773c65b19f54ff362b +1;
assign I4b15910b07c427bfb666057cf4700947      = I197c0cd576e16ee2197a28c86397f801 +  ~I86e495dc894d2aace15c1aff89798bf7 +1;
assign I5694aa90f55816a9ca217470b70f29a6      = I197c0cd576e16ee2197a28c86397f801 +  ~I0d53bb5344cabe5fa5ce3ecf7122a260 +1;
assign Ia1d3638756959bfb67f32a37c58fe190      = I197c0cd576e16ee2197a28c86397f801 +  ~Ib2f5f5fc77ea8b529f2471c54388f2d1 +1;
assign I3e81666362b0209c98c5337a74dcbfa9      = I197c0cd576e16ee2197a28c86397f801 +  ~Idcada1bfb3c0d1f2a09aab58a2071a57 +1;
assign Iaa723368e8f531ae9bf99c9b99fdf0f7      = I197c0cd576e16ee2197a28c86397f801 +  ~I814b62120953991f9da055f118967e05 +1;
assign I3713f644fba6dd9d4bb4dc3b4c91fe77      = I197c0cd576e16ee2197a28c86397f801 +  ~I123a212546a8ac394051425db4924812 +1;
assign I5a3e3131db6fdd74e5c822fde6a8f2c1      = I197c0cd576e16ee2197a28c86397f801 +  ~Ie95f1a7e0effcec0aa423dc803056a13 +1;
assign If18033df3d6ee029fdecf3323ad8d62d      = I197c0cd576e16ee2197a28c86397f801 +  ~I106deaff50b8480eac31ddbae2ec7c61 +1;
assign I7514cd65da98bd214b4e1da34ac358f1      = I094a178e55425f27ac1ff6195217396b +  ~I68528be9951f5b8805411711cd11ea59 +1;
assign Id947f3ca55c826ef94d1ac4ad2a227bf      = I094a178e55425f27ac1ff6195217396b +  ~I0f034a8f077b0ab231727b6298e366d8 +1;
assign Ia6f83033bc647143bbf5377056c7072f      = I094a178e55425f27ac1ff6195217396b +  ~If9c12f8662333fb54a45cfa1bc5da487 +1;
assign I21dd15d84c5abe8d2ac53f65236f587c      = I094a178e55425f27ac1ff6195217396b +  ~Ie1681d905517daafcc7584725cd6014c +1;
assign Ia88c70253514b080daa27d2df0aef202      = I094a178e55425f27ac1ff6195217396b +  ~I2ff3edcdb6158f1e3c9a555aeefc0850 +1;
assign I3cd11d85b17ce4c2181dfd2430ff4595      = I094a178e55425f27ac1ff6195217396b +  ~I43b380be6df7df0d354223d0a0d6d6b6 +1;
assign I9817361d029cc98d7407cf3b8b020567      = I094a178e55425f27ac1ff6195217396b +  ~I23eb1dc4d1c992f804dd04a2d823c778 +1;
assign I47a6f2033a2356ac604133d12d7e0c0e      = I094a178e55425f27ac1ff6195217396b +  ~I7f90f96c0260560ad5e6dc7448b2670a +1;
assign I3da1998324eb1853e5ec747b112095aa      = I094a178e55425f27ac1ff6195217396b +  ~I07b417cdcc99eaea3413f563e26ddc73 +1;
assign Ic729cdba5f8a3933121a0ef35da99f8c      = I094a178e55425f27ac1ff6195217396b +  ~I2f3ab9654e515a54e22e73d6c130ccc3 +1;
assign Id7542fd1fe3a099d7274f15c008f1cc5      = I094a178e55425f27ac1ff6195217396b +  ~Iebdc41368d57498a04fa73e30b10a966 +1;
assign I1a91347d29cd64af8941a3e042228a52      = I094a178e55425f27ac1ff6195217396b +  ~I5b4305bef5b4350c1d7ae143667afddd +1;
assign Ic6b16867c426103b3e53db94469de2cb      = I094a178e55425f27ac1ff6195217396b +  ~I2795d21d343b83a69146314a2407cfa2 +1;
assign I7361a720882c68965c1c28c2d6ba1dff      = I3177408f7d08b431be99297fb10586e6 +  ~Ic6386d7d8813731d612e24b715740275 +1;
assign I668a239256c66a858129b4788b0001a5      = I3177408f7d08b431be99297fb10586e6 +  ~I4c366a57920ff090a98a2cb8b9caa00b +1;
assign I73a72fba51f575f80ded2357a6b71af0      = I3177408f7d08b431be99297fb10586e6 +  ~I14cf5d43fc9864820a8a25efcc5c6d86 +1;
assign Ief9131d8e69f733c51e9f9167ad5fa4a      = I3177408f7d08b431be99297fb10586e6 +  ~I33b99994abbb5ecf8eed4de39033e4f8 +1;
assign I1e6904544c93f0f4bf403793e50dbf99      = I3177408f7d08b431be99297fb10586e6 +  ~I7c3291f0250d13ca94802b0b071a95c6 +1;
assign I74f9e6de534920d70eda17b59206a4af      = I3177408f7d08b431be99297fb10586e6 +  ~I2c926fd9d306e9ae13364e07c4b0395b +1;
assign Ied74515bab35cad5e94048a9f210b7a5      = Id4948c876d48bdbf317d32f135e645b4 +  ~Ib23edc35fa5bbfe0415fcf0861a22d9b +1;
assign If38f871a7b021ceb84cdb3010d08f667      = Id4948c876d48bdbf317d32f135e645b4 +  ~I3e0e682047f7cc36142e668828cbff1e +1;
assign I12a578d51082c42fcc5a9e769535ac0a      = Id4948c876d48bdbf317d32f135e645b4 +  ~I99fb9030e8361e57818c07511479a9b8 +1;
assign I404f31fea404e730a9c4e04bec369c1a      = Id4948c876d48bdbf317d32f135e645b4 +  ~Ic87c3d7762a18772972552162e1d1a8c +1;
assign I915d15cb464b6e78cf9939232618b14c      = Id4948c876d48bdbf317d32f135e645b4 +  ~I7e393e6c1d1bc44daaab120d55f5dd59 +1;
assign Ia8531e691cc60dcc32225eef6d8e8a2b      = Id4948c876d48bdbf317d32f135e645b4 +  ~I448f126fd3932d5065abbe7bb2d92c56 +1;
assign I5f7cd38f8b6c42a3dcc52664ea7c08a5      = Ice5ff01d4fb4583898498651a0ac0171 +  ~Ifc8c6df8904b97674f2970ebc95b523c +1;
assign If3f0f6acad563083949c5116ad78ce20      = Ice5ff01d4fb4583898498651a0ac0171 +  ~Icd0622a90782b9c451950e7ab0399567 +1;
assign I2b8c7ab8f53d7fbda984ab8760e05fd3      = Ice5ff01d4fb4583898498651a0ac0171 +  ~I6493b3c087d4685a6b3f98c73dc2ff49 +1;
assign I29d486911dcffddec336f69b981e1e50      = Ice5ff01d4fb4583898498651a0ac0171 +  ~I20c2057240417146df144b518b43d052 +1;
assign I893881a7874f85e519089559ac4604bf      = Ice5ff01d4fb4583898498651a0ac0171 +  ~Ied029d0bdea3bf134744c99426fa72dc +1;
assign I0b730d0a75cf72482ffc5b0d0267fd83      = Ice5ff01d4fb4583898498651a0ac0171 +  ~Icb82c9ff4cb58159a1c3115c6fdd5f8c +1;
assign I9beb581fcdf85cc7302da093363e3b02      = I0fb33a5ced3d15622c9aefa188052e24 +  ~Ia3450e134e4086c35acbdee1e6042396 +1;
assign I0e35fb521572c6f87dbd06a8ce213337      = I0fb33a5ced3d15622c9aefa188052e24 +  ~I5a0f27df5158309f32f0df31e8ae3ae3 +1;
assign Ia01e93b03cf0ff22e2f002f2e84eb9d2      = I0fb33a5ced3d15622c9aefa188052e24 +  ~I17d9e19854cef197fd3267618617efc3 +1;
assign I98a2d427581a73c639cbc9f4bf4c8802      = I0fb33a5ced3d15622c9aefa188052e24 +  ~I2993acb61f1abe529f8a60c94a438550 +1;
assign Ie60ba6ee53f7a01764001bc74fb90d61      = I0fb33a5ced3d15622c9aefa188052e24 +  ~Ic8be2c94235fb40f78da33179ce4873a +1;
assign I508e632bacf8c083a8376f73cec11bc6      = I0fb33a5ced3d15622c9aefa188052e24 +  ~Ib3367565e4456da15e7c2315dccdb5e4 +1;
assign I47ac3c977bbfad06ee1782b8eac6d9ec      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I15a1671def323cd294591564ae6ef8b1 +1;
assign If8537bb117e0bebd25ece101a23674c8      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~Ic512effb493a06ece58a2af155135004 +1;
assign Ica8f952cb456e825c608f2e73ec9abd7      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I2c72248cbe49ec0a0febac2437b8a6dc +1;
assign I1a332ceae6f1a640e4577c82b2bf4511      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I964e17c41a134c080e9c43412a514f3f +1;
assign I82c5b5deaae0b927c14adfa3b477c8df      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I94f1724740defe5bb7e40041d0e266a0 +1;
assign I37b08ee3258fb8359ba4c1653101e03c      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~Ic19486b6ab0373b9c0ad8f7597782d8f +1;
assign I58fa785303fe60b1f1c596420aab4b5e      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I31243de90dc2a1656ca9d5e03bdd78da +1;
assign I1ceca376c3f4cd24c22cf8672c9343ba      = I0074e1c3ca0ff903a9201ac5fe7ca841 +  ~I242a30bdc8699d8ff550b25dd53d6c59 +1;
assign Ieca948a12a0806b9fd483ace71c8b98e      = If65f587e987a51c093e8dd4df532e26c +  ~I9d15f76bb68b214057566cba4b511214 +1;
assign Icd2579fee72faaa432876ec8fa124d40      = If65f587e987a51c093e8dd4df532e26c +  ~I9cc16a00912e7dfc05fb505a9db23cd8 +1;
assign Iec4164641d5b71630d9d5aefb1ed5676      = If65f587e987a51c093e8dd4df532e26c +  ~Iacf9640cbf486411d6ceb8fe1a2fd5c9 +1;
assign Ie43841b2ee3b5369c3863417b60e5851      = If65f587e987a51c093e8dd4df532e26c +  ~I9015033ab0caf3fa41dae4de43f24a82 +1;
assign I1e7346a531973e40fb2582a68f96e383      = If65f587e987a51c093e8dd4df532e26c +  ~Ia630e59cbce82a570ae3890a6c0221e5 +1;
assign I53b62438d1bb777cf10761bf95b22718      = If65f587e987a51c093e8dd4df532e26c +  ~I4904ab14b19fa1b6befc218bc7be3842 +1;
assign I6b8a0d9d8fe6ac6fa08c495b0d0d5264      = If65f587e987a51c093e8dd4df532e26c +  ~I282d2eb4e74e034694e33273b9cb19d5 +1;
assign Ibcec436bb431239047a99c495262bf87      = If65f587e987a51c093e8dd4df532e26c +  ~I3f33901c407a87e10d86c13c83dd52eb +1;
assign Id9d1f164781aad87bbb332ef7c0b5113      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~I43f41bf07836cee48069e9890c1de2a0 +1;
assign I76a91ad2a7f0323b5874f857eb914d67      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Id88480a0a350bb5fcf01ed5fff0bbd4c +1;
assign I9aab2781bbd57dbe4381c695f130d5b7      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~I1d9b9ff357667a362f0442f19986f451 +1;
assign I11c62ef31300f66f787bb7285596b995      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Ice73589836da9028def6efb24a04dbbd +1;
assign I7e62705e1f1e7abb04ee4a94753183b4      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Idb72c046c5996fbbd80b706666ffbd92 +1;
assign Ia4d8ab77dd8598d550c4b3c57f02b328      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Ie5757e7b1647ab7d43cdbcf98cbb77fc +1;
assign I23c2886f2707bae85fe967379c105eb5      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~I6072331f838d82329a07a4ffa340c7b6 +1;
assign Idfb980ae7487145d65bdf83b97751e6f      = I33d7e77d08590f0dfb1867e741dd8b6b +  ~Idf6875955525d80dc660ce956f4a84e7 +1;
assign If7916cdab9aa2621009bc0671d985133      = I678c22563e0273403b046df4261f21cf +  ~Ia96955d9c0a8a587e0afab37c8415d8c +1;
assign I1969f6d312f67452ec24690813fc07ae      = I678c22563e0273403b046df4261f21cf +  ~Ifec374bce7f5507438f550df22d61a01 +1;
assign I6b3c96ebbba2bfe8c549caea4a266656      = I678c22563e0273403b046df4261f21cf +  ~Ief67e897e57b96e2ec200e82bbc7caeb +1;
assign I73172f8b4bcb0bdbe27a09cd7ec204e0      = I678c22563e0273403b046df4261f21cf +  ~Ide604e9bbe35cb55892a4602e18b2527 +1;
assign I96acfb8f7e6c42f616a880b3657f42a9      = I678c22563e0273403b046df4261f21cf +  ~I262f2390e77ec486ccd3a6ed05816e2d +1;
assign I5cdce64ba621df381f9efbb8b0c8e10a      = I678c22563e0273403b046df4261f21cf +  ~I280e20c20c0b4f26278b3de9b2ff84e4 +1;
assign I61389621065261b79f16e6dae7c7cdac      = I678c22563e0273403b046df4261f21cf +  ~Ib3a0307176d424a4733720416d71069d +1;
assign Ide44caca4eb1b6edc9b55c584239ff94      = I678c22563e0273403b046df4261f21cf +  ~I76060709de3ea188748849f043c59ac0 +1;
assign I892e07e7e972dd521f273519694e4ee7      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~I8be20605d26d218911e80a883a90d085 +1;
assign I43c8950bb200a93cec12c09af4a38dae      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Ieafa9d74d4a61d28ac4a913db460bf33 +1;
assign I591f0a636f176d5a398cb6ed6d67f627      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~I6fd1b4395af175eff85b3bfeef4c329b +1;
assign I8be467496bf21fa2c46fc5db2442a339      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~I39e6d3fb468aa40ea73535e81556ea65 +1;
assign Ifa0294e878bf5a4f1c6c7cfa52c46e7d      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Iae449b74e50e0907feae9e60f2329426 +1;
assign I35a8b04ecb2c6d2d7bd52a64010038ff      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Iebf769a6bdaf214c1006c55c608d4eda +1;
assign I38629158c9fc8600b05a3e32589cbeda      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Ia030c08757123aae947f86ab8bfb6d94 +1;
assign Ie20705331f5fabb4c9f720a5c6592c7d      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~I8c35c5b343b552c22000e194c517ca12 +1;
assign I425d66a6ead3859f364e20a797b0e4e2      = Icca700c12ae2e8155ca6b41e692e8a8c +  ~Ibf80bb564263ea85bd886a8617f09bb2 +1;
assign I66a2577a791bae1f31c5b99b0c3f324d      = I5ed74e81d2497681af5a0ca13fe23088 +  ~Ib8dfd9b8badef282ca00a4f793c3c868 +1;
assign I77350e171f060c2d49e50c636fab084f      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I596ad7e132f272cb196b74faa8c75aa4 +1;
assign I2101d085d5e55ef5b8247de3898a80e7      = I5ed74e81d2497681af5a0ca13fe23088 +  ~Idc629414f6d0236ce0714cfaae23f065 +1;
assign Id38879e0d52fba6818597bd60dfc2b2c      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I157fdf8775206858c08682db3039b084 +1;
assign I68081efdf01e540fe5e07643a2bc3463      = I5ed74e81d2497681af5a0ca13fe23088 +  ~Iacbb4daf5ce5c7eb1a2afe30d0cb5382 +1;
assign I2d70e6f392396c2ee505687f5a950a6f      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I4e08021c0235fafb60200aab97827a8f +1;
assign I6e6eae8e8a955b80abb7cb722a940e27      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I730634ea15ac94d241f3ad2d6393a227 +1;
assign I54cfd5f12219687ba48be0c57a979add      = I5ed74e81d2497681af5a0ca13fe23088 +  ~Iee367c535d9c39f872d2ec043e7e7b33 +1;
assign Ifda70e49dbdc4b5511961649914ecc71      = I5ed74e81d2497681af5a0ca13fe23088 +  ~I68bb1f26f878862f288c1f57049cf58b +1;
assign I0feba37f523d6c6371bd934796519c59      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Ia9b5d9ede006c56a6d83905529c77b7b +1;
assign Ibaf70dff036e0bc11df75e2a1fe4fb34      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~I1487170cb1f3370ad45efc801cefc8ab +1;
assign Ib00eb8856f044c3af325f0134d16a970      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Id88568dd34fbee42c9cb8cc15ac5c31d +1;
assign I4e89f11e414b55e9574f5c3d79dc4506      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Ia30539545e66c4cfc16828140149180a +1;
assign If25b7447f1f34072a597f70a4234a16e      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Icbfbb37bad6344005dd233b3605a784f +1;
assign I76ae0b929aefad162304529ea04b725f      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~I91a6408a11fab36a8ba3dbd3f895a803 +1;
assign Idffaf5edec0ef7b25c24f3c5e636fb75      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~I47b878f27c30f79a37e97e022307e9e9 +1;
assign Id041de10db620915a3755358fc2d9a41      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~Ie76b0739aec66f8860870e66e87a6445 +1;
assign I92ddd31add3c914ce6b0271e77cb67a0      = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f +  ~I50383e3d7c172eedfa00aa50a9faac4c +1;
assign If80ebbd3419cd9fd63a745412b7233b6      = I26010e26e22d8a2ea831e86fae34a24e +  ~Ifeaa99e03bda8ded058f98387de3d49d +1;
assign I0b67c1f8e03165404e0b76d1a05d88de      = I26010e26e22d8a2ea831e86fae34a24e +  ~I4255ac1af4367c321567c4e46b06ab25 +1;
assign If78c15d7c2dc19cef26743eccbb52e6c      = I26010e26e22d8a2ea831e86fae34a24e +  ~Ia445bdc7def7d8c1eec31ab892c25c41 +1;
assign I228c0b3c3919aaf70ea24874f314eaa5      = I26010e26e22d8a2ea831e86fae34a24e +  ~Ic3b4752136ac08e343933ccc3a4ec47c +1;
assign I986ca3b0590709588c3d9d2274a1fd34      = I26010e26e22d8a2ea831e86fae34a24e +  ~Ica6707efd6d44ba6bbb87c0593a3d828 +1;
assign I765867ea6452d51f31e96ec83f68f9df      = I26010e26e22d8a2ea831e86fae34a24e +  ~I739267bcc50c54b8a685cb3c6afc5cc1 +1;
assign I6e970e7bafbfa1866203483ed18a7db7      = I26010e26e22d8a2ea831e86fae34a24e +  ~I9160d11439c5140c0109b5190eb82e6b +1;
assign Ia31bbc3e099eb2180960917330d6b2e1      = I26010e26e22d8a2ea831e86fae34a24e +  ~I6ff7b86cd7f63f9243646f1be10b2577 +1;
assign Ibc94d96e529274004dfed98c98915827      = I26010e26e22d8a2ea831e86fae34a24e +  ~I165653ab165cfafe2b74cd441331f9e1 +1;
assign I60eb0a19c8d75780a4dae7d33ba46bd4      = I578efe5c2c504f12c8f2466a7f734215 +  ~I08a8cd6965c23af6650568b654831b20 +1;
assign I701ff10dac46e4482b3bcaa387c9a725      = I578efe5c2c504f12c8f2466a7f734215 +  ~I9b6a674dbcbfcf65f1ae0deb8fc3566d +1;
assign Ifd170f2b9fa5df9a7d0817307b5586a2      = I578efe5c2c504f12c8f2466a7f734215 +  ~Ie3a336de822ac7baf8486b1618ef1126 +1;
assign Ia5feb8ce451f12382cb66853e948047d      = I578efe5c2c504f12c8f2466a7f734215 +  ~I5fc3c26d6c5aa893dfd5caa0f677233a +1;
assign I3a971f30fe10de02e604402b55c181da      = I578efe5c2c504f12c8f2466a7f734215 +  ~Ie22b94121b58f17af14c75bfb27f96dd +1;
assign I3350d782125dfaa1c32d06e6ede68e0f      = I578efe5c2c504f12c8f2466a7f734215 +  ~I0d9f8c99194d9d6e187b4ad02fcce8b4 +1;
assign Ia07581cdc470c8ba833acbc8a58f7d0e      = I578efe5c2c504f12c8f2466a7f734215 +  ~I71e101962e766a4d1484b3235359a4b5 +1;
assign Id91d824405f52636dc30344bf8c088ec      = I578efe5c2c504f12c8f2466a7f734215 +  ~If2539da6722562bbf31786fd0036666a +1;
assign I36beed9320665d5988556ea089ee26f8      = I578efe5c2c504f12c8f2466a7f734215 +  ~I22c8ccd4a9018ad1c129aa058bf579d8 +1;
assign If05d018c797e7d4348fe5bd5423b23cb      = I578efe5c2c504f12c8f2466a7f734215 +  ~I83330fef69470d2f5def8e6d7d9c50d2 +1;
assign Ia78ed58e20602b99c01f2208cec79dfd      = I578efe5c2c504f12c8f2466a7f734215 +  ~I0539d598bbe3d50940329a282c801328 +1;
assign I229890d0e3576523fabea29f8594a853      = I578efe5c2c504f12c8f2466a7f734215 +  ~I202f88fdc946494d55fc8831c2e8a34c +1;
assign I3f0ac12bf9d4014f5418383146bcc1ab      = I578efe5c2c504f12c8f2466a7f734215 +  ~I3ee10f6a7785a236db317515fdd23a2d +1;
assign I38e35040b0a7e5476f308d265b7fbf67      = I578efe5c2c504f12c8f2466a7f734215 +  ~I453fdf4fbb5af5bd28a20d7643da9eb2 +1;
assign I90c35b33579355f50d23995dc25cc2af      = I578efe5c2c504f12c8f2466a7f734215 +  ~Ic4a6c02880a9aead7353332708e3f388 +1;
assign I19a71e86490479795328e31521b6b842      = I578efe5c2c504f12c8f2466a7f734215 +  ~I7fb3b66cb48521f8715f66bf5642cdb2 +1;
assign I5505d84d5ef89111fd375ce986e33c52      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I2fd872df07f50688486c0d602cfc5549 +1;
assign Ie47404148e49f0bfa2775b3573dee999      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Iccefa45795486757515d95e5908b306a +1;
assign Ibae1afc3891aaf6fa2751a693cbf5e1c      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ib1357cb20f471f1670ac2448f964f8eb +1;
assign Icbc45a900f0692fde798caa8c1b9b223      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Iab953a8974a1eb619dc0f074c003b5f9 +1;
assign Ib8aaa1d409ba2d09187c3cf4ad4a1fec      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I6e37582849c2c98fd15ad92d22c222da +1;
assign I6a97c95991e02e0e36ec0a1f7c006626      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~If004de0cac6e5f7701a1fce48c6936d5 +1;
assign I30c34fb37caafa3e5870ae3ee43693c1      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ic1efa395cc1fd2c5a1d1559fb169a5a0 +1;
assign I8f23d2c62e919062678a00aa98eff7ea      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I8e96c69e7d872be23229353808c34953 +1;
assign Iaddc9a87ebf5cfb7bbabe07260c592b1      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ib6aded6c73a8cc3cb964b0ae895b859e +1;
assign I24abea8ce306ff137aabea504932da94      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I939368b76d98b43826c68c7f468a5632 +1;
assign Ibee212f9caef9ff8a725aa08e2e955bf      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I544f6263f16cd5e0b7cf28c511a8f6e3 +1;
assign Ie62effeaea232e1a8a50ac3f744f3f3b      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I484545c4d2c869d79eb17f51e11070a3 +1;
assign I6712564d12398f5407fade724db8792c      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I39289e6385a9bc378a9b8dd440249a7f +1;
assign I5a699ad31ee84bb49eff73572bcaf84a      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ie9cce5746a83479a567bbaeac6dbf497 +1;
assign I63f0b04113e2c8b0cf0474f8aa4fc1cb      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~Ic044d7419cc43736d278c2df33b4a3cc +1;
assign I0dd55598c5774df690bb002eefd62dae      = Ida86d05f907d23ff9fed06927c2ec9d9 +  ~I6714551e8885ef5e4490673fe1b2dad1 +1;
assign I361cee04efb7ccdb28fbf44a7f9c3467      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ie9ab3c88ac62369e3d92d110165a94a8 +1;
assign I26225a10fd6209094b91ed34531ca2b4      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~If38feb4f76f761dce6145731ad235d7f +1;
assign Ib269184699c52eafef7d54ca1fda31d7      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I6359856a1843d8c8b65dc478bccb3acd +1;
assign I586e24737da989e9591444e6d260cc9c      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~If6f3d91c3c7a43622b9a522492cd83d3 +1;
assign I01fe0c5ce70d18bdced623e1bfeb55c4      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Id023a6298e65da1f4da3831f5136afc2 +1;
assign I31e6b870600dcb417653fd673d0c1a55      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I6b24690f394792edb0d82b3b9e110851 +1;
assign Id79c1fa529c3b719ef4534d1c3abc975      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I5b55c285f7e3e78447fee68532ab9f7f +1;
assign I496765810959107754d8f764be715da4      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I32701d9e4b96853c53f0ab651a6a4ba2 +1;
assign If1b62fde8c7b6aa858dff5eba22d51a8      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I82f266e5792cdb6e7ebd264e246161f5 +1;
assign I5a86b5c97d7b531c201169167a720d2b      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ibfacfe5b83819afe7fbd4bffa2d6d4e2 +1;
assign I8e0d580b0f875a9373a3d8fb5523183d      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ib8e68a77ad8b9e7cf415bee17645c3f9 +1;
assign I0a35c9a4f7596b64d8a6e39878fbc83a      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I644ee0055a55f54ab3544bb532e39c61 +1;
assign I9eed09a7c7b86123ee154b783cb7e720      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ic5467e42aa377c6ffd8f70673808774f +1;
assign I45efcc842b324efcbf828c6d68f19e84      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ic57eb4a034247a4c952d8224ea9f2bac +1;
assign I4922b2f4381eb54d365a270b32c944c0      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~Ia642db613c0ec1ca4e69afde7a14a839 +1;
assign Ica29fa9ccbb761ae142e6ae7186aa830      = I9d9f8c7a23d9750ec44e706bf763df76 +  ~I432aa7cb844286c442356954f8814260 +1;
assign Ie1e5ff68116424c122e4763955e243ac      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~If520c1cd27f9d4bc52d0d029f693b660 +1;
assign I1c817dbc1d0d04ab8d417d31ef477daf      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~Ie87075ac979410cc11099a356966b8a2 +1;
assign Id4bf2c50adae02e36a8c7a862a470efb      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I6fab46b1766878b26b53f352fee98223 +1;
assign I11f3867bc6c57b2f58b19c0ffbbc0827      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~Ieaf14683f40374c4531326d228cb43c3 +1;
assign I630f6f37116aab84814e74017b6d3c4c      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I5149125aaaad943d891df6a3c2be93a0 +1;
assign I3b0edd5d01b89026be06cf00b6eca7c0      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I770dff588ee1f52f58bea1921cb23383 +1;
assign Ifad4e44440835f78f56065a3aa29ad3f      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I8f0a90e761111a613d2488285534a500 +1;
assign I93a1ba64d41cef26b742ba06755d77a1      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I765a8825e42180a6c63f7b33703bb483 +1;
assign Ib2531654b83ce43d8f11a08c36cca4f7      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I512cc8f6519aa08aee18225b56d47c9f +1;
assign I984fc2e5cd03bcf452fd7eb62be1b5b6      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~If08370fd0e8af818c6db20f43e74034d +1;
assign Ide09ff97f4d7b3049872064c78fd2b14      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I0ff382edfc8051459657ffa3899f5f73 +1;
assign I99c143788bcb9dfcb14e29b1f9117770      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I9d2864024148337277523ef7fa2e1600 +1;
assign I4c4a40069ce9f6b40b8a1ec7787cade1      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I1c85a2d1df6749a194072eb731506bfe +1;
assign I5a345140c4181b5307ea3c5b79e62b11      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I3e3ce8b4ead150a6eae2e5c701c7b598 +1;
assign Ib9e2a08275b9e2571238c39945aba5d2      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I45bc13ae0e0554a79c62cd9c6aa8f2a5 +1;
assign I203718fd22ec9e6e4ac7a9c1973d6837      = I0b41b002a32b8e9e2fe68e819f228fb7 +  ~I92678f5b52c9c55556ff7f17f0f607b7 +1;
assign I8fa60b209a1ac0d2738e58662612206f      = I0e872d4c07169cac84549178fa144274 +  ~Ib4bdc9069d0c08655f5e87f705943eda +1;
assign I579c31eb0b51668db2b1edb1f10a372f      = I0e872d4c07169cac84549178fa144274 +  ~Idbf9094c94c931f16fba468b9dd59a25 +1;
assign I425545d21b0a9447b41481b5874c6a26      = I0e872d4c07169cac84549178fa144274 +  ~I1c3c4ce44610e04c5eef2fcbc2ea5114 +1;
assign I2d1670c45bd1cc15172a12175f7fb906      = I0e872d4c07169cac84549178fa144274 +  ~Ie84be0ae8311d906eff08f7f5b214943 +1;
assign Ia4c9bac1a64e1a17f7964491d880660e      = I0e872d4c07169cac84549178fa144274 +  ~Ic90b98708faa8c8b75d4bd9a52c292f7 +1;
assign Ibff15c9092ff0ab60ccfd9528d5477bf      = I0e872d4c07169cac84549178fa144274 +  ~I8eba6f14f42701d22859fbea94bd1871 +1;
assign Iac2e396e7f63a651c52c6aa372419808      = I0e872d4c07169cac84549178fa144274 +  ~I6d83efa9f988328f487e9232bf2633a2 +1;
assign Ice856d92219493a98683a6e36f6a81f6      = I0e872d4c07169cac84549178fa144274 +  ~Ic23e01562c8a753fd70c343297be288a +1;
assign I5e784ab32ea84026fa63ce432c6f604f      = I0e872d4c07169cac84549178fa144274 +  ~I5669856f88f5e2c98f64df696db76414 +1;
assign I32251a5b768526c3599f145a3eed1949      = I6f4ef0f404ae046519b8436171d51e09 +  ~Ic3a608b850709286ea0ad2f67425d9ac +1;
assign I6357b0d86d75dc1018fa50248f3e2deb      = I6f4ef0f404ae046519b8436171d51e09 +  ~I5267fa34449e6eebe891017fc32d0749 +1;
assign I8a50948f1b1f5589972c137e91e4eee0      = I6f4ef0f404ae046519b8436171d51e09 +  ~I599d01cfe6e54d8e45d64446c446818d +1;
assign Icce2cc29f7ad95af1a9605954033fce0      = I6f4ef0f404ae046519b8436171d51e09 +  ~I8f94dbafaac589ac9f14b56d4556ff96 +1;
assign I276997085c2cbcdac1c886e74bc2e530      = I6f4ef0f404ae046519b8436171d51e09 +  ~I754563caea429d3d0e22df5d193b84eb +1;
assign I7299d046eb7c80908def7e3ec9665c88      = I6f4ef0f404ae046519b8436171d51e09 +  ~If7f373506cac70f8ba1222db135c27e8 +1;
assign I8f993e6b8e7313dfb4323ebf4ccdb640      = I6f4ef0f404ae046519b8436171d51e09 +  ~I69f563e7b7ad483893ac9c4684349769 +1;
assign I2b75fcd754488677526db195256ddc06      = I6f4ef0f404ae046519b8436171d51e09 +  ~Ia0a02781c674fe5d769206448d475245 +1;
assign Ide04235316ff1098fd97e125d76797c2      = I6f4ef0f404ae046519b8436171d51e09 +  ~I1b7a401bc11741e6f011fb9895b5c797 +1;
assign I39755c95fddbe19ae343164be78b0fff      = I4d04e66ad9103a685fbe088b74517452 +  ~Ieb528d666fdb708279184bb59eac25d9 +1;
assign I37d4177c1ea3ac376d3906e49a4a3224      = I4d04e66ad9103a685fbe088b74517452 +  ~Ic3ff7ce12c836bf0693252b9a7a7cfe8 +1;
assign Ifd04130d9f32af7f7debe20de6b6fa57      = I4d04e66ad9103a685fbe088b74517452 +  ~I19bba6a58ad3ef959b33701f82761984 +1;
assign I7ee40f0225ba9aad10df1dec7a0f25fd      = I4d04e66ad9103a685fbe088b74517452 +  ~I8acc93b34974c1e708b0e1591f7b2d3d +1;
assign Ic780d894a72f9111937594d50a9ce311      = I4d04e66ad9103a685fbe088b74517452 +  ~Ib60d4ac0fcadcdfce5a14fb92f58423f +1;
assign I36feeea802ed7e4122a43a71d976b7d2      = I4d04e66ad9103a685fbe088b74517452 +  ~I039f05d5be891a37e04556f1eae674d2 +1;
assign I698319d790c8eb982fb1b113437d93be      = I4d04e66ad9103a685fbe088b74517452 +  ~Id0f75e19b94541ed5c5c352d13390d2d +1;
assign I69c4cabd4c61dd816fbc44ae02f3d8ab      = I4d04e66ad9103a685fbe088b74517452 +  ~Ife1190f76c2e251704c2960c23330a48 +1;
assign Id504dcc780b333a51585556c4b58c610      = I4d04e66ad9103a685fbe088b74517452 +  ~Id3e0c98bff2636e216b4d3a0ffd51054 +1;
assign I0c8aff3de7ee8ede0d8755cb4aebe427      = I988e525020c1e43d238fad41dab4e6ea +  ~If4d3b31b87c0f723241d35ce7e854eba +1;
assign I1898ec6433c0e994bf697eb3b7ae5eb3      = I988e525020c1e43d238fad41dab4e6ea +  ~I72369dedfe36cb22269033cc305b730c +1;
assign I41b391dce086564a0de53aa3f82b510a      = I988e525020c1e43d238fad41dab4e6ea +  ~Iec71fe7fcebccf1ae0d10a5d187fcc44 +1;
assign I90c35450751e2a9607e95ebe3115c51c      = I988e525020c1e43d238fad41dab4e6ea +  ~Ie11da10808c4ca84f399535df6261307 +1;
assign I02be13e15f91f4957ba7086ee96c1ca7      = I988e525020c1e43d238fad41dab4e6ea +  ~I280fa9d114e227cd649bf0e55e845651 +1;
assign I02cc4624a6245c0c54b079dfe50420d4      = I988e525020c1e43d238fad41dab4e6ea +  ~I94c4e11670b4233fa072517a8f19c901 +1;
assign Ib0942c283a523d31d5d11a51f01fa016      = I988e525020c1e43d238fad41dab4e6ea +  ~I4dca2dd40a7127ce44f83b430a34c738 +1;
assign I93ad63d6294ac100b7027b8190f15387      = I988e525020c1e43d238fad41dab4e6ea +  ~I1a24e98165afa62bd14986911a36fb6e +1;
assign I8b92187b5833150d05b4b09f74441a20      = I988e525020c1e43d238fad41dab4e6ea +  ~Ife1164cad7cda4aa9a08d94dfe86add6 +1;
assign I02846f27754a2fbc493cc1d0848b9090      = I90d92887cb2526a2956d5e8c9fad760c +  ~I8d8d95ff26f33f69a182b32ccde23905 +1;
assign Iea2573c99c098c5fe2ee97a9c1aae44d      = I90d92887cb2526a2956d5e8c9fad760c +  ~I2508854bcbab37bd09c9465c377c06aa +1;
assign I8c250d6e46e2d8a7f2f77035526c1f8e      = I90d92887cb2526a2956d5e8c9fad760c +  ~I140078292f7209eccacd53a8bab18016 +1;
assign Ic968e5570985a076b609845c9968110c      = I90d92887cb2526a2956d5e8c9fad760c +  ~I141fb1cbe09f9abe282cffd4de815d25 +1;
assign Iccd14e61a9147bf5aefe4a196485ef03      = I90d92887cb2526a2956d5e8c9fad760c +  ~If79d1d378f7c6fd29fc3335ec5f5c51d +1;
assign I4e09b4d678ce7239bad645b57535df20      = I90d92887cb2526a2956d5e8c9fad760c +  ~I4a41999cea9357a85c73a0af509eeac9 +1;
assign I6bdb1743d21a19cf2ce13b056271d1b0      = I90d92887cb2526a2956d5e8c9fad760c +  ~I8e517c401d62dbb10dcc96ab536f6afb +1;
assign I6259bbd85d21c216632a71648eddae35      = I90d92887cb2526a2956d5e8c9fad760c +  ~I8ad3627f171eadcc960a688ac0afcbc0 +1;
assign I8a654b2420f09bd4b14bc5f5faa7d40d      = I90d92887cb2526a2956d5e8c9fad760c +  ~I85c4d3d6c8408c6f38741257ed177ca6 +1;
assign I50d163f8fe5bbb86e3843bea768f049e      = I90d92887cb2526a2956d5e8c9fad760c +  ~Id66c47fd69c175a4393e975a269cf053 +1;
assign Ic3e2b4869f7ac3d189713dcc40a1fb30      = I90d92887cb2526a2956d5e8c9fad760c +  ~I37dca40506d61bdeab1255ed4892ca20 +1;
assign I3d8f79c5f5af5112dc5f7fdfaf0a2434      = I90d92887cb2526a2956d5e8c9fad760c +  ~I340c98b886123c541a1b8d9fc8a6d48c +1;
assign I0544d6bafecefee496a6227c698a4d1a      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I2dc64c3b06588542b027f997437bee63 +1;
assign I6672e8613ad03882a4b7f4141a56d535      = I00fe3792cde1eeab36e576fd6634c4fa +  ~Id92a37c091100e9df08e24498ecb4022 +1;
assign I1542f0db2447a8b733077daebe1d2321      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I74a4b9365391fd20c34588002ad40547 +1;
assign I3038115e5ee2b90df4a7ad7e25d5337d      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I461195b7ae78743e09ee50486ad6ebe5 +1;
assign I758ce2910b56968ca8ebc74c19f2cb47      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I356d747600182675699a2d2634d4c5ce +1;
assign Ifd3191045c45b2f46fbbb63b1766e9fb      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I87d6a5d30c3e4202cf51f33c7a770c51 +1;
assign I5a15f4c8b810f7234d421967f4d926c6      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I960768a84aec9d5b8bc7c1c523024a25 +1;
assign I6f82614fc25bf322e359b929caa86025      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I09b5273bb15d48a7fd78559930fa6d1c +1;
assign I4dcffaa8c903a955a4c4b5197cd2d728      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I5814a85c45fd0f7be21ed325235fe4b7 +1;
assign I71dbc37567c4c703f28c39b97c44d1dc      = I00fe3792cde1eeab36e576fd6634c4fa +  ~Ib06b60cf9933dd8952206c5f3ccced8e +1;
assign I224678d6b3b2a1ed8f2368d7035134d4      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I67347c413b5efd8ff9e0d5bc7ab2a047 +1;
assign I6942bdfb9c73af7b24e91f3cc2c40443      = I00fe3792cde1eeab36e576fd6634c4fa +  ~I72b1bb104bf2843f161448baf7aab44b +1;
assign I8eae50dae3f5eadae891e7875180bd47      = I6e586c5ac59a28b30c377e51287bf04d +  ~Ib23d889edb5a6d9f27de977d3b1a2616 +1;
assign I5ab8c899cb9e33273d3e5758757dbdfd      = I6e586c5ac59a28b30c377e51287bf04d +  ~Ifaff9dd032cf96487be819c59b03000a +1;
assign I23890d77a1b1c3fea977146599cee178      = I6e586c5ac59a28b30c377e51287bf04d +  ~I028ce03be0618b816e0ecdf43d4cd6e6 +1;
assign Ib311a6a7fc40711d6920e3c43b31c5c2      = I6e586c5ac59a28b30c377e51287bf04d +  ~I6ae2523095237282533e0b5f1c26b488 +1;
assign Ifc3cc051690f3d687caa05e26dde6d93      = I6e586c5ac59a28b30c377e51287bf04d +  ~I5aba6218461e8d571be03a3ef041ebaa +1;
assign Ida60773a931859ee7e5e2db24b9bb72c      = I6e586c5ac59a28b30c377e51287bf04d +  ~I6ca8a1fa2c72b1c61d11dc7d1ba5f37b +1;
assign Id5e39679bbe2407407a53366e77aed13      = I6e586c5ac59a28b30c377e51287bf04d +  ~I3ec5819176ad4b0895a9118d90ab22b5 +1;
assign Ie3eab29a9004627e296a198708459545      = I6e586c5ac59a28b30c377e51287bf04d +  ~I49b64469d298012dbb131d879bff38d6 +1;
assign I86c0872f8ce743bb3fa7b3fca2dea33b      = I6e586c5ac59a28b30c377e51287bf04d +  ~I95361d5f524ccb9feb42811af5c482e2 +1;
assign Id1aa022173e0fa45a3f26b4d31e113a3      = I6e586c5ac59a28b30c377e51287bf04d +  ~I9c4b34b5fb1d59c132bcaeb6258675df +1;
assign I0bfd4314a81f9f0930e549a09ef4c68f      = I6e586c5ac59a28b30c377e51287bf04d +  ~I613d4b1e3b9e812b785c9cf14fefdfe6 +1;
assign I2e90a66f2eedee35927bcb8c5ff26fbe      = I6e586c5ac59a28b30c377e51287bf04d +  ~I848ed394bd4f0b199d11c0ff458394a7 +1;
assign I9d6828434155b5672b44a1172ae9b6eb      = Ib5dc74106d8841d25a793010fdac599a +  ~Ie65a0634454381e24bb3223a333e3ad0 +1;
assign I0483abcf888b35d85e8a62c901b6021b      = Ib5dc74106d8841d25a793010fdac599a +  ~Iad166146f7df5e8068fc6efe4d3e4141 +1;
assign I8f6514c2e33675cd94350a1e1b0b5f80      = Ib5dc74106d8841d25a793010fdac599a +  ~I63e45abd4d27219bddcef06108b72021 +1;
assign I23d3830f616b3be90cd63e45b606fc2e      = Ib5dc74106d8841d25a793010fdac599a +  ~Id1bacd13718f7c29c26b63c239d04dd8 +1;
assign I106ef13f4b977bc5b978b5977cc06eb7      = Ib5dc74106d8841d25a793010fdac599a +  ~Ia3104c69fb4f7abfb5efa3874169a7ad +1;
assign I3fdcbddec1b193cc85d20d4796aef72b      = Ib5dc74106d8841d25a793010fdac599a +  ~Ie1b7257c99831ec5864f65958ecf14fb +1;
assign I3956ec3a4f9d8ea94a760b5c6388f2b0      = Ib5dc74106d8841d25a793010fdac599a +  ~I4accbad1b451ed2b622e15ef9ae16d13 +1;
assign I5541cea9c0da962da2b7d9154c66de98      = Ib5dc74106d8841d25a793010fdac599a +  ~I5ce8b2f633011e89356243a1a71edeb6 +1;
assign I0c1edbaa3c2f47d66034fccd799b5387      = Ib5dc74106d8841d25a793010fdac599a +  ~I3e5139f24e3d082eb31b0e61ea9fa1aa +1;
assign Ia6eb0c9c2e6c3a440defef2c3879de88      = Ib5dc74106d8841d25a793010fdac599a +  ~I61cc8a0f49e393721a62a776e4793deb +1;
assign Ifcef7363a6ecbb3b3248cb65bb6b0d17      = Ib5dc74106d8841d25a793010fdac599a +  ~Ie631e40caade823a196370fc3358f042 +1;
assign I5e36ed7643bf47aef14bd47a835e1a01      = Ib5dc74106d8841d25a793010fdac599a +  ~I4c971e714427664c59c6371e14781bae +1;
assign Idc662c9332f4a6cafe820ad2bc0d16e1      = I3eaf142d2734d2d0decef084dc037b50 +  ~I36ca732e811d67cd742d24fd4cae887b +1;
assign Id51e465dc2adba5eedf6ad37d0a25aa3      = I2d171ad83e27a3745d204849a6f46954 +  ~I354fdd241d5d07f0d8380fe8924e0a8c +1;
assign If0d4550f2f3884c49d1cf5a40251cd58      = I977f1083f5e4f6f8ac38e2c5aecf1b79 +  ~Id38b705f5d2863a020a475ffffc8afd6 +1;
assign I3af1a3cc1733db0dc42ab6214351aa99      = I9bcd673a4293e14fd20b48fa20492df7 +  ~Id6e5d67e7bb7c4b999459374ea80459a +1;
assign I022b7b4693a7e7b654b8bd85a94f0d9c      = Icb7422ea46b22b9330c123b40fe343fe +  ~I05341013abd4206eb66fcddfd63bfe26 +1;
assign I5bd1d6563b4acb8dc10d348ec0a2346a      = Ic414cdba230d7ea73972b0eda1ec6b1b +  ~I15da71a21f5842cb65b543d9bc3e267b +1;
assign I17bbbddc2ace71bcd660f93fdf5e32a4      = Ie4e1e00503dba189b0f871c3c0810d76 +  ~Iccf255fb3422c558465e45226068a16d +1;
assign I4eb0952c6dd9719774c57b76d3cbe87a      = I721c43ab62b42a18c3f5228fc0a73262 +  ~I1c2674b2e6b269ed539827412c5199a5 +1;
assign I6fb63afabfeb4cc43c164e04d35a6c76      = I1f7cb03cf806b247be1cace4d75de942 +  ~I6a3f405bb4a0c4448d9b9d3dd95d036c +1;
assign I91ba6681ef5a1092784cd98b48dc420e      = I775cc766b069022bc00220050feee4e4 +  ~Ib528bb7a64cce4f694081d151fa6fa86 +1;
assign I6eda15abfd6c1f377d25d70e35373596      = I08b78f774ed494fa7f119977bd92679e +  ~Iaa40bd3abf668a21e0f87c7bda7b3f69 +1;
assign Idf9a54c3bd991a031e09982424a8054b      = Ic7dc7f94af108ca7c8003a2d07e1e168 +  ~I919d36a7f6ad42c4bbc23222beb73106 +1;
assign I5d7b50b4839c16d1c7010ef2c8c535c2      = Ibe1327961152cc2d26b3f19476a6e2c9 +  ~I648d2a279dd1f587b1e45eeb35f2fa90 +1;
assign I821836ca9d1bcb5e0d12c348bb323c9a      = I5ba97de444af4e8c9744c3b707502edc +  ~I194a64bef92ecf6714141eaa5d41c9d4 +1;
assign I31f94bb809811efebb378517c2138b7f      = I3e4f1314042010b5d7384693b580da7b +  ~Id332e7f482524adeac7f7cdafcf5ca46 +1;
assign I3f203b62c645fd01c54ed43399b390e5      = I4a47ce6e21c1a274578397e480c184c9 +  ~I226383d68f89db716cfd8d08b837865a +1;
assign Ic01c569fbe524a2fe3626e4d22414e62      = Id184731beb200ad6a53ce273b963bb3e +  ~I2bdf5d319ba9089a4da34b108f5c5ae5 +1;
assign I5a30e151cf8a2259d8cde3fa76389e78      = I3317f2f6eef9a8ef1fe1ff68b47c5d03 +  ~Ia91800792941ec7cc60415c3f844e4ed +1;
assign Ic5340f7fa98175b85f475a03156a04a6      = Ia6b9fa10c79e6f3847f89b35afb4cc59 +  ~Id7c507d96098ee7a955af8a48ee5d72a +1;
assign I0b25b22531e117125c9dc82b1fb69166      = I91e98b804ef82eea53c5e8eccfec827f +  ~Ie15e4c1bcdb0e18085d4b320ac6a925c +1;
assign Ic0c22023bce6b4e011b52acb0ac89944      = I5f1e0d0c6b50f70a6f5584124e095501 +  ~I5485d9edcafc6202f6e5f0969979802f +1;
assign I7f474f465227aa0e2aaa3986574ed756      = Id61fcc605b4b581f5d42024c2610c8b7 +  ~I7fe364f9f537cbef782e7007848a1c10 +1;
assign I8869bb7415e726932972a16630d4090a      = Id64738b7668931553151dbadd5605b71 +  ~I52dcf5bace9cadcf8a895aaa6a8c1da8 +1;
assign Ic1afbad56abd1a486de1d72dc835ea03      = I3bdfb451eb96d256da542864d39024df +  ~I13a9eec6175e695ab8bc4516cf57d6ec +1;
assign I0cc174ebcf049214088dd4a7dad9ebf0      = Ia740d8ccd8230b28d078b2ea3e58d6ba +  ~Iee73a7c685a4cee03f33d3ef379b1c8a +1;
assign If9a4389e51bb56f222cf06e66dcefbbb      = I574050722f82569d34bc2cfae1eedaa9 +  ~I740dc91716e3906ad078e2c7cc3c925a +1;
assign Iff6098f0561da4ad6ee64dbcbf7a8b94      = Ic8f7ec6ee09fb9ee2467e3cea30a44a3 +  ~I514d2dc697e9b39ba027c418a6df6cb9 +1;
assign I26a679e345a21470331cd4fb2512dea0      = I2b77d922a74fdcef0d57debc789bd539 +  ~I782726e317a2aada9e755bcbc4b0d3fa +1;
assign Iec11498f4ab0492570a3454760ed5679      = Ia1d8127af4944b23475bd7deac91d60e +  ~I11eb26cf0f0b3a334e8f7317bf8d9eb0 +1;
assign I78154c0ca0236b79bb58bc2942b0f51b      = I247abcede9914633c0a33fc402bf58ae +  ~I26cb63ba20245b2c332b09e25c4409aa +1;
assign I3a2c3112d5ba223b037baab170e9da79      = I1f413d3e081c6aea012b122fc94f73d5 +  ~Idd7691d31f8d0c09ee988116d574ec59 +1;
assign Ia56b6d58ede63ec2b56533f0804b16df      = I1b812fb764d3b48511c0d15a7efaea29 +  ~Iecc02842a2d2b9b9e8187f2d39e62e05 +1;
assign If8bafc8e64df4d25c725f8c577e6db43      = I88882bd8a9f8718411564221ad85b223 +  ~I5551342f1751fc64f32744a46b9649be +1;
assign Ie7452b79bbda04bebf83147d7f2ddcec      = I232f24e2798488ee66003f3b8cc294c0 +  ~Iff7c29299f005c1cd5a16b64601e727e +1;
assign I29a84f35944a4e286c267c60d9899c62      = I856284e951773518eb6c4232ea7f3d40 +  ~I17a5446e942bcc1dc2c96930e0a87a70 +1;
assign Iae0a8cc0afb8366a7c9df146c0d08eb0      = I82cbeaf5b3e4796b2aaf33dcbd119f4f +  ~I719b67f84e07e90dfd29a8cd5d94cf39 +1;
assign I39d0497d0550115c6a2c08676c451845      = Iaa7791bbc193412e5fe25000ceec23d6 +  ~I2c835dfb3596b8bf057a7cc21122c81f +1;
assign Ia96a79462a86a7ed9e337df66d99bf92      = I44bdc0baed3d51ef54ce2728618ad339 +  ~Ib71b3d357c98dcdfae5c777ca3082275 +1;
assign I8ef19b31ec6d7e52e78b0c673f23ce12      = Ib6bc7e75ce750a26113cbb8895c2f024 +  ~I086bf19f620c8a8f6888e775cb1ed7f4 +1;
assign I8081b1486e6def0f6ae514513c7ef4de      = Ib4188380f7e96d5afb99f5045674193d +  ~I802c554d5b04af6b949677819a4966ed +1;
assign Iee5a68c2d52ef1cdd3f19b0a912603cf      = I5bba219c5024301e420e9a5acbdc5845 +  ~Iceefb06cb3715e1b41e6f7d89420e5ba +1;
assign I4b5525780a9259b57497235bd0bc69a4      = I1bb52988c9ba03e16b1b69335d3d7e7c +  ~I56948bc48c0220893d68004615a6ebaa +1;
assign Ibd65f08dbbf43d438c3a985c7b17f2e3      = I1b9990aaeae716f66b0f89fb02be0a74 +  ~Iec1368f034655d61354ab5b5e94d7d89 +1;
assign Ifaa5785a3e04cd1e3be505042347fe26      = Iceec2cf6aba9138648a3340390f39fe9 +  ~I1e43c0aeeb8a2461d208eba24967af30 +1;
assign If0cb8cd465ff1f65de99688abd92aef2      = Iad7842f3d4672f42c1064c28d4c8ec4e +  ~Ia6eb85b127cf9c1a437611556296b967 +1;
assign I10ff180c115b9372f9b4b12df313372f      = Ie5a53cf9343fdcdb5788667c45fadc83 +  ~Ieba89aa901e61218074af53a2484a74b +1;
assign I64f177202fe847d13a8a12bd80a45946      = I30e06d190906bc9eb6f1c3156c47f9f1 +  ~I8b3b875c6c07bd97ba598a5139156fa4 +1;
assign I5df97e26d5887da447669b8d932fbdd9      = Ieaaaced47e22029ad2945eac9cc45e6c +  ~I7b33ddad346077928620344542b9481e +1;
assign Ibdc07eb6a0a66e1393cb2dbd9ac77c72      = I08dc6f8e837b1f6b80bd3fc742290dab +  ~I11d967a5c5d14c88b5587d4cfed1d05f +1;
assign I3d353247a021629a4dd38a784eba5c1e      = I8eb6a9c907c5909dad6cda98022d70b8 +  ~I27458d76b3ac6520fb379405c6b2956f +1;
assign I20d77ee5328ef46daa4a54c0ae98d31a      = Ia5067b1b458af82c3c2cd50653099854 +  ~I2525111a2fb5f10d64bbd16e148653b8 +1;
assign I8284c3a4664f99934170474b8e0e73bd      = I198c6753cf12d423c709d1512e66fa9b +  ~I7b7cbcd1c6d2a2eeaaff474536a69eed +1;
assign Iaeb44f2b4b78055f103df8070110b5b3      = Ib600dd8a39fda48d28e1289d44d49a84 +  ~Id2a7f0781d18dccc7c4e0b383b7cddfa +1;
assign Ic8242c1f7d2f582c63c3cea63d929945      = Iabf09191227584c76d7fbc634b706d12 +  ~If8bc141d98ebe1be7fa81cde5c65868e +1;
assign Ib9dfa491b9914f9ac567ae8681a2cd6c      = I4869ba08cab90a6dcbc454b0001a7a20 +  ~I8645e1326c66f5efef4b9c923599d1a3 +1;
assign I029b75f94f58485022bf37590df82900      = If97974406672507f8c9a1c507c4b6951 +  ~I0426ef66185128dd1ef4dbb68dcda585 +1;
assign I1cc49a7f6f5c1ecd775d2734c3321364      = I4210341f99ac7cb08245137999739114 +  ~Iddd954df5bae9b4240e0512f746669a9 +1;
assign I596867e7be52dbcabd95cdd2600396a0      = Ic24f4dbd99c8f4d88c8450d4fef762b8 +  ~I29e940970d87e8e09b26ab1b0b8f2286 +1;
assign Iec0928bbbc2730b835fb20d75a988a7a      = I68dffa1a13eb6ab54615347729c1d6af +  ~I488f6d9676aa85a55d030bf12e8997a7 +1;
assign Iabaf04fabdf2dc5fe29d1eae22b23f7e      = I10153d5548b184b9ac2cecdba4ec4b1a +  ~I99d761b75ade1fb2e8afbb1a77752609 +1;
assign I678858a018330bbc4ddb8fe46ff09f49      = I104b7f0512440cffc0fcce25e477f537 +  ~Iac4e3d20178049f9c59abf374752dccc +1;
assign I453a3e7067a9421392ad43b673f203e1      = I18b6758319272eebbe76e1eee5ae55b2 +  ~I618d33f26badabfa578908903a613bce +1;
assign I1a3dcf633defa34860b0db5fed0d710d      = I780263b10b98f9bb0eaf66c045d8d37c +  ~I822d7973afe090b2764335f1b72dfd0e +1;
assign Id4ba510039040276d71a221b3468977e      = I37b772442e55cbcd44ba892a0608d662 +  ~I12c1035353e553b3b6a13bb174ce6020 +1;
assign I7b9204a45b89e3800944d49a811a930f      = I0ac256a6659ff5c6673fd110a8bf578f +  ~Ia6d61947d36fc128c689808c82db80f6 +1;
assign Ia9d671775a9c5d0c1c0886abc70c5100      = If134e1d27e736005e5a390e7a2ea1f4b +  ~Ie9b042f686381739b9ff219041f1e0ce +1;
assign Ief6f4ea0ada586ed46ce19d0761edf66      = I7b37b8f908cd82683832536e02faab0d +  ~I0c4268c01aed70ce4fc71531bf4bb862 +1;
assign I02e35fcbb30d8951f129525146af7f9d      = I08b4bf60c9c7e7229bd1952cc88bc7b3 +  ~Ia34e42f8de91fa4861b0c6cac5dcfc29 +1;
assign Ia55f4e6ae1e56d5aee09414ba7617fc5      = I267d637eb63fef9f4723f7978fad88f0 +  ~Ib7c5850b4f7cc77be2048d114a2128d9 +1;
assign I4f077fadda92556acba301e0990a8d47      = I4fb56a70e5ffa71f58f715da36368e04 +  ~I32bb50faa2b246b2d3b462a79be597c5 +1;
assign I8fc930fd14a7605288eea0d3f7561930      = I5e9e2acb258baf96ac4b525bba54a462 +  ~Idc6d40a49f05c5422758cee50f787eb1 +1;
assign I29eceabd1f5dfb4cc3028ec248645616      = Ic40f61443a4d8f87769067fc39381cb3 +  ~Ide1d7dc22a4b271ef764df14ac22366a +1;
assign If55674824a5a3574ffb2f7da75e2f2d3      = Ieb36710c9a3726f33407436d62639c8d +  ~I7ace6778ac86b3e05939a3fcc716136f +1;
assign I12b13bd78932e54099144478a82ae60d      = Ic804af393da2e4b9c8ef25d4a3b4e8d5 +  ~I044e01e8d2df46e03f00a0af2beb0bf5 +1;
assign I09a98ded5754d5439ec3a384635d63c8      = I52e4c446693c29a42bb3b665f72d382d +  ~I45a7ddcda2662e36b7617dfe64514346 +1;
assign I802fd7e7eb9c1b2fd917b1eb657e71b9      = Idbf02cf10add496d30fa44bbb18458c6 +  ~Idada779a1ac7b844867571d77054b657 +1;
assign I264cc4045cfc24b211d08488ad2eb105      = Ida095585ad26e215f1c1bf989912da89 +  ~Ieeba01b18a244ab8c0ac263c138fabcc +1;
assign Iaa96c298cadeb650acccbd3e548cf281      = I19f1ffa05c7c9a0df5e7014044024c7b +  ~Ie4c9797a955778694dd8615219cb51e7 +1;
assign I463f424b1cc557868a77721849b635a3      = I4d68a2fe778fa93faac38b138138291f +  ~I28a5ed4c239e64c76bb6e566b50cfd23 +1;
assign I5fe371b91ca52980957e017a6dbd2308      = I54393ada6f76ac82c31f2668e228e29d +  ~I79a705ee1e414fe4a5fb14e9b3ce9597 +1;
assign Ia301618cac1f678b17595d3e87a85068      = If5b9ef84f09680f3593250b13a852c1c +  ~I04f90a907f10a7fa1ae3591b48094d5c +1;
assign I0ce7b89ce37757be43c464793608e6da      = Ibb759bc4179e5b7aa759d850c7cfa467 +  ~I31d25b1b49e65216e90b39aa27acd6be +1;
assign I8abcaf2ec878673e81c94be11046e97e      = I05e8b5f8b83f07b609b5ebf272bb2229 +  ~I1f6540c5f037d861dee2c0091cba01ec +1;
assign Ie394af0713a3eb30d9d5c0cb38414b90      = If6ac15373ec1146d38e7aeb71c3ece64 +  ~I9632bb500b7faaaaeb649d74c21cbe8c +1;
assign Idc8ef4846c1f33c0510b0d4c1b027c81      = I2ab3675e1eede757af80716ba980a4e6 +  ~Idd0217a35c3adc8abc7bb581a5df7a2d +1;
assign Ib0e1198c7bb8c8bd611fd9afed1bf0ac      = I388c271687ab31b57421ad57192273ed +  ~Ic05b46168884322644db4e331d37d759 +1;
assign Ib2224de3f3f6f644c9e2278ca159eb90      = I6121679cec8caa51dc5ff0d1a61f9821 +  ~I53c88dc237bb2cd02d50fd7f0a168a48 +1;
assign Iad987f88aaf1b32bee71e96904d0c51f      = Ia0649b990bf5716cfab230127cd5d47f +  ~I7450d4ab3ef0227e93a02bfd620d047b +1;
assign I0831e757dd5e5868bb023dd9004fb68a      = I867a0626ca22108b16267d95c0aadf4f +  ~I2b16e5b4e279bb29c3c675b72083e5fe +1;
assign I64b4330df88134dffb32e0dfd8d4ab36      = I1af54bcb73d7c6b93e55450871207976 +  ~I70c92e8ada46476d15ef4b3c620d2601 +1;
assign I5066c1fb5193c037de084c7463947151      = I91883553543d0425e9c6dd726dce3d27 +  ~Ib193b07804d6d5f111b06bda487bfa5f +1;
assign I76c57762b38b9546bc862bccfde73a81      = Ie95405659701278e3f87bf1f823a037b +  ~I885433b0ab16c6d87abe45af13c9e529 +1;
assign I4720972ec687864e66b86780a4a03e47      = Ia42392e2104b50c0908aad82738a5ee7 +  ~I198c055930cb89d0390c336eda8fed4f +1;
assign Ib0da91fdb282ea40f13881671d9736b3      = I68ad63230a51b9b9e3daffb307ea970d +  ~I688a2c72e69b217d2673e8da75146a83 +1;
assign Ifac345df39972bcecf0cf454e30c0cea      = I7a052d63944ccf42e598efe3a95b88f8 +  ~I3b6fde4ed14cd68af1468ae1d4cc1a22 +1;
assign I47ee2c7239716a56029d9d7dd2efeec2      = I2b3c6d69f79c8d51e4d1614c62c44fcc +  ~I5d3df1e7563630311f56143ee6d97a8e +1;
assign I02398b40df5e80a6818d7f7c20896897      = Ifcef0e92f50e3920bf1208af5d64c632 +  ~I90a7ea789d3bf7f9126c786474a56da0 +1;
assign I5943d30c92a0938ea3933ba61819ce91      = I111340a19625901a3c1b95fd0bd1570e +  ~I5029424c9d9fe923eeb858b1e62cd758 +1;
assign Iab0a2d1699d14959918590a17d221dac      = I11aec4fa85c30f6fe1fd9fa72542ef6c +  ~I1e805c70d50c2765b4a03ad2982dc421 +1;
assign If30544b94b0d43b30a8e4a1a6f67e461      = I80cc333c181c16a96b7bd6501c27c2b3 +  ~Iba58175a7fd5c5da650222193caff0b3 +1;
assign I4d6cdcb3b63c51d9dd8b915eb0645255      = Idc6354325a6280ae9890da33c06c33ec +  ~I7401a0501ba69c5559fbf00c77e58dc5 +1;
assign Id147fa768121368db44934717c87f635      = Ibb04cf82acc4ac16599ad3ddb0c2ada2 +  ~Idd9f7ea657ea9cdcb45a7e4b573b9d50 +1;
assign I7f67e05ed60a537f26feebbbe643a67c      = I3ed096dfd8a14f4acb4d53a70cf8aceb +  ~I53f275395dd6be17961a5edc3e8da7f2 +1;
assign I376c401480a2d8e6131123a91e6fa1cc      = I0fa07f95e96326cb0599c0c3f76e2b48 +  ~Icab010d78cd66b02e089c74f04bf4e75 +1;
assign Ic33856f32df0ab980accff5678cceebb      = I87d98fbc97d9a78c2e7d6a6280e7a49a +  ~I376a48b7e0195a5aacc76a0ad8bd14b2 +1;
assign I97e41b86305179e201cce4d69c2ffa21      = Ib7ddc4dca877f7cf5697a02c3d1915ba +  ~I241622b0367dde514f96ece55c8c3964 +1;
assign Iecaf532a526a0f689b65a6dd749d66cf      = I3612ef280891f6017fad205d0484bde7 +  ~If94a1abfb972f63629d07e64dc23863c +1;
assign Ia54ab64aa44544f38180c57e0864e071      = I561547649aeb5b4c3f10d9506db1f3cf +  ~I07b9b1f4fa01b16cc69356057d3b6154 +1;
assign I8ed5770ee3c9a504d934506743f6b427      = I84cc76c0079b86da7b994844c3ccb875 +  ~I2288a6ad3b748b716249f4adc42d52c4 +1;
assign I7541c0e729546e0e13e98f4658b95a1d      = Iec013c508d0c6401d7eb856e7eb60446 +  ~I022df337bcc05ac5648b8ae2e42f3a76 +1;
assign Id861f8b6cc578cfb1d83d065ae78dedb      = Ifd8979aac6b6b24aa560b46b18240e92 +  ~I60d9a7f95fb8623753002ecaf9a4efcc +1;
assign I6fd4a37bc3b6eb96e6b7e814b203ed21      = If12394e78dc913b01890b56650856a44 +  ~I23a74ea5e7174d95e6d16a5e85ac236b +1;
assign Ie31fceaf1518af42616d21bd8247577a      = I94d18aa10695f3f22b23246884b72822 +  ~Ie697d28d757df82b3901564bda43251c +1;
assign I89ecfbed8d99ec79402dd5f3f1e64100      = Ic90b38835dd7e760dd54067b196f8470 +  ~I8572aedc94f7243ce5eacb332c81eae2 +1;
assign Iddde66a99ea9a0caa45b06e168194488      = If3691ea51f6efe9b165a31964854d2fe +  ~I6734123aaf6320da75638b212812732f +1;
assign Ib645c9e05a543ca3e8ce0994e56aac70      = Ic2ce582555add38a14f5006d3c87eb15 +  ~I7f6dc6f0f403c58f9aaaa70c2383a666 +1;
assign I29fedc646a3ba823d0dcbb3ecb9b9ad6      = I58cc950ee2cbe56b7c5a619be3792511 +  ~I66391978843c39b6acbdb4847a01050a +1;
assign Ie89f6128d6d68c146ffcecb551618321      = I0d8e329ec5873db96df1ec309445a096 +  ~I4f756e4125c8af5c412944b273e01cb0 +1;
assign I3388d6fa5159183888944f2951de9361      = I106325488e2ecfdba1cf9e5201e6bc8c +  ~Id2c9f7ac95de07148c54803f69347f56 +1;
assign I3575e2d60ee8b0b71c67d53b496e2775      = Iff73a0085541a511d3912b64686a82c5 +  ~I5061e13a179d27e1ba5f89ce8ee0fd4a +1;
assign I52cf4fceee16d75ea59dbb574ea7c7b0      = Icdab59de68f2870504598c9ea18f1d2c +  ~I0f7c32fc1548fb49b8041f55c157498a +1;
assign I59cfcae849791453127d60b213ff7355      = I75604d727e82c977741f90113719183a +  ~I89ffab735ee30423c82e079ed98216c5 +1;
assign Ic218ffc97e5e89851d44554326aa5bae      = I6f50c4d0d2639857b2dcca300c2d7b04 +  ~I9494921d8487ee0b314f75cf0380fd2f +1;
assign I6886b93a81c52c7f93b506404b6a4252      = I5cd013a2be2e761c10c6a957632517de +  ~If2b3e7d1541cbd8ffc2b4cfc3ad13a57 +1;
assign Id9c9ac52a48ef3207581bd31c0593b22      = Iafeedddd02428bd2610c576e68d4ae25 +  ~Idf3d79da44f2d686f5bd43c3c1427430 +1;
assign Ib3c08e618350ef723607b4ee58bb4dd1      = I912d6325e34180e0f668f0f024e63581 +  ~If8125ad3c9e7f0a2b84106064d320996 +1;
assign I2481f5b76264c857df96942bdaa941ca      = Id1e05294dfd02df499ad0c08bb5c191b +  ~Ic9018b88fa91fb638bbab0613795ae13 +1;
assign I3a5aa34be4c3adccf4aad2772c38e972      = Id3bb9b100ee4302473b49ac14615e9b0 +  ~Iad4ea0196eb32f9a152c9e6fe5059e46 +1;
assign I95b6796cf442383290a32bad614664e8      = Ief32db1cfc443119b6202b0cc7bf70a2 +  ~Ia8ff29ed728e7f2ae4213f00328b495d +1;
assign Ie45ac55c4add6c3390924c54d2e8d65e      = Iad7dbe9909b5eed3261adf92d3813acc +  ~I70717726200ec02929f679ef05496455 +1;
assign I0935498f4dd90c1fed52d2246ebe326b      = Ie7daf0789c35caaadbba06cafabd2b70 +  ~Iaf1e4c7dae6ad89567836877c08f57d2 +1;
assign Iac314ba0cecbd52f3992323dbce81856      = I2bd1f9b75d9ab94af9ddceb7528935e8 +  ~Icd09aa81e9b43528af73e23b2f0f80cb +1;
assign I2f8a71c2c9078e2581087c7662c961f4      = Ic3d9f5c6677758810e4865779ec303e3 +  ~I6ebb2b94f0f80425f8401ae823d92a1d +1;
assign I38c53b94ea9a59a52cdcfe6681491da8      = I00af04882a25e2832d913a67d4d86d7b +  ~I4a2c3204a6a9936d4a215b46c0ffd045 +1;
assign I5c2c6a0ca07e820e699062299b7064e3      = Ic9db631df0a1a9108c10c3e0eca7bf15 +  ~Ib02c0694762c4815448b2c8d3df767c2 +1;
assign Ia962052eea10222a1c16ce5800e1c063      = I749f9ed1fb2dddd40ebc28f638e02935 +  ~I98cee6efbbe565d3a4de16703189782f +1;
assign I33ecd2de3fc7f48821e40313b5dc2093      = Ia45b2a24df24bd5e3c95885c8928686c +  ~Ibf981c01a9d44cbea3c6d8ead92bc2ab +1;
assign Ie4d5fc4a5bf560bf75561f7f6baa761e      = I7427464fde340780aba7f9847b4ad564 +  ~I864c33e8ea204d20a9baef4584f22d4e +1;
assign I57de351c4dcc2f9c6bacdf1f39961723      = I33fd1ae225e2b881b2b41e0358675e22 +  ~I6ad3228e0e2e1f19648d73e83ba5a229 +1;
assign Ibf1a5a90d4a7922c4bd6273c9a3f1701      = I2e21a35d1cf560936fd19b944a208b6b +  ~Ie099210a99a4899c53baf39559592690 +1;
assign I8a9e51ef30c6434e44fe23412d20425a      = I249522a3d42cc75d7a6b9ede1222ee76 +  ~Ieeec71d9df4613555fade2ced7b3baf1 +1;
assign I796d4045b29e6c1100dfed4a78dbb912      = I68b4c43d9f40ae4bfd70d2983594392c +  ~I4931884e3544af182bcda9061091a42d +1;
assign I32551e388a1ee2ecc7d7da3a4646177e      = I63145e0fec15c7e7c0de105f348bfd31 +  ~Ib3fb10da528d450251764a9b9ede0dba +1;
assign I6c266cffd4d2836af16d4d81bbd11250      = I8af625de86c04016c3424d116fddab5b +  ~Icdc9e676957b2223d60c413331fa982f +1;
assign I9feff48bffd8e1f9eee0a587b4b026d5      = I54c9c10527f83b4ee4e1e22f1e4044ed +  ~I381f6051282c062ccf53866830344cd4 +1;
assign I6c540a2cc92ae1fc269a3a395504a08d      = I972559e47c7f83bd9000ca1cfc14d8e0 +  ~Icfc21935c007fbbceb2a67ebe1a68a0b +1;
assign I683c93eb9205a2272d286e4ad0e998fe      = Ib97a7f941eb7ce2a867503a04ff86a67 +  ~I120d597a80158374726e064fb0f099fb +1;
assign Ic92cbaba339661a83c8bbd3f8377c105      = I5979b55f607c71017537f2b48b40cbea +  ~I2520aa556aadf851f58f0b1820498730 +1;
assign I81850f6963cf07be478907b167cf9206      = I6a56760b621f238843b091279c69897f +  ~I6203f49a08107f7185ebadeecf2c16b0 +1;
assign I6d94790ac6714bb8c62a82bb06960fbf      = Icec45bf76c241d37c9a50a5cd092da9d +  ~Ia706fb593b63cebbee0321c154cb859b +1;
assign Ie19542cb6dc9324368b1ea75a5d5c274      = I2f6d3f61f2890e584d3063a09587e99b +  ~Ia4b5f2b07556629673fc6576bc49a5dc +1;
assign I6c96e6686c458cee66b9d93d6d71f350      = I7c396ea2e959d84fd9a6964617cb29c6 +  ~Ic532c6b85b156f821e0742f47239a65c +1;









   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
            Ib0973b6e90e7678addcb064fded7ce0f <=  1'b0;
            I5033323484d90d6bfbe03749019fc6dd <= {MAX_SUM_WDTH_L{1'b0}};
            Iee06707670e19a82d911c1750bcfc811 <=  1'b0;
            If5dad13ac41b3034bdb034bc86c9b348 <= {MAX_SUM_WDTH_L{1'b0}};
            Id8d5df9e869aaeb107a41a6bca3b89bd <=  1'b0;
            Iac428f9f798618e1ef495c626c41892b <= {MAX_SUM_WDTH_L{1'b0}};
            I507f8602a99a1096e4c293ba3c235bbb <=  1'b0;
            I5a6427c8f18b36d2ea18fe60a0831ef1 <= {MAX_SUM_WDTH_L{1'b0}};
            Ibdf2178bd18783c4797c21e642388d16 <=  1'b0;
            Icc29441eac6ca7a138d45743d37505e3 <= {MAX_SUM_WDTH_L{1'b0}};
            I2c690809d9b9e3482fe5a133b5c00afa <=  1'b0;
            I0e7754dcbc04a4850e052ae4a2fbe328 <= {MAX_SUM_WDTH_L{1'b0}};
            I369ffa98995ba0834f8029ecce705c56 <=  1'b0;
            Ia30c019ed8ce395556494a92e7b42a92 <= {MAX_SUM_WDTH_L{1'b0}};
            I9ccef4c47ae7cfab43584de0f2e193d3 <=  1'b0;
            I9799695ea8244992a6694eaf5c8ae64d <= {MAX_SUM_WDTH_L{1'b0}};
            Ief31fe169c1b360d5933558208dbb602 <=  1'b0;
            I4524cd664b4cb41f642c675fa484c84b <= {MAX_SUM_WDTH_L{1'b0}};
            Ib8c0317dafcfb91b3da5eb5afae1f2e2 <=  1'b0;
            I64e959d80af111ed2fcd54a5407d21bf <= {MAX_SUM_WDTH_L{1'b0}};
            I54e3f08f6f4cf784da57ac39f246b8fd <=  1'b0;
            I3e0da4bcbab4804b5397fb3aa2c94f51 <= {MAX_SUM_WDTH_L{1'b0}};
            I16c7f1b874b0d05c6d120bbede254416 <=  1'b0;
            I3740b30d31f3c61d93a14a46e3199c4d <= {MAX_SUM_WDTH_L{1'b0}};
            I0c3cb2de514ecab0dd311e86a4dc3cdb <=  1'b0;
            Ibf0a30abfec9031737eada436ac1a0d4 <= {MAX_SUM_WDTH_L{1'b0}};
            Icc5ba4554d7a44bc3b43377efbe3b5f8 <=  1'b0;
            Id36e8953a02400a5ab1f4dfdb0422e6d <= {MAX_SUM_WDTH_L{1'b0}};
            I5e51f49adb6dce65a9f19ff736526c4b <=  1'b0;
            Ica71108a53bfcfd1892b4d03ef68110c <= {MAX_SUM_WDTH_L{1'b0}};
            Id57092394c7cda397f42374df4aa3fec <=  1'b0;
            I7c97629ec6e594f9b2160815ddd133cc <= {MAX_SUM_WDTH_L{1'b0}};
            Idd6a4f8ae94c431f2fa3312b4fd287ba <=  1'b0;
            I4823c8239ace86dc399e906c1b5a0d74 <= {MAX_SUM_WDTH_L{1'b0}};
            I9f1f8590dcf596097bc81001d51684b9 <=  1'b0;
            I10ad572ca72c2ea991487c39f7eabd7b <= {MAX_SUM_WDTH_L{1'b0}};
            Icecd765baa87877675b0f3972d78c02f <=  1'b0;
            Ie9f3fd3a6d16316e55addbe0e336519f <= {MAX_SUM_WDTH_L{1'b0}};
            I401a38ea1d71dcc71d17a4694ceb0988 <=  1'b0;
            I07965bca84276dd56da1af98e64b0adc <= {MAX_SUM_WDTH_L{1'b0}};
            I3db9b61e28a51e974e2d5e323ad53c1e <=  1'b0;
            Ic2ade31b8bcf68c4dcc1a371ff14074b <= {MAX_SUM_WDTH_L{1'b0}};
            I96d0a4387f9b959bc779ac13351182cc <=  1'b0;
            Ic0edcf240048fbfde4e938c3e4c5e281 <= {MAX_SUM_WDTH_L{1'b0}};
            I64082bc75fdbeb69a52a4361ed2d5883 <=  1'b0;
            I8b42e89ff5f780d4ef8cd1cd5c99ef61 <= {MAX_SUM_WDTH_L{1'b0}};
            I62929057b7c214bd38fd532e20ba5623 <=  1'b0;
            I70b1b8521b36920707e95fc9418eb8a9 <= {MAX_SUM_WDTH_L{1'b0}};
            I641179f37fef63e7deec603b3291381c <=  1'b0;
            I4fb1c32a62cbbaeb585c6564a3c938f9 <= {MAX_SUM_WDTH_L{1'b0}};
            Iff04b7ec87148f5bd408b4ec4b0590a5 <=  1'b0;
            Iefc37daeec14e14ef2fe0716f73109dc <= {MAX_SUM_WDTH_L{1'b0}};
            I198bfb18d6f91c8f62777e6f592a88fa <=  1'b0;
            Ibd15f164f6d2ac9e5721a21464bc2c5c <= {MAX_SUM_WDTH_L{1'b0}};
            Ia1562c88b4f56d8935c3a5d6ead0f816 <=  1'b0;
            I951dfff9507bb70214d48e03a0ebb3a7 <= {MAX_SUM_WDTH_L{1'b0}};
            Iaccba3030d9d9f8a56f86d6e34ed6325 <=  1'b0;
            Ie78e30b2a2eda75d0df7d10fd67b5e36 <= {MAX_SUM_WDTH_L{1'b0}};
            I953dfeeacee8c44c08d0a425fa549e49 <=  1'b0;
            Ia0b83a372dd4115dc4d61eb8ff0811b9 <= {MAX_SUM_WDTH_L{1'b0}};
            I214a50bf9f879fe747904f4679fdd1f6 <=  1'b0;
            If5c5bcbbea01aa22f242b913f0d01929 <= {MAX_SUM_WDTH_L{1'b0}};
            Ic88f2c344a8ad254fc7d7034cb594f6d <=  1'b0;
            Iccba58cd3519fb4cc75a61b50da1d562 <= {MAX_SUM_WDTH_L{1'b0}};
            If299d1a4e044acbc70bc3b7bce9f86e9 <=  1'b0;
            Ibc0999e4d0b3cc2650f9348b8c204b14 <= {MAX_SUM_WDTH_L{1'b0}};
            Idb373d2cf788f6a93a0e5df7f9179292 <=  1'b0;
            I2aeff1fb4b839a581acaf26f90f9113c <= {MAX_SUM_WDTH_L{1'b0}};
            Ic73b8c8f76a985330d4ac1fa0cc28e7f <=  1'b0;
            I7d60d53f883f8187700c4e78b4c22f1c <= {MAX_SUM_WDTH_L{1'b0}};
            I134dfb2c57d8cdffd2789e2f442c3247 <=  1'b0;
            Id6fcf4b7af4a37c854a12e2ae80851fa <= {MAX_SUM_WDTH_L{1'b0}};
            I0c735e43be8030078ec10bdb6882e79c <=  1'b0;
            Ifa5e5f7d753964f14f0f16dbe552fd85 <= {MAX_SUM_WDTH_L{1'b0}};
            Ie9951415c1d599570af1787767caa2dc <=  1'b0;
            I900d471b087cf5a436c2ad66a84d8280 <= {MAX_SUM_WDTH_L{1'b0}};
            I2630f187d63ba9b0af52c77093e6b760 <=  1'b0;
            I6d1434907f0292ea2ee47cbc5b52bfb9 <= {MAX_SUM_WDTH_L{1'b0}};
            I83db667ace2f04ef4950e2c186e0e6a4 <=  1'b0;
            I938bef7ba7ae1739d8e6a6a7c117a1b1 <= {MAX_SUM_WDTH_L{1'b0}};
            Ie818c5ea3f3b879fded32e6cb06ca546 <=  1'b0;
            I6384a9416b2d1da01df1b2d7b16c5390 <= {MAX_SUM_WDTH_L{1'b0}};
            I3a67a175863091a52844aae6ad277da0 <=  1'b0;
            I5097a79e7cf7a30d38ba198d1407119c <= {MAX_SUM_WDTH_L{1'b0}};
            Ia3aba80aead67feab12e4800fef82322 <=  1'b0;
            Ib113c26c8dcf49c972c41a938059a787 <= {MAX_SUM_WDTH_L{1'b0}};
            I1181d42b560fca7bb5c924a81a5db1fc <=  1'b0;
            I970c4a25a8bce82a9d2846679029fcab <= {MAX_SUM_WDTH_L{1'b0}};
            Ie4e5f3d7c5d2df30653f5666d14567bf <=  1'b0;
            Ibe2af096ad2db26e54d8b4b3bb05175c <= {MAX_SUM_WDTH_L{1'b0}};
            Ifd9345cf219c58291c0b437aac093d78 <=  1'b0;
            Ie48569c467fba0c1291f71d6080ebedc <= {MAX_SUM_WDTH_L{1'b0}};
            I4f2d7bb48918ce51efe6b3b12f9f8e65 <=  1'b0;
            I90e7ded06617b49cdb8b5301fe9c6a20 <= {MAX_SUM_WDTH_L{1'b0}};
            Ifa612e6208151c616c3a0319182a96f1 <=  1'b0;
            I4920014f5d017f4e840dc3b88526955f <= {MAX_SUM_WDTH_L{1'b0}};
            I9cb28a0cc6358610854c8f8d1dd3c707 <=  1'b0;
            I03b70553f1c501609400574ae7cd73f5 <= {MAX_SUM_WDTH_L{1'b0}};
            I40bcc924f5cf1f7d587aa35267022261 <=  1'b0;
            I63c9bf68b43ed66c51b0f4c0ed92e9ab <= {MAX_SUM_WDTH_L{1'b0}};
            I5238f7273b05b8b9f376314acdc6cc42 <=  1'b0;
            If408dfead07757878cc878131bc7d6a3 <= {MAX_SUM_WDTH_L{1'b0}};
            I7137f56eeb4c4ae08bbc238db4cd3441 <=  1'b0;
            Ia0857d63d309807789b6ff4f6028f1b3 <= {MAX_SUM_WDTH_L{1'b0}};
            I02335be013799e2560a98b6a82a0c528 <=  1'b0;
            I53921b825c5e434b63bee0e1ecb7a517 <= {MAX_SUM_WDTH_L{1'b0}};
            Id327bb65156c8307901dfcb4184bb65f <=  1'b0;
            I5e68f84e123c37f19a03c13892c77e19 <= {MAX_SUM_WDTH_L{1'b0}};
            I56331cb7b310613016958553732cdf40 <=  1'b0;
            Id5270b57c6fb4b18db3bbd0a523e467e <= {MAX_SUM_WDTH_L{1'b0}};
            Ie3b00960f8af88a5aba7a2104dfca9a7 <=  1'b0;
            I3c18a84617eb21472d53e598700d7f4c <= {MAX_SUM_WDTH_L{1'b0}};
            I7d1ef47f35b7a4c3ea2e4383732de398 <=  1'b0;
            Id36663e7a01fff3170833ecfecac1321 <= {MAX_SUM_WDTH_L{1'b0}};
            Ibb013f036fc42687a04bdcbe2d0bbd8a <=  1'b0;
            I8d3be15109c7007a79fecaac0d891626 <= {MAX_SUM_WDTH_L{1'b0}};
            I77eae49d321f1d1e39dd7c75829aaedc <=  1'b0;
            I92169cc57291f20d336a479e392ec271 <= {MAX_SUM_WDTH_L{1'b0}};
            I420a4d69a077dc1996ddb4b715d63e15 <=  1'b0;
            I6178b220b469b40dac39168057023a1c <= {MAX_SUM_WDTH_L{1'b0}};
            I652202a4dc8f102d29334b4811f5628d <=  1'b0;
            I55342938216a0ea0889f96c2f6c05ce5 <= {MAX_SUM_WDTH_L{1'b0}};
            I0e33e0cdf39fc4cc99f6696e9f2784de <=  1'b0;
            Idf28431c76a84a48dd895979d2b11a63 <= {MAX_SUM_WDTH_L{1'b0}};
            Ib9479328689dec62f900946e56ba0eb4 <=  1'b0;
            I1ef61124c8d62e8f6a82a729fb091694 <= {MAX_SUM_WDTH_L{1'b0}};
            I2728682c0f749d1a9e8afeacdf44bfb7 <=  1'b0;
            Ib8bb96f0372323e6a8072ca56fb9396d <= {MAX_SUM_WDTH_L{1'b0}};
            I07da3bb5f943db6271fe1867a358df35 <=  1'b0;
            I432f74dda4f6b1cebdf5ad59c659080b <= {MAX_SUM_WDTH_L{1'b0}};
            I61fc44808c85a75909b9d9fd4035f147 <=  1'b0;
            Idc689442305acd00f0f32416d8fb3773 <= {MAX_SUM_WDTH_L{1'b0}};
            Ic5075ee0ad355c20dd45ed594f2a8c3f <=  1'b0;
            Ida03738adc101c03c2229756bed2469d <= {MAX_SUM_WDTH_L{1'b0}};
            Ic0a651f45a502ead495cf14f97d65bfc <=  1'b0;
            I4d14c75f28f3e516c259ea288996131b <= {MAX_SUM_WDTH_L{1'b0}};
            Ic1c05ea22f708f620f626cc8c5ca309c <=  1'b0;
            I6e6cbbf430d57f347a0d70558af143d8 <= {MAX_SUM_WDTH_L{1'b0}};
            I61a18378aadae4556da501ce997321b4 <=  1'b0;
            Ib7487df45118e44acec6b9d07bbd5969 <= {MAX_SUM_WDTH_L{1'b0}};
            Ib1fc521709a1ce2198fd8df5b41d0177 <=  1'b0;
            I492f382fea500462b3d0866240fb91b2 <= {MAX_SUM_WDTH_L{1'b0}};
            I1bb5511c9cda1a595c45ecde48e9ebc7 <=  1'b0;
            I3fb3ebddaf28efb56092d19a1b4695de <= {MAX_SUM_WDTH_L{1'b0}};
            I4a29c37ed36b6e12f1f8e263c92bdbc1 <=  1'b0;
            I22a26b7f0b1c8c16b00597732ce2ab23 <= {MAX_SUM_WDTH_L{1'b0}};
            I4bf02a07719402890405fb2e7b679ed9 <=  1'b0;
            I2ac08a2d8c917ecb37fbaf5325cb0473 <= {MAX_SUM_WDTH_L{1'b0}};
            I75bd82990cb60b6d7ccd7aa2982da7aa <=  1'b0;
            I50ff8f51e75fb9ce3db983c2a0f57196 <= {MAX_SUM_WDTH_L{1'b0}};
            Ia6d3e38249f8a1208540b68f54c46769 <=  1'b0;
            I444bc340ffb7ef7b72d4d2e761d58872 <= {MAX_SUM_WDTH_L{1'b0}};
            Idf548b72357ab28fd956791e84e5d65c <=  1'b0;
            I039c6cac5830759529595a958b7f65c9 <= {MAX_SUM_WDTH_L{1'b0}};
            I50b6f2e0ef2831535ac8c18cd7ca9379 <=  1'b0;
            I0584de7d919236ab138e288a27d08ff1 <= {MAX_SUM_WDTH_L{1'b0}};
            I4003a2515229ca8eb6fefa2bef289ca6 <=  1'b0;
            I086402c82ec67ae09a9e6360c58904b4 <= {MAX_SUM_WDTH_L{1'b0}};
            I48672f8b83eef8c406694676746469e7 <=  1'b0;
            I1cefdc831c146187c77f861b3e2d1af0 <= {MAX_SUM_WDTH_L{1'b0}};
            Ia14a60c9497c0faf3f1f448ff2abe553 <=  1'b0;
            Ida9c16ae57d17b6faee8a54838860447 <= {MAX_SUM_WDTH_L{1'b0}};
            I0ef3962dd323e8ec64c4a881bd4b3044 <=  1'b0;
            Ia3b9fb112f39dd0ccbf7555659369efb <= {MAX_SUM_WDTH_L{1'b0}};
            Ie9b64c34e31dab63c03b3de4528d53fe <=  1'b0;
            Ib1bfcdc0c972aafc99116ed8c0511445 <= {MAX_SUM_WDTH_L{1'b0}};
            I5941476ded9f6dc25d7394f5d133955b <=  1'b0;
            I7adff505c50450a04f1717cac1adebe7 <= {MAX_SUM_WDTH_L{1'b0}};
            Ib46c78ff661ee6fb69c704d39235ffe1 <=  1'b0;
            I699feb4382974a02b21cb387c13f7f3f <= {MAX_SUM_WDTH_L{1'b0}};
            Iadabc5abc7dfbc1dd747179ad7e37850 <=  1'b0;
            Idc99c3b23e49aca3c98f0685ea34441c <= {MAX_SUM_WDTH_L{1'b0}};
            I97a6b5f0976feceee3a5b5890d4d76a0 <=  1'b0;
            Ib67318fa6954ec8f3247927d34e74f8c <= {MAX_SUM_WDTH_L{1'b0}};
            I7217d4790fec9797a1eb8cab1ebce71b <=  1'b0;
            I8774ce3f11362915c4331d1026e452dd <= {MAX_SUM_WDTH_L{1'b0}};
            I3dd024db4130c105a6817e8a4935de0d <=  1'b0;
            I2392b2d17ffed6073875fbe8e92534cf <= {MAX_SUM_WDTH_L{1'b0}};
            Iae502e5a5ae518fb7b817afff28b7932 <=  1'b0;
            I3a4f0d3e32596ef05477f494768d4266 <= {MAX_SUM_WDTH_L{1'b0}};
            Ib8b2b1d90204af5b100379ecad20fc0f <=  1'b0;
            Icd08ff59cf6be3ba97698dd55703339e <= {MAX_SUM_WDTH_L{1'b0}};
            Idf0e651d0b13e167df3c0cc40d149c29 <=  1'b0;
            I985fb7ed22a8476ea322c9e3c2b3851c <= {MAX_SUM_WDTH_L{1'b0}};
            I89daaca029498d05ca62c095db439eb5 <=  1'b0;
            Ib985709316b1b0a9d3fa3c1eaf6c641f <= {MAX_SUM_WDTH_L{1'b0}};
            I0fe5a34ceda936d0924efdd07fad11e5 <=  1'b0;
            I4be898887dff6e2cebe53f135ece131b <= {MAX_SUM_WDTH_L{1'b0}};
            I7876cbb2b5d8aba3652ec8b218080dff <=  1'b0;
            I004db04f61fb57aba81e15cc015442b3 <= {MAX_SUM_WDTH_L{1'b0}};
            If692ff56ce90d22d7af881599c54df75 <=  1'b0;
            I8f7e3dfb2f728d4cd1e79b82b62b0406 <= {MAX_SUM_WDTH_L{1'b0}};
            I18a7a4fe8931c79df3a69223af46c440 <=  1'b0;
            I991054370345e61638ddaf81785505bd <= {MAX_SUM_WDTH_L{1'b0}};
            I8eec3538b8cc9c046954b6804cc656b0 <=  1'b0;
            Ifa1f503965270d10e7a5c9a15576069b <= {MAX_SUM_WDTH_L{1'b0}};
            I653767e659590c1676edf6c25fc0e253 <=  1'b0;
            I24f773842a4742fb58d09cae45717b2f <= {MAX_SUM_WDTH_L{1'b0}};
            I5ff863be142b92dff89f7916d0d088c1 <=  1'b0;
            I5bac7e0d778a547a0ae764fe259b6f7a <= {MAX_SUM_WDTH_L{1'b0}};
            I49f9fd0e0719be527f2a54814dab83ea <=  1'b0;
            I255577ebee6768871df0224fc1db2db3 <= {MAX_SUM_WDTH_L{1'b0}};
            I945f2476eb599844cbee0cd89038e392 <=  1'b0;
            Ia7fb4af3d3529a32f902a52cf5598474 <= {MAX_SUM_WDTH_L{1'b0}};
            Ied0c5f8a9243cd9d93672ad6cc907d21 <=  1'b0;
            I2c98806141f064c9e92935b23a84ede1 <= {MAX_SUM_WDTH_L{1'b0}};
            I9134c7f579723c7615af60b4344efe76 <=  1'b0;
            I5680847bc8d224fa4ed93b2fc0d841e1 <= {MAX_SUM_WDTH_L{1'b0}};
            Ie92388a9d1e71d73c07ed86e9bf6c887 <=  1'b0;
            I365254279ebb10dd7ba0b3482d5e34cd <= {MAX_SUM_WDTH_L{1'b0}};
            I6804fecdf59233c6cf14409bf2f1e430 <=  1'b0;
            I57bf4ad773cc058ae1bb7b1911dc3174 <= {MAX_SUM_WDTH_L{1'b0}};
            I9e777a342bf53eaba0280737ae404bc1 <=  1'b0;
            I57072dfb29c4a3d2e2b40e46e62f0d95 <= {MAX_SUM_WDTH_L{1'b0}};
            Ied53820aab06b5c3423b1d878c71948f <=  1'b0;
            Id8cafb6f76321bdaba9711133be7be99 <= {MAX_SUM_WDTH_L{1'b0}};
            I24cceded372d782c67b33f3a78b16045 <=  1'b0;
            I6344e71ca2b0fd39d36caedd889c3085 <= {MAX_SUM_WDTH_L{1'b0}};
            I2e78d36bca5bfb016af674c343f9c041 <=  1'b0;
            I0c99a68e0bed90afce18807acf7d55bb <= {MAX_SUM_WDTH_L{1'b0}};
            I17a9a995de58643dbbfb78604f26198b <=  1'b0;
            I1c95650979c86310ae2a949961c9db11 <= {MAX_SUM_WDTH_L{1'b0}};
            Iad642c4c62766e8f8bd5a1e9e73bdc80 <=  1'b0;
            I04eaefa5d133e53494fc270b07be7043 <= {MAX_SUM_WDTH_L{1'b0}};
            I96f92481be1ac6cf985b8ab387d326bf <=  1'b0;
            I4a64fa2412eb8058c2dfd9351d7b297d <= {MAX_SUM_WDTH_L{1'b0}};
            Ie03c09039ccafb427153d2347c1caea8 <=  1'b0;
            Ie8bb2fcb752c6a33254963d1ebb4130d <= {MAX_SUM_WDTH_L{1'b0}};
            Ie7381a8294b4cdf669b9c57cfe4012b5 <=  1'b0;
            Iac05b7e3ae18f948b72c356ccfb8000f <= {MAX_SUM_WDTH_L{1'b0}};
            I61c9e3f8e42f869f4c9c1386325100b3 <=  1'b0;
            I27da3f75cca6c49e55db90306aa68e94 <= {MAX_SUM_WDTH_L{1'b0}};
            I24c5b2de59eb1f43fe1efe687231c4b7 <=  1'b0;
            Idc7fed723190098341225fe01ba65ced <= {MAX_SUM_WDTH_L{1'b0}};
            I43d43acde5f831fc32b7bf5f10b9b3a9 <=  1'b0;
            Ife9065805598960919ee4f14c3cc6fd4 <= {MAX_SUM_WDTH_L{1'b0}};
            Ib06e93161fc8ca3be232f4261b04feb1 <=  1'b0;
            I717c5c2d6a2be61593492ae5f17a112f <= {MAX_SUM_WDTH_L{1'b0}};
            Ia0dd00f83afc805036f2c6a0e38f725e <=  1'b0;
            I4c31fa8e6eb648439cdae1de1afe0d6f <= {MAX_SUM_WDTH_L{1'b0}};
            Ib0a0f924fe3757a1e0aade7017ad9277 <=  1'b0;
            Iead549a9af27f1fced7d9c36e7b5c3f5 <= {MAX_SUM_WDTH_L{1'b0}};
            I1ca949071d734d230cdb8adda46c9d79 <=  1'b0;
            I10422eb79364e7d0e21e1643d9060331 <= {MAX_SUM_WDTH_L{1'b0}};
            I40170922c652fa7fa42abc6f580b5e3d <=  1'b0;
            I914cb87eba8baa40cd515334e59f26b2 <= {MAX_SUM_WDTH_L{1'b0}};
            Ib1ad0b531ac9028971d68f533e7ae566 <=  1'b0;
            I32ed679af4ab759901aee43c9d93eb67 <= {MAX_SUM_WDTH_L{1'b0}};
            I0ab0170c7ceffbb58377b65d2ad92093 <=  1'b0;
            Id376dfa5141402f4d41a8858180ed87e <= {MAX_SUM_WDTH_L{1'b0}};
            I9ac68f228a93bbf4aa4a559b1364e42e <=  1'b0;
            I98a384bc62ee03f5ad7df20ef2d9af95 <= {MAX_SUM_WDTH_L{1'b0}};
            I375c5f7eac92d853e85e0606011f3fb0 <=  1'b0;
            Icfed259ca2bb2732d8e0c26ef67cd4cf <= {MAX_SUM_WDTH_L{1'b0}};
            I94f9b1f2e63748c21ec7222c9641366a <=  1'b0;
            I20861535c450d6e6bf11c45dac120454 <= {MAX_SUM_WDTH_L{1'b0}};
            I55500c1d85c4970932be67cc5cd2e023 <=  1'b0;
            I013929385ad819ddfcfcc59c22902ee3 <= {MAX_SUM_WDTH_L{1'b0}};
            I36b487cd1a57a3a503e587fdefbb19e4 <=  1'b0;
            I34fffcb07fe82f11fe142f7c37f39155 <= {MAX_SUM_WDTH_L{1'b0}};
            Icb5350e8c55a2adb370078a7575e28f8 <=  1'b0;
            I61ca60fde05ed88cce714dcd8c13b827 <= {MAX_SUM_WDTH_L{1'b0}};
            I8a7a31327c9e4cbd88ce39fea8971caf <=  1'b0;
            I4907dd45c158dc7e0041c64f1fb388f6 <= {MAX_SUM_WDTH_L{1'b0}};
            Ied069655ed3775819d0bcb722d6d0488 <=  1'b0;
            I2c8f6a9b9f655b317bb0af4d60fdbc4b <= {MAX_SUM_WDTH_L{1'b0}};
            I78a5fc80d42e8db1b56cce5f4c97e325 <=  1'b0;
            Ic7dff631559304ec59f0696c66436d62 <= {MAX_SUM_WDTH_L{1'b0}};
            I3ade7e345432319c1a9c91d4068b3ec9 <=  1'b0;
            I6a239d3e55b4a9a3be9989a85bbec545 <= {MAX_SUM_WDTH_L{1'b0}};
            I88aed46f6dad7a81006562a720670654 <=  1'b0;
            I630f905e55f08e7d1569a08e937ad216 <= {MAX_SUM_WDTH_L{1'b0}};
            I79e574dc9c7e18b695c9a2619b71b995 <=  1'b0;
            I8d13eb3669785c4279c685763d4f3fad <= {MAX_SUM_WDTH_L{1'b0}};
            I800ef583bec1d46d3d4ffdea6b312ef9 <=  1'b0;
            I25a6f3de9a9a01cbbdd32ed848561aa4 <= {MAX_SUM_WDTH_L{1'b0}};
            I56cc5cd6d0a5a4e4601fd48e838fdaf3 <=  1'b0;
            Iba3dd4b2c2c85c4cfe770d9b52ef4634 <= {MAX_SUM_WDTH_L{1'b0}};
            I21047a3955b8b89bdb9013d571b2bd0d <=  1'b0;
            Ie1b744387b5200a504e4874e14d2f282 <= {MAX_SUM_WDTH_L{1'b0}};
            I56eb529a34b484cd20e29958cd6878eb <=  1'b0;
            Icf76cb69aedf4db01cd3444f4c4ba471 <= {MAX_SUM_WDTH_L{1'b0}};
            I74588df6399af2c1112e3fa557e89e17 <=  1'b0;
            I4857b5b50556c8e7fff4b2d3e08e4b28 <= {MAX_SUM_WDTH_L{1'b0}};
            Ic8eae1a92f46db040eb22d726c3a0e6d <=  1'b0;
            I0a1e9cf99f1d4725327615f50fcc3ad0 <= {MAX_SUM_WDTH_L{1'b0}};
            I854a15bc7e9728b01c9a1960f6248dc9 <=  1'b0;
            Ie844f4c446983ce381b0bc4c0e8ef7d7 <= {MAX_SUM_WDTH_L{1'b0}};
            Iae332cfd000fd0529684ab787041b5dc <=  1'b0;
            I6067f47cccceea96ac46ff0d457b25f2 <= {MAX_SUM_WDTH_L{1'b0}};
            I70148fe95244eebf7f0ec953703398de <=  1'b0;
            Ifd6fd1f3cbf8884ca7f64bc42278e4fa <= {MAX_SUM_WDTH_L{1'b0}};
            I24ee2d953e65fefdc73b3d3c4c0ddd05 <=  1'b0;
            Iaec9fd9e79371676bfa8ff14b4feae52 <= {MAX_SUM_WDTH_L{1'b0}};
            Ie3a5f8eec283fd4f682b5d0f909b051c <=  1'b0;
            I500757c4eda5d3d899aee47b87da585b <= {MAX_SUM_WDTH_L{1'b0}};
            I781d986d7fd6c2fec3a8cf3f29545174 <=  1'b0;
            I47bf091b0fa74ad511a760bad9d2506c <= {MAX_SUM_WDTH_L{1'b0}};
            Ib4db8131350f8605e00907234aff901d <=  1'b0;
            Ia4c3d0cd9957f678880de5775de76e0d <= {MAX_SUM_WDTH_L{1'b0}};
            Ie093f0750b60d3aed75705637933f34c <=  1'b0;
            If5f957fa2f055b1c2c28e8d7cfe3e9ad <= {MAX_SUM_WDTH_L{1'b0}};
            Id2fba7c1b3dc7a75a5e0d90494d56962 <=  1'b0;
            I3608378a5da8c66bef58528d56192530 <= {MAX_SUM_WDTH_L{1'b0}};
            I9ecee74c445711a376133636ef414666 <=  1'b0;
            Ie6dead855e00ea0a8e6a9b7503aaebb8 <= {MAX_SUM_WDTH_L{1'b0}};
            Ifb3cf6b88835d27220df837682c4dc93 <=  1'b0;
            I3bae5e6862e003a8b9a476f72cc6858b <= {MAX_SUM_WDTH_L{1'b0}};
            I386fbb3bd550891d682e137044e8773a <=  1'b0;
            I4431adecba8be9e5f21bc6b3e1f8cb10 <= {MAX_SUM_WDTH_L{1'b0}};
            I7ede7d2e1c2730b3b71340b11e880f5b <=  1'b0;
            I21c7a2885126d532d00484376588a469 <= {MAX_SUM_WDTH_L{1'b0}};
            I64c65fad4a7d958d625c783626808175 <=  1'b0;
            I2c4d7339ff2fe68d060dd8d961dcab8c <= {MAX_SUM_WDTH_L{1'b0}};
            Ib2e0cd0a2b51c3a265bdd20834c0ed2d <=  1'b0;
            Iee518b15b067eec58cccfa37f7432ea5 <= {MAX_SUM_WDTH_L{1'b0}};
            I67be0b66c8d0680eb23290a4b3885af3 <=  1'b0;
            I42145be9c2a80288ba4a2edd91f661a3 <= {MAX_SUM_WDTH_L{1'b0}};
            I01148401f7d058614dc1ae6ed3c8bd94 <=  1'b0;
            I9dc297ad41fafcda77f5347f331cfc25 <= {MAX_SUM_WDTH_L{1'b0}};
            I3394319c370daf6102be00d938d55769 <=  1'b0;
            I846700c79f30ca954cc2933fc94d355b <= {MAX_SUM_WDTH_L{1'b0}};
            I24d6a334dd15ccdea558f32cd029e6d1 <=  1'b0;
            I8af96a91457316e49e3f7dd5e57c82da <= {MAX_SUM_WDTH_L{1'b0}};
            I3a41f68bca2d7edd1f5738c4fda8e73c <=  1'b0;
            I7d1c247500d7d32e406b2a5f7e2b745b <= {MAX_SUM_WDTH_L{1'b0}};
            I9ef1784d165492f3482d14f475732451 <=  1'b0;
            I66d85c030a8864505298919046056305 <= {MAX_SUM_WDTH_L{1'b0}};
            I9d9378337a77515a4e8d04fb88938808 <=  1'b0;
            I4841257ae596d9d3e4eb1e6f886956b0 <= {MAX_SUM_WDTH_L{1'b0}};
            If0e20ef9aa69b77ae0e58ca3dfc9998f <=  1'b0;
            Icd6f7ec117f9ab4eda8c5eba41386ffa <= {MAX_SUM_WDTH_L{1'b0}};
            Iec2cb48bb1b58f268bf164d5e8a8120f <=  1'b0;
            Ibc0498839d1d9b6dc853b8e5d7a88fa3 <= {MAX_SUM_WDTH_L{1'b0}};
            Ia4ae7c98720d43a604f28dfc5dd67d50 <=  1'b0;
            I142ebca7f155e287e38ddf45423ab0fd <= {MAX_SUM_WDTH_L{1'b0}};
       end else begin
          Ib0973b6e90e7678addcb064fded7ce0f <=
            I5b177dd5c14ad082516b47f550875682 ^
            I477326720157df2503149125a43ee987 ^
            I319012bc6fe93d78de57bcace0caaef5 ^
            I174b6c36f2af82f8047cc76543a3b4ee ^
            I8fd5787ebf758919e7cb75d7419441e8 ^
            I413b1c1985a6c9c6f202e85ff901e3a8 ^
            Iea3e35ece9fdb3aff3b9ff5369e9a7e0 ^
            I30c0fcd89e0cc7c5fa348df7b4fa2ccf ^
            exp_syn[0];
          Iee06707670e19a82d911c1750bcfc811 <=
            I77b05a8aa92c66a235195a66dc13c0cc ^
            I876fdba97e755b74532f7ab191fbac14 ^
            I5590d801fd7fb496019d4c31b7c6d898 ^
            I25f1ee9cee4d04bd8fec1fe601d016d7 ^
            Ifebcf64858d5e2d07ad7894d6182eb11 ^
            I163cf58b9a308e0439a8dc7c1526e6b5 ^
            I3347717ba9556e69de30ce7533d4f5a4 ^
            I5f96a68d20e3ebc71dad4b43305baa20 ^
            exp_syn[1];
          Id8d5df9e869aaeb107a41a6bca3b89bd <=
            Ie117f6ec475f5d6444998af151ce4e69 ^
            Ia538dadbd6ae3711740595a18c89b65d ^
            I141cda06bae0c5666e3bc61c6fe5ad66 ^
            Ifb70a30f8bade95f402e71f95fe6644b ^
            Ie50aca688b3433fad7565998cb900155 ^
            Ied33f18cbb778d5ba744d249f91c950b ^
            Ibe97860165dc5d9a076ebd935385ae51 ^
            Ie46b71f55aef4d00168202431d47dce0 ^
            exp_syn[2];
          I507f8602a99a1096e4c293ba3c235bbb <=
            I92cb615e2c439914e72ce001256518e4 ^
            I7d6a6026eb3c4d06e682523424f9628f ^
            I06ad520cb02e46d34c45f207d42a9243 ^
            Ifa3df8b249467cc1e827c69925ef415f ^
            I4ba41864bb1d2130c6971e0b2903027a ^
            Ia67f9b902a21de0414eb8dda52171991 ^
            Idbbf2ce4a30787c5f07c3b908a73da75 ^
            I71d3a999d88e591e102398409b3adebf ^
            exp_syn[3];
          Ibdf2178bd18783c4797c21e642388d16 <=
            If7f3174da35dd39af7f4792aaa649bf1 ^
            I953b975a89adcc88039284970e9b3404 ^
            I5a247475beb737d470f03507e55f5b24 ^
            I93084ccf5b5e4efaee968b497bb2a775 ^
            Ibab55499323660588ec82ebd07ab0572 ^
            If9285bf7611bcc5ea6432215c349e021 ^
            I3566033cf5c9a06977c9182925750707 ^
            I87b10521099179c18652c86d5887c908 ^
            I13a98f98c54b2e412cd88c96f016c41b ^
            I6f7a45fe64ffeda9ed120be3a4519aea ^
            exp_syn[4];
          I2c690809d9b9e3482fe5a133b5c00afa <=
            Iad799775eb657f8973e6dfcf70a9875c ^
            I5ec1e530b9007a75a778af4d82ab427b ^
            Idd59a5357d4c835379ed180ac0924bf1 ^
            I7a626ec321bf963a5401892a7e3891c7 ^
            I3342fe0c5d3ee5021892d53eb45bde21 ^
            Ia858ff5551286beffd4cf82f876d30ac ^
            I5402fd208dc7ca81dfd2920a9cfa2715 ^
            Ic32c6734132776c290155a80025fe366 ^
            I5d92fdff96b9cd64f3af2b28b13e9956 ^
            I221524a69e18854f029cad30e8f94e8a ^
            exp_syn[5];
          I369ffa98995ba0834f8029ecce705c56 <=
            I55e4ad2d71a29ad63b4999d64ac0dc4f ^
            I592a495aecc800236c3470ff8e6adbb5 ^
            Ifdb5589982db805a0416e1c01276249a ^
            I0c47ccef4b55410286248884a7249703 ^
            Ib68deeb7bec4ca3585d1a4dcbf8793f1 ^
            Ia17906696bd0e095d7a5297da2e049ea ^
            Ic11a6b77b84c44180eb99220a0c4c9f6 ^
            Ie08ad9bd71329858c1742c8f571a1c36 ^
            I8c0c1a0a35f4f7a688f516c567242d39 ^
            Ib105151d91678f81978495ff94b1e651 ^
            exp_syn[6];
          I9ccef4c47ae7cfab43584de0f2e193d3 <=
            Ie92110d19f4886cdfcfacd0920c06a4e ^
            Icf3ad912aaeaa0c5cd1ab0edb898d6e8 ^
            I857d3155df0b6dd704514b039c66fa97 ^
            I3bc094d67805664859fdcb66f1360e64 ^
            Id14074d5230885c38b89b09b130ecf68 ^
            Ibf312ae4f51fbc44b43848f9df62a45f ^
            If6ce2fa9f0b8bc74442ed8262b5089cf ^
            Ibabf61085ca7af8dfc7927b3656a76f7 ^
            Iebecd2d19f9174d87deedc1a273e7baa ^
            I94a9de743d5bedbea3876de954f479bd ^
            exp_syn[7];
          Ief31fe169c1b360d5933558208dbb602 <=
            I59c5da6338f431a626c86a065a355c35 ^
            I8edf1a08ef943f06ee28771c6e140e28 ^
            I1c8024aa9d81704d2dcf63e34853f8cf ^
            Idc1b8aa2f81a7fbd87e4f5821d14bf01 ^
            I02812a8a833bb69eb168a1004b6fafdf ^
            Ic44eab478be232721e7a43d14beca32f ^
            Id1dafb7e45b860d506e0c2c91b28142e ^
            I9db50007841762c9a10f6b7e9d40f858 ^
            exp_syn[8];
          Ib8c0317dafcfb91b3da5eb5afae1f2e2 <=
            I36ba87b69b5b9dd919319230f697dfad ^
            Ie7d9730b191781c78391141d95d4f8bd ^
            Ib774f380e3d7cfd1f5f064e93d8134b4 ^
            I13b0c9578f7b6b3b7e6704d7b44079c4 ^
            Ia01c82761aeb124cd92fb15ee367ee8b ^
            I2db290170ddae8dc52ce07edaf48b365 ^
            Ied764ee7730ad129b6f62837ef50774a ^
            Idc5dd6caa4ed17a63746d30d381a944e ^
            exp_syn[9];
          I54e3f08f6f4cf784da57ac39f246b8fd <=
            I719a892ad54e63b217c7271741b29cc5 ^
            Ia0c192e590d8c914555b434ce5a634a8 ^
            If2b40d249c531e10cc22d1335f350441 ^
            Ibe7e5c2cb9c50eca34a3859d13e83a92 ^
            If0970d9f7b053fce3ced3521b4885588 ^
            I777ee54ff20d0544af18ad8a870d6915 ^
            I4edd64d1f1da865b1eb886e22726a033 ^
            I4dbabfd592b74aef93b819163130ef5e ^
            exp_syn[10];
          I16c7f1b874b0d05c6d120bbede254416 <=
            Ifb064c69c7110c014593149ae69c75fb ^
            I2c741a5fed7d88e9bdd6b7459feac649 ^
            I8a9e516aa824260998d10db758642bb0 ^
            I8bb5522183b65583fda83067990b3e94 ^
            Ib0001d7298ad1f3b1c7603173a70d8b5 ^
            Ibc9a860879ccc58c815b9f6caa23320a ^
            I17c9d8f658dd6b2916b645d103f4702a ^
            Iba283e99a57d0a3b78ad2e309c316b65 ^
            exp_syn[11];
          I0c3cb2de514ecab0dd311e86a4dc3cdb <=
            Ic98c8641d2022080297c54ff2539e75d ^
            Ia9c273b32d0701c7f185ab2de9e57829 ^
            Ibf5c141c5cc0a6a20c05b52bf8282476 ^
            I2518ccf385b3b677d95983bc550282e8 ^
            I86fefad34d3c864dd0e725133f303b4f ^
            I180d4f3b23b518271d7cb8189fbeadc5 ^
            Ic7ebdc317c978eb275eca41d5b9106a5 ^
            I84057a3b319ab3d6a2ed8f2310f970fc ^
            Ifab075b1437495268b6a3be4cb022e71 ^
            I89c5af1a6176cefa1f77ee69996473cb ^
            exp_syn[12];
          Icc5ba4554d7a44bc3b43377efbe3b5f8 <=
            I17a6511072c7fb4846be5844decf17d6 ^
            I9d18ff3465afd8cae63abba68487542e ^
            I1e77fe6aeaba852aba34ed37dd53add6 ^
            Id38852415486e6989b89a0d85ad6771b ^
            I89af7644c48a80d7d22f50b008d35841 ^
            Icfc03646b36b971b9fa57d04a26dbfc4 ^
            I05e739fc87e962848f265e2c73338cac ^
            I624958486d181501c7a8ec2642cb503c ^
            Idd775d9fe6fa8dbdbfb07d4071b9caa5 ^
            I17086dc5193aa55e5c6f56ecd365cc00 ^
            exp_syn[13];
          I5e51f49adb6dce65a9f19ff736526c4b <=
            I7e12ad8a8ef857e02f4563b2f3a7f0ca ^
            Ibb35bace971548c9fc98d773d1aff712 ^
            I68b585571699a57bc6ba5e8955467119 ^
            If76f04fe0baf171d7df2c0cd849aea2b ^
            I5134b762ac428bed07ce102d8927a418 ^
            Id277f5f05551eeb5dec1701056330da1 ^
            Ie886c5effc85f1fe0b6411db4a2cde77 ^
            I3c10d579f80bd0106506ad047d75f188 ^
            Id18c5a1d4eaa73a94e699e5f9e3c3d35 ^
            I9ece87047aec25abc02a5eea72f0e647 ^
            exp_syn[14];
          Id57092394c7cda397f42374df4aa3fec <=
            I12f2f886517647044cc251861721bbb9 ^
            I27e1d2e0e980216b27b90ea48c061025 ^
            I41eff06fe1dea8be4613945de596d3ca ^
            I94e4041b482064334fd0ed92b91bde89 ^
            Ida3d808d100e0bba290f96ed9e744e65 ^
            I4c66570630a650fa7b9bec543f685487 ^
            Ib1a40247057324b0bd810c844bf11f51 ^
            Iddc5b5b4501f9f13bcaf22081e5a70f4 ^
            Ia71cf07b645c58cffe33be1a9a960eb2 ^
            Ifba3e46933049cb093d2c1809f3a8a3e ^
            exp_syn[15];
          Idd6a4f8ae94c431f2fa3312b4fd287ba <=
            I4acf6d84471cd237f65c9b2391b7a20c ^
            I17b3a9df6752da6cc987e902e6bbad48 ^
            I168afc1863f909dbcb6a9230db9f3e00 ^
            I989dda9add29306d7b3c0f376822763a ^
            exp_syn[16];
          I9f1f8590dcf596097bc81001d51684b9 <=
            I7f7b30f2acbb8e31f50b58096b738254 ^
            I615053b36a1851a06125e2ed5ec7f880 ^
            I9890f7fc708c7b8cf460849b4a30025b ^
            Ibc929201e2eeb3e61cc8f0acbade497a ^
            exp_syn[17];
          Icecd765baa87877675b0f3972d78c02f <=
            Ia098bbeda8b755ece6b88eac83d03e55 ^
            I87f34821cd0b58f8855b25c75f2dd32d ^
            Iab2f643f81921ed8464e1bbd9fa8c68e ^
            Ib0dfbbbca2d3d264065f73b4241caed5 ^
            exp_syn[18];
          I401a38ea1d71dcc71d17a4694ceb0988 <=
            Id20e72ac258d1d1b6cdca1e6c9e3596d ^
            I5ebc3047985651f4b9a957d502a97e95 ^
            I53222c82827cab7c770e057ae91bc10e ^
            I339786aa60d4c71d12c65db27ac420fe ^
            exp_syn[19];
          I3db9b61e28a51e974e2d5e323ad53c1e <=
            I7a387a1f887c32e9d0f8e89912a8618c ^
            Ifa09fc1b009d073d5a9973b430c63469 ^
            Ia9c8cc5e3becf3d48feedec8fa2c93a4 ^
            I4f134c0669b5a6a8c7e03be7eee30c6c ^
            I1c4b29e48d0effac4839037ae5688334 ^
            I3ade020bbdf8f954821f737439513043 ^
            exp_syn[20];
          I96d0a4387f9b959bc779ac13351182cc <=
            Iefe4099ff7e457f6b9fefc83e176c1a0 ^
            I487496233a32f657171b3789590d0522 ^
            I39d3bce4060032a81e6b6a1c1805cfe8 ^
            I9963d0b24763ed8038b1f3922b8f9548 ^
            I5e69e930a318dcb0594a823b3129d650 ^
            Ia50526cd3a3174bebc5a7a0889fda661 ^
            exp_syn[21];
          I64082bc75fdbeb69a52a4361ed2d5883 <=
            Ie7470dd75b54d14038de19e4d3043ba9 ^
            Ifbc6aa14cd448bbe416897a3671ba857 ^
            I7547c56b32513ad45d775b4502596d9d ^
            If10f33385e236eaba56cbab8c2883399 ^
            I17d7f36fdade16dbcf621fe302bd7e57 ^
            Ie9f37dba0791359bc426a73639ce33ad ^
            exp_syn[22];
          I62929057b7c214bd38fd532e20ba5623 <=
            Ifc34f5d6b7a7d0533439794958959856 ^
            I87211ac14d832ad3205d47fb83cf256a ^
            I17cf58ef5326978c62c03c56090a299f ^
            Id79636d195efff260c430978f0bcee9c ^
            I8015717cd36aabbf2cf4aa3a5c234690 ^
            I9518532a8617fc8290eb6a5e981dea94 ^
            exp_syn[23];
          I641179f37fef63e7deec603b3291381c <=
            Ib862ac63c230ccde7fae0e62f9d047fe ^
            I013d84bfd582acc7accf07ec522961fa ^
            I7cb58e4c486e683faa4acad4756815d5 ^
            I67d57e38df8cb35ca686ac2eb44e233e ^
            Ic0c13c9a929c8c46e8702cef74de8955 ^
            If66524125bfde5aa48ac70c4e448b38f ^
            exp_syn[24];
          Iff04b7ec87148f5bd408b4ec4b0590a5 <=
            Icddb43f9b760a4597a0bb637fb405616 ^
            Ie41ca18c7d11a47e274f9c33f75393ec ^
            Idbf4ad11ab2a27044193448c8739fec6 ^
            I04864c28351edb33b61a103add6fb875 ^
            I431fc2e9533012c8571d8158d4777dea ^
            Ic3ec6375998b05a3e48f6c5fe7b3910b ^
            exp_syn[25];
          I198bfb18d6f91c8f62777e6f592a88fa <=
            Ie95662d4faf6b5a4cd5ecfa41697b983 ^
            If3b77c41fabcdb283f2c6fdacaa5e9a4 ^
            I6c765e677f42fe600b848698c8a78349 ^
            Ieca2767ac27170058499d83016447aa7 ^
            I403303228c0df825f67436f4a7e64061 ^
            I0ac421af6e311b6005c3e02e93ff94ce ^
            exp_syn[26];
          Ia1562c88b4f56d8935c3a5d6ead0f816 <=
            I849ee5d34760be03d4285185136aa52e ^
            Ifb422c30663eb4824caa72326b238df6 ^
            Ia98de3691917dfb63bebdc3f8655c8be ^
            I67f87fbb746dd937fffc534c596f36c4 ^
            I23afd747ecece714e32fbb896b5c022a ^
            Ib9db80f43718305a8a8774d8d80c86c9 ^
            exp_syn[27];
          Iaccba3030d9d9f8a56f86d6e34ed6325 <=
            Ie6212a29c7c6b035cfff4c869f945b68 ^
            I41ab6fb6ec6ef7ffff70e50f25f217b6 ^
            I0bce960fcc58938e6a1e01b912eabbf2 ^
            Ief72606c77113ae37845e4aa4a2ae5e7 ^
            I5ede62333e0f7ddc5446b653ba9a2382 ^
            I3b775b06b5d78fcd7373c966a62f44ad ^
            exp_syn[28];
          I953dfeeacee8c44c08d0a425fa549e49 <=
            Ie34534dfd435b3d1cf35e82ca71e83ba ^
            I0ec27b590ee6dcdd9c1086105e3b6c23 ^
            I452e51cca9acec44e36e4efd21b43034 ^
            I946246be5b4745508b7d4b578f83aaa2 ^
            Ib2fe0f68044c11f879e512a200f8099e ^
            If2372a5956f21f97eeb9c76281b6675e ^
            exp_syn[29];
          I214a50bf9f879fe747904f4679fdd1f6 <=
            Ie596289582a73e37f78f4ca4cab21e3c ^
            I7b80b4902fe98c10dd72c9eb082346e5 ^
            I3051f561a5e1131ebf167cb6ccb5adf4 ^
            I388528eaf83566cc56b23485a9c05962 ^
            I3ed6426fbdba8aaf1c948cca7442b3a6 ^
            I7b32c2b108e24750e2a24785668af3ea ^
            exp_syn[30];
          Ic88f2c344a8ad254fc7d7034cb594f6d <=
            Ib81431cfb3b281555fa7e5b4582a2524 ^
            Ie5373b01a92f2ff85be8077cfef2175a ^
            I284b23051c85300c2a1e3afe8f25e99e ^
            I71d7f72d83b7410de31e09ea96adb95c ^
            I4af3e2bf2ebc913ac902b48da672c5b6 ^
            I8ec99197a7d823f5745d382c10161430 ^
            exp_syn[31];
          If299d1a4e044acbc70bc3b7bce9f86e9 <=
            Ia3559d98eb372b7307f30ad1f7c4c7cd ^
            I0e8679271ba733bb87c44b6b9f0b6ed2 ^
            Ia7c9c24f8e993526e76c6915e56908c4 ^
            Ib895fec0b3756932b85962c1d129a03e ^
            exp_syn[32];
          Idb373d2cf788f6a93a0e5df7f9179292 <=
            I8f1a8a22637d37c3692e808d5eb3d543 ^
            Ifad8c7bacf72583f91be27fbe5b7a1e1 ^
            I384e50fa8daa639124f083dda56fac00 ^
            I76aab345d13c6678fe37a4a7133cfd7d ^
            exp_syn[33];
          Ic73b8c8f76a985330d4ac1fa0cc28e7f <=
            Ic76e72b434b47c10ebac3fac4ea50bde ^
            I835b902949c2c4c09b757d4d35574a76 ^
            I5f1609647f1e71cef4ba2d605c6c8445 ^
            Ib4f368fa3d3ec11d9ffb2ae9a2ae6310 ^
            exp_syn[34];
          I134dfb2c57d8cdffd2789e2f442c3247 <=
            Ia1b617e3d141263b51e58c5ef0bd7a89 ^
            If343015b4815b01dae88bbb6f2017b3d ^
            Ic98f33c6a4613534bcc9b6bc4b4f2d17 ^
            Idd0f3cfc5599481c954a2bfe69f044e5 ^
            exp_syn[35];
          I0c735e43be8030078ec10bdb6882e79c <=
            Ie74c72742807ae4243748fd27d80d626 ^
            Ied8bd4b6fd0e4fbcced6d20eb7435f55 ^
            I6cbc06919b9c695d99621db6f8d768cb ^
            I641539560711ff1824bd90baa0f21f96 ^
            Ie624c4dad5036a25ca314b94cf3c4b95 ^
            exp_syn[36];
          Ie9951415c1d599570af1787767caa2dc <=
            I8510240df7dc41f85ad58a39868a1fd7 ^
            Ibe3d3e6bc58efc2e9d9eb1f96cdfe424 ^
            I72939e49bf2d9c6a84e404419fc644a1 ^
            I95f0acd4f955058041c035789c3a4d99 ^
            Ibf4b3caa5655cfb6663f9b7e2383bbbf ^
            exp_syn[37];
          I2630f187d63ba9b0af52c77093e6b760 <=
            Ia0116a3cebf94318ed5b287960957ad6 ^
            Iaaaf373f7e6f55214915b93da9bd71d3 ^
            I0ceb14ac0187d804f9692e0c55b8e941 ^
            Iea424dd9d8916c4951b8746408b8a521 ^
            I049d1c09c15def12ba7bae95fc1c3d55 ^
            exp_syn[38];
          I83db667ace2f04ef4950e2c186e0e6a4 <=
            Ic14760b65c6fe150c3c48e64389a41d8 ^
            Ibab1d13cd6a4f7b0c79c9f845339e53f ^
            I2919272e9ae3996a3e1d602ff72ba86d ^
            I1db4ea6916125702e7fb09d0f742e60a ^
            Ide06ba186ddb179b489ba6e3e209e3e8 ^
            exp_syn[39];
          Ie818c5ea3f3b879fded32e6cb06ca546 <=
            I6f420c64640dfb0c001f57df7e3b4504 ^
            Id75c23e80cdf25d883806ed20d4ae783 ^
            I4d4901ff372f6820ca9c8c29cefa664a ^
            Ice0234f25de4ab1f03a3cb01a2d61dbf ^
            I1b78785ebe2e7f77a3125a6334c4dc54 ^
            exp_syn[40];
          I3a67a175863091a52844aae6ad277da0 <=
            I9eb87e62d23bc87d7cd82c0f329f247f ^
            Ied6c684cdd280b41ffab93a026d27282 ^
            I1ca188bcdebbf41d84f7a5220bd1d195 ^
            I9322a2a61900943075bbc23c72a3f65d ^
            Ie79c93f1703121713fb9401617f349a8 ^
            exp_syn[41];
          Ia3aba80aead67feab12e4800fef82322 <=
            If9a5d830e3ade0fd96b98f5949f165f0 ^
            Ie7a68c2b368a295f95571bc4a109b9f1 ^
            I0152dc6e6a7acd72a2144623e63998ef ^
            I9b560d9baf8a7422b0dd84720e924ced ^
            Icf25f076eec2bf81c899c66f6cfbebc0 ^
            exp_syn[42];
          I1181d42b560fca7bb5c924a81a5db1fc <=
            I7332e088bbff69db19c62685e033d26a ^
            I1b6abc8fbab3849b285e9f88a4fe867b ^
            Ic14f948884da19a272a4760ffaab9ea9 ^
            Ice5f7168aeb940d48093cc9df7cba36b ^
            Ic5c837a0556d1cb66edbf0294d08283a ^
            exp_syn[43];
          Ie4e5f3d7c5d2df30653f5666d14567bf <=
            I3600031716c2b4e21c9f577d34e033dc ^
            I859d795a7d141eb777c1f3c038203794 ^
            Ib9c194ec16f435a9357cb344cf25bdcc ^
            I69d82ab774d52c219509e993e7cc4deb ^
            I51ff4bda38746682e3cd4c68118c3216 ^
            exp_syn[44];
          Ifd9345cf219c58291c0b437aac093d78 <=
            I2eac5b39c6f485c9ae0bd341f894633d ^
            I12a18a1f8d4416e9bc8abee6ac3dacfc ^
            I45bdd0cfe107da0d57cad1333bf95e3b ^
            I768720af835b02a8dab376ef23d17a15 ^
            I1c074a53e6c0f2467bcdd7c952f51670 ^
            exp_syn[45];
          I4f2d7bb48918ce51efe6b3b12f9f8e65 <=
            Id3de87169c440f95d406693ef77cacd6 ^
            Iedc463e359dd3003d9f7e50f3e858e93 ^
            I23955b54e486f0f0d21a2809a9472b86 ^
            I24075f37c6bbd90c83370de1a2e58af2 ^
            I37c49c5a2af240496f5a5706b0d42ea6 ^
            exp_syn[46];
          Ifa612e6208151c616c3a0319182a96f1 <=
            I44daa5992b00e7af19adbee70bf01f2b ^
            I457ae11ad90c8478751eb4b42764e158 ^
            Ida3dd5e990ce3c237e9628a9a090901e ^
            Ifbadefd3a7ab50719a703400ddd742c6 ^
            Ia94c439131e1df5c95fc8ad3cfdba473 ^
            exp_syn[47];
          I9cb28a0cc6358610854c8f8d1dd3c707 <=
            Id88a7edf897eea1b4a137141789a04f5 ^
            I70dd1350d65155ee7b562f4c79024a3d ^
            Idc445d3f5b3b62562b0ac83e5f17e92a ^
            I723a6fee3b2496f23c48b3584f8bf9ce ^
            exp_syn[48];
          I40bcc924f5cf1f7d587aa35267022261 <=
            Ied638fee34f8baed4154b0b72e43a21e ^
            Ief03713f5cf37200373a20d42c7fc9eb ^
            I3ac0799861144b599995318bdade2114 ^
            I648b62fa0bc2185c1756ee531e8e34de ^
            exp_syn[49];
          I5238f7273b05b8b9f376314acdc6cc42 <=
            I1b43f29e0ddb72467befd6f3a9c1c829 ^
            Ic07c650e6e49892a41cfaf3a37471426 ^
            I4082b3564c1949a19ed35bd5a88e1ef4 ^
            Ife631f9a3c4c64a3d92aa9586ae75f3c ^
            exp_syn[50];
          I7137f56eeb4c4ae08bbc238db4cd3441 <=
            Id0f4dbb72da33748d8baf723c5a32567 ^
            I44ccc3ae897109dd51f9afeef93daca4 ^
            I73bbf90b625d56f663ad10f9d21d8e76 ^
            Iaac1d82f0846fce1bd88ebf8e60300ac ^
            exp_syn[51];
          I02335be013799e2560a98b6a82a0c528 <=
            I002820a37fa7c6c504c487df4368e2cf ^
            Ib0bb71b1f8829347b3a9a7543f9dd964 ^
            I1dd4671765f8826c2fe20c592c5e32c8 ^
            I3175159add7b814df637c2db8feb43f6 ^
            I48cd09f035f668536cd288a23010b07b ^
            exp_syn[52];
          Id327bb65156c8307901dfcb4184bb65f <=
            I76992221b1edff5684c482df7ac4693d ^
            Ib13436ad16a37d656d6b1ee95b9aee20 ^
            I47b0847946b0e00961233ac0101fa2a7 ^
            If2042aede3390bd208a281f0380c95a4 ^
            I119b2e5c2fea5338244c4019884af26f ^
            exp_syn[53];
          I56331cb7b310613016958553732cdf40 <=
            I3751f191f5009322acb7c9be4f8d7129 ^
            I14fa7aebb608d4a3d67176ba27d34d9a ^
            I7b813d83b13bb7bc13940cf5714c06ba ^
            I0eaa22f5eca8f33dd254fe241017a098 ^
            I2bd34b2fd12f12bc301fd0d5d69c0fb6 ^
            exp_syn[54];
          Ie3b00960f8af88a5aba7a2104dfca9a7 <=
            Ie517386cb5832e406fefc5e85eb2e7d1 ^
            I3fd0fa3b774d30a267d61e9427d09f3f ^
            I4ee312036de8c08300c358edcff1e1e9 ^
            I1d98943b01a6a2d8c4db18b98dd62f5c ^
            Ib715b1e0061b84ce614a30d961a83e7e ^
            exp_syn[55];
          I7d1ef47f35b7a4c3ea2e4383732de398 <=
            Idc07dc30c0a957e474546ac7a60df38f ^
            Ifc640243288c9b37b7eb9e00351b23f0 ^
            Ie83fa8157a7cce44c2e25f46ce897dbb ^
            I570c036d0237c53bb069c52d621e539e ^
            Ief8c2838abac83370fd7ec25c06d509b ^
            exp_syn[56];
          Ibb013f036fc42687a04bdcbe2d0bbd8a <=
            Iad90879acba3fc2101829549264960f3 ^
            I951dedd7af44c3865a8f36888432d0c9 ^
            Ia7606050c683ecefc510ba92ac539a9c ^
            Id3b089fb6edd5bcfdbca142fddd5ff89 ^
            I561d79eb079915c0b1732cbddb119c2d ^
            exp_syn[57];
          I77eae49d321f1d1e39dd7c75829aaedc <=
            I2eb08ebaa07a1004638cdd61a7209b7d ^
            I46e1047bca2b38e62b4de80d1d2249de ^
            I41796b587316c600bf583edc62649bd8 ^
            I0a569f6536789efb7ad2377c11842830 ^
            I8bb75bf828d5ef337fa6a965808e4638 ^
            exp_syn[58];
          I420a4d69a077dc1996ddb4b715d63e15 <=
            I47cbb92d2284aef7b9e56e88f0ba6f7e ^
            Ib99e1b93fb7fbda260d93eea3d24c3e9 ^
            Iee6e52d75c093a24eb4e5e0b45feb256 ^
            I19b73c5c93a71e90f620572f23f0e6d2 ^
            I11ba339c8250d07b497c88a39a6df1ac ^
            exp_syn[59];
          I652202a4dc8f102d29334b4811f5628d <=
            I8a4c1f23212ff846400651b100add502 ^
            Ief18a19d451f05f6051e3cc8de16d73c ^
            I7009c18515dd43d8dd2e5d1ee6779641 ^
            I173aa69cf52114e223ac1410d90b4bfe ^
            exp_syn[60];
          I0e33e0cdf39fc4cc99f6696e9f2784de <=
            Iada5bc4a51dc1bf57bb9cca11326bdff ^
            Ib6fbe376477afa58bfcc17a8564f78b2 ^
            Id48fe0672aa98f987162931527e9f9bc ^
            Ia4e89e99acb95f4183474b94798ca35d ^
            exp_syn[61];
          Ib9479328689dec62f900946e56ba0eb4 <=
            Ic1927bb3335f6a28c0816eba12d3975e ^
            I5b8a1e1a6b904b0f6822c224ee0486e3 ^
            I8be4711146486fea913843e497065b50 ^
            If4c36727ab1c29bf78f72e8acfc00d7c ^
            exp_syn[62];
          I2728682c0f749d1a9e8afeacdf44bfb7 <=
            I9b096ce09467c10f448496fda13987d2 ^
            I57b7b48f13436b19a8d6a47e014eb41f ^
            I5446c1c323774715371c73bd1be66697 ^
            I6426943b4ab66f17c2b7b399ccc7a6a9 ^
            exp_syn[63];
          I07da3bb5f943db6271fe1867a358df35 <=
            I595665d8128bb87ab62741d7ac520a4b ^
            Ic920452d5997a8477724fa78c86c0fba ^
            I3a8e9e7d2cd6751e8500a5567cef5acc ^
            Ib0dadebad37d9ea9d01350054872863c ^
            Iddcffa815489773b3688fd68dba18bd8 ^
            exp_syn[64];
          I61fc44808c85a75909b9d9fd4035f147 <=
            Ife0952b85f14a960007b67646b0cd969 ^
            I4d54dd2ee2f32909098d3cc2b6689220 ^
            I797c9cb725f88c07be28f017871d17f8 ^
            Ie165d0729542c81ca89f45d15e0afd3d ^
            Id00642563679fa9a6696f8e7bbdf6576 ^
            exp_syn[65];
          Ic5075ee0ad355c20dd45ed594f2a8c3f <=
            I258c45897919cec5c6acaddee7f3a41b ^
            I1e11f0088959aa40b4ad1a047b59caf4 ^
            Idce46f6d03376bea1ba361e8c59f8bd1 ^
            If17c0096ce34b88007247bf4c429d5c4 ^
            Ifda1c55899cd3506853cc82b450b3936 ^
            exp_syn[66];
          Ic0a651f45a502ead495cf14f97d65bfc <=
            Ic69094123b75ae36e3e54f179a9f2cb5 ^
            Id182a776b03f48fb139c28194ae7ab6b ^
            I65171c9ee8449407484e5c82d13c6751 ^
            I92eb6f60c14ee9eecb01718b01ea980f ^
            Ib5d1a7cdbcba0b654c12063d4f1768e1 ^
            exp_syn[67];
          Ic1c05ea22f708f620f626cc8c5ca309c <=
            I07abbbd75d91018ac53f53e64cffafb9 ^
            I4cdc955fa9afc75c2c977de4ec540e1e ^
            Ie79ce8adeef2c3c24a3386f054d0cf5b ^
            Ifc2963762403a00c4f3662b2863c991e ^
            I5e8ed024e2f2548bb375a2ecf1918a5f ^
            exp_syn[68];
          I61a18378aadae4556da501ce997321b4 <=
            I256050251d23250854ff337bef28e460 ^
            I20ffba20af04b99954bf719589e90d1a ^
            I7353ebf3a1cde89d2bb3fa667f7f5485 ^
            I97e82e5f6775d1e31537b891597223bd ^
            Id25deba967318f049de8163e67262f4b ^
            exp_syn[69];
          Ib1fc521709a1ce2198fd8df5b41d0177 <=
            If876ca6a14ffb4323503ed46666bc25f ^
            I5109afc4dc91780e05704ea5e1399e3e ^
            I621b20d29d3a9a9f41065bc3c3bbd2d8 ^
            I76fd9005abd511c3c5bf6c77de8bf2f3 ^
            I925f6b549a25cdc8f85152eb21ea3b58 ^
            exp_syn[70];
          I1bb5511c9cda1a595c45ecde48e9ebc7 <=
            Ib42d37576e3aff3d205f1f8822cc58b5 ^
            I3ce10718a2211184999663c3c2493cc1 ^
            I06b48093d4c9b0327c3efc6fa4ca7daf ^
            Ie8e29053f122a9247b0dec291c6ef4f3 ^
            I9b49e1acb81ef5b088b808d2e4ce9954 ^
            exp_syn[71];
          I4a29c37ed36b6e12f1f8e263c92bdbc1 <=
            I364ed3f83c49626bc3b939e53524d9c7 ^
            I8188dd7cb03854c6f709de06ff785d91 ^
            Ie7cfdd25541414ff3f8d6e5d7677fbe5 ^
            I6386a4dd26e7c36165dc265b3a2c93cf ^
            exp_syn[72];
          I4bf02a07719402890405fb2e7b679ed9 <=
            Ia659126b51468cfef48c97a135a71500 ^
            I866b30a63b3b5fb708934a1cbb0e1d9a ^
            I2b7822d5d77aaed61eee87570564df76 ^
            Ia20709f08cfff3a51d4af1e81d640400 ^
            exp_syn[73];
          I75bd82990cb60b6d7ccd7aa2982da7aa <=
            If1c0a3726041f70e508d68cbf6e40e04 ^
            I019e399a1cef87745e025a7d74e94db0 ^
            I0dccb8eaad52ce4d780696a8485420f1 ^
            I1ff042bdb52aac5d69791e96e2f9706c ^
            exp_syn[74];
          Ia6d3e38249f8a1208540b68f54c46769 <=
            Ice1ce5b4c30841dd92268559ebadafcf ^
            I3d149293f106ae8680c7f4702daa0bd6 ^
            Id17ada8dae3f9810d1892d34f2288859 ^
            Iaa2cbf59f6f61198b4fcf5a741cd5bc8 ^
            exp_syn[75];
          Idf548b72357ab28fd956791e84e5d65c <=
            I3eeeb1949945032d6c1759875426b733 ^
            If2dfcbf493b761fb5d7c622e739b23f3 ^
            I3f5053e519a928640ae49cf4e5b39d1e ^
            I01c94743a11042e75638ba6618356203 ^
            exp_syn[76];
          I50b6f2e0ef2831535ac8c18cd7ca9379 <=
            Ic2b000c3b2ca3beff2d427caab04701a ^
            I1c2ee281cd47a8414851c5e1c758ea65 ^
            Ia3ef2f70c5abaa852586a33c505aee0d ^
            I0a0340a0e52145f3597accfe4a4e8624 ^
            exp_syn[77];
          I4003a2515229ca8eb6fefa2bef289ca6 <=
            I3c3c22bf63e55a81ae91b1dd1ef615a0 ^
            Ib02268d5048c7c8e83118070e927453f ^
            I30be0b18e4415ca50f2d8149efaaafe6 ^
            I3bb4d24caaa0882a75125e466070f0b1 ^
            exp_syn[78];
          I48672f8b83eef8c406694676746469e7 <=
            Iaf36ce8598a29573979c683a5e2cf9fd ^
            I82f0e5a32d1bcd761a74f1f9ce8c88ba ^
            I659322a9fd0d5eac514437b02e0491b3 ^
            I44ead0ab5ccc53226fccc03024643771 ^
            exp_syn[79];
          Ia14a60c9497c0faf3f1f448ff2abe553 <=
            Idc2a9c6dd8d2aa912548c918c8a488f4 ^
            I08f22261d5713c0636d77c7938f592d6 ^
            I04c734eb876aa722e84d6b9edd297978 ^
            Iaded125f7fd5c833e7206dd7071069be ^
            exp_syn[80];
          I0ef3962dd323e8ec64c4a881bd4b3044 <=
            I98febac90cccb5fc1f3d966b6e38c4d3 ^
            I0038305f94aaefe2cd1a243580d95932 ^
            I0d41bef808860bde56d48792764612d5 ^
            I373be7c3f9511a2906584e33e5048abf ^
            exp_syn[81];
          Ie9b64c34e31dab63c03b3de4528d53fe <=
            I2c8f4a147b363d9c5ef0e080d9a9ed40 ^
            I9171019227f35760d02d0c8ce786f4d3 ^
            I669d34b955d2991ebbb31c149ad1b6f8 ^
            Ie0b5f51835ebdb508a596eeebf0e4847 ^
            exp_syn[82];
          I5941476ded9f6dc25d7394f5d133955b <=
            Ie644d131c4f2c603e8e64c5581fdf822 ^
            Ib70e99c3acc76286a6811bcacc9284de ^
            I263aad78110a1136eb7012c6983b2a8d ^
            Iddb75e0197b9a76b36a59ac2a7ccdf3a ^
            exp_syn[83];
          Ib46c78ff661ee6fb69c704d39235ffe1 <=
            I8e873fb2321eea82bb590a92411e2e2c ^
            I6cde57127c5bd2732e71ecb7738fad6d ^
            Iae6ed7748692f2edf1aa9d73380075f0 ^
            I08c03198b9599b2f4590e3022e398f7c ^
            exp_syn[84];
          Iadabc5abc7dfbc1dd747179ad7e37850 <=
            Ia62832d325f86160285c4d1a790a32cb ^
            I2f23d4cdb6f5f827513aa60266936e4f ^
            I4b99891bed4f5c149cd4a5b4f1dde0f0 ^
            Ia4f3cff223e24815ee1d86bf41756f06 ^
            exp_syn[85];
          I97a6b5f0976feceee3a5b5890d4d76a0 <=
            Ice82cfe55a5f226746e59e5c8beb46be ^
            I09031235f61238b0e32ff52641aab70e ^
            I9d7614d286377329eb3999213889b707 ^
            I56592e1452c4b559af19465b30230ec0 ^
            exp_syn[86];
          I7217d4790fec9797a1eb8cab1ebce71b <=
            I384d5377ee6b8f7eb2db23a2e444ddbc ^
            I477a920e2326828bf026b0a6b6a18e2b ^
            I5196382b75d16892d550f17893de15ec ^
            I213ce488e5345fa405a9c5df297d6f74 ^
            exp_syn[87];
          I3dd024db4130c105a6817e8a4935de0d <=
            I5ad7eb9d3ce7c712515254f892d1670d ^
            I914dedc1d5e5e21c9b8d07ec0ecc01f9 ^
            Iefac1e428116a797c2c0803410ac5601 ^
            exp_syn[88];
          Iae502e5a5ae518fb7b817afff28b7932 <=
            Ib534288c2cf976b6ec85db743bc2a823 ^
            I90023493600924a76d2192080cf6194e ^
            I8b419d5827e5b1af9649d602401c189a ^
            exp_syn[89];
          Ib8b2b1d90204af5b100379ecad20fc0f <=
            I485f9d1104a965d5d035feef912a2ca8 ^
            I474f6bd977f4197742d0bddb3bece684 ^
            Ie989550c9101de382056dd60d5da0e01 ^
            exp_syn[90];
          Idf0e651d0b13e167df3c0cc40d149c29 <=
            I9b76f0121a3f7e887e7121db50024ab4 ^
            Ic3fb524ab434e80b3289c9241b65d224 ^
            I259010e323e1e8dcd9dd719091131f6c ^
            exp_syn[91];
          I89daaca029498d05ca62c095db439eb5 <=
            I30d615203b697787ead37394953925cc ^
            Ic9146d8b3dd0c612073b70b8a8791e8c ^
            I3e0b41bee4c76eb5f3340ad23bfa01ad ^
            I389ac86954fd70464c9550e3fed4ed33 ^
            exp_syn[92];
          I0fe5a34ceda936d0924efdd07fad11e5 <=
            If4cb744ee52b6ae793431cd038069b57 ^
            Ic3cb34aae74c5f1a870b3635f8a40764 ^
            I877e8d94236c3d8b0a31858a98fba5d6 ^
            I77371f0e55b4684d1af196ed52d3d997 ^
            exp_syn[93];
          I7876cbb2b5d8aba3652ec8b218080dff <=
            I83c7d177eec2dad0a924557cdc91ba77 ^
            Ib1073489d63ea33d7f3892f4ff875358 ^
            Ieefbb5d6f4ac1e586832c5c0f513c5a2 ^
            I5a21996f5724a2a49fcf8e928c01b062 ^
            exp_syn[94];
          If692ff56ce90d22d7af881599c54df75 <=
            Iea1297491d1dfe98f395d8c73808a893 ^
            Ie9236599cea94cfb603c6b977fdbb44a ^
            If8fe5af7e5c3c97b5a713f6bcf919f1f ^
            Id46108963921efa50aff64d4dd7d1701 ^
            exp_syn[95];
          I18a7a4fe8931c79df3a69223af46c440 <=
            Ife25829fb3c5023b7d69bbaadf9cf77e ^
            I3375fff5ee0d4b4b12c5a70fbdee59fe ^
            I68c35d63dc95baff41b4dc27a86d2342 ^
            I8da50e5093acefb6f809aed64564a53e ^
            exp_syn[96];
          I8eec3538b8cc9c046954b6804cc656b0 <=
            If988b82b86db1f4ff6d3695f7b0197e4 ^
            Ia9f5ce4603af279bbd9b486b67016482 ^
            I0c5539373b3868d0664a92157b4b4226 ^
            I03b0694777d0160a83cbc82ac1397736 ^
            exp_syn[97];
          I653767e659590c1676edf6c25fc0e253 <=
            I10fca5f2cbf5e2bc3433c0dda579a051 ^
            Iaa1e981134f5a5c02983c49562683bc5 ^
            I6eea5fde8e2517554ad6ba25018572dc ^
            I85c2bffb93569d9fe1b1bcb10b98bcac ^
            exp_syn[98];
          I5ff863be142b92dff89f7916d0d088c1 <=
            I9eaf4e9ebe07717503ff69b51f0e1905 ^
            I23c8b64e433af0bd00cef44e38df99f8 ^
            I7bfb4c5d9e22d1bd8811844d9c74dff8 ^
            Id00274c88b93867a80606343add1cdab ^
            exp_syn[99];
          I49f9fd0e0719be527f2a54814dab83ea <=
            I7741e239c16828889d488cc87647c154 ^
            Ic828cdd5dfde844df4c150921af2a443 ^
            I61e829cbf7d6c0ef8ddc11677981e2cf ^
            exp_syn[100];
          I945f2476eb599844cbee0cd89038e392 <=
            I7050adb9d06f767549b7f35c4679e391 ^
            Idc5fb0f3a04ab32948e249e088a11b11 ^
            I9e8ae2aed048068b01b3bd46f30baae8 ^
            exp_syn[101];
          Ied0c5f8a9243cd9d93672ad6cc907d21 <=
            If43dd31198c8a0da6fabd194cf13bb70 ^
            Ic0732810fd355d59a3168be896a0f9ac ^
            I7dab71adbe62687846fc027d2789451d ^
            exp_syn[102];
          I9134c7f579723c7615af60b4344efe76 <=
            Ib16548d471f0a4f4625852ea04335dcc ^
            Iff2f1716cbd73b406d8f07c22dc79fc8 ^
            If1295608bd218ed60922a0b95bf1d098 ^
            exp_syn[103];
          Ie92388a9d1e71d73c07ed86e9bf6c887 <=
            Ib051eb1091a85f85a1e50007f1b27cab ^
            Ibdad0ab78e4404c852e60a2b04c3a5f6 ^
            I5fdd8e1550feaecd81b82069fe73ed7e ^
            Ib4ae1cedd09d72c235765a6cd7e91366 ^
            Idf04e08c120ed116af14a62659675b44 ^
            exp_syn[104];
          I6804fecdf59233c6cf14409bf2f1e430 <=
            If6a5dc79c0f6ce348956286737a369d8 ^
            I6d4fc81ced37c159303c243af04d345e ^
            Iba1c0ebd9cefeb0dd7f690bdbbbfec58 ^
            I3472ee8c06644490252e606b62bf9bd5 ^
            Ieb7614ad1b1bfed3e2b0089a72fe214a ^
            exp_syn[105];
          I9e777a342bf53eaba0280737ae404bc1 <=
            Ia8e304ca12c82e41cb8e4de7be199394 ^
            Ia2c5fe53cb5b318fa63d09881609655f ^
            Ic124975d36a292816146a2fe61ab3ab9 ^
            I3eab1582cc42db0ac7739386cce2a712 ^
            I589062eca318b25dfe5735da455b6fe1 ^
            exp_syn[106];
          Ied53820aab06b5c3423b1d878c71948f <=
            I05721e06a1acdcc0571907c7d853f18c ^
            I1e93f0470d2818249f1c28ef2a399a0e ^
            I453dd7d7c0a2f003f0b67e909630d641 ^
            I6387919f2426c283e2d70e471cda54a6 ^
            If3db87afb3ea184c9e4020c5e45cb161 ^
            exp_syn[107];
          I24cceded372d782c67b33f3a78b16045 <=
            I7979161aa1e2262ebea862004c387697 ^
            Iaddc1f2e822fd2fe9d9046d759a82cb4 ^
            Ia14bc1fcd5bbdcb60b8e68298f7d716a ^
            exp_syn[108];
          I2e78d36bca5bfb016af674c343f9c041 <=
            I04aacd95d9e44657f616e01c9053f0fb ^
            Ia8974083bfd064f2c27dcd421490fcfd ^
            I268b60cb371b3d46dc3f8b0009f541b1 ^
            exp_syn[109];
          I17a9a995de58643dbbfb78604f26198b <=
            Ibeb8c72b90b50c6897224ca1a792fa56 ^
            Ie232799bd6c4ec99e24c78f3ad798265 ^
            If2cd93b57cd1c2b91ee7a73a97dd19f2 ^
            exp_syn[110];
          Iad642c4c62766e8f8bd5a1e9e73bdc80 <=
            I0987c561670b7b2b6683303c1be39561 ^
            I3b30b4ab00a49e10a75587aa324d6132 ^
            Id81305359a07db527e49fda05cd2784f ^
            exp_syn[111];
          I96f92481be1ac6cf985b8ab387d326bf <=
            I8b2a79aa4ac88e6b4ca8188a7852022e ^
            I6b5645cdde4b35a16fe3e91d90caaa4e ^
            Ibc48fabc172f27ebce18d0a9b5120dc5 ^
            Id8292eca087c1a17dc8b5a572a76f21f ^
            exp_syn[112];
          Ie03c09039ccafb427153d2347c1caea8 <=
            I6ef260ef75e47b011a46ba2080ac3684 ^
            I34e6e9d2153e4a70ee36ab85e72d5318 ^
            Idf1ecab26889c4adcb835fda6b1cb368 ^
            Iddb19725b093506e5e521d8d68dcb8e1 ^
            exp_syn[113];
          Ie7381a8294b4cdf669b9c57cfe4012b5 <=
            If8572800d5d80cc92dd917b60447b63b ^
            I3566f2779e860008b1a5d305366a07c9 ^
            Ia9f1e580e8f441394d719d52a7bad688 ^
            I0b573d3a86a3111451da661e46384876 ^
            exp_syn[114];
          I61c9e3f8e42f869f4c9c1386325100b3 <=
            Icb0841ecf142687c3aa23e68f01c927c ^
            Ibfcfd3151af0d82bfce293ada44059b3 ^
            I220e32641265b46527ca61111f7ebf1b ^
            I0ff479e61d1a0cede88ebffb073c60be ^
            exp_syn[115];
          I24c5b2de59eb1f43fe1efe687231c4b7 <=
            I8e87530a131b5a73cad6df68b9e4967f ^
            Iee17ece482d04964d3c21a092ec955a4 ^
            Icd6f8f5df6b4ca4c81855e974db76526 ^
            exp_syn[116];
          I43d43acde5f831fc32b7bf5f10b9b3a9 <=
            I2bdf4736022e5da7294a0e851006a124 ^
            I1c7e41b9cb1bdb6f649c88c0ed3f4100 ^
            I7ce064a756dad56d37684d5d7d168047 ^
            exp_syn[117];
          Ib06e93161fc8ca3be232f4261b04feb1 <=
            Ic62fc602da3d16fe13d03a49a21269d0 ^
            I5364deb983adc2ae505ed2b8c57f876d ^
            Ied2ea62cfb21602645babc36e27b8218 ^
            exp_syn[118];
          Ia0dd00f83afc805036f2c6a0e38f725e <=
            I2ff317d57f59747c4524ef4278d51092 ^
            I6e92a48aaab94074a555efa9bd1e7243 ^
            I79b85da6e5ce0b02ebd1619115c98e24 ^
            exp_syn[119];
          Ib0a0f924fe3757a1e0aade7017ad9277 <=
            Ie68b31360c12a83c6095254b6f14603c ^
            I00d3f14b20e1ea7d726533386e0eba27 ^
            I579c7926e7b78f4ffc606adc10522f53 ^
            I837183265ee22d080e81fea468ab0887 ^
            I8e1ddd7e4185c28caa71d30bc28138f3 ^
            exp_syn[120];
          I1ca949071d734d230cdb8adda46c9d79 <=
            I9539fcc40d26b13015a864718b116d5b ^
            I02849282dd1bd663fd39baccf41762f9 ^
            I5d6e576b0fa7e3219aaf9ccc345085b8 ^
            Ic0191941cb968bbd7644c21767423d2e ^
            Iab0bff1633e2f3ea0bfbc291f3ab5d29 ^
            exp_syn[121];
          I40170922c652fa7fa42abc6f580b5e3d <=
            I8850ab26807dcd55fefadf6310729ca7 ^
            Ice59d2af73d0b0f2ae91a2ef0c2b7f04 ^
            Ic4efba3932e598784f5b9ad6ad04772d ^
            I9ad2f6fd2d7f68011fc926ec9abd5c34 ^
            I5f0751fceaa008feba5c6867ced453dc ^
            exp_syn[122];
          Ib1ad0b531ac9028971d68f533e7ae566 <=
            Ifdabf743a8cb46b7053000ff48ea0c60 ^
            Ie562ebb336e476a81f20a652d4cb20f1 ^
            Iefdb8bd28839af9413a3906cbfe715e6 ^
            Ib9d58222da98f29fa302b4896594fe26 ^
            I9f6751c15237c20b0cf2175575195ea7 ^
            exp_syn[123];
          I0ab0170c7ceffbb58377b65d2ad92093 <=
            I081e2595b18f306a74d070203447ecf6 ^
            I3b84dad6d0dd8730312b3e20c6d5a2a8 ^
            I6ea50be10bc990a1206cdc9e28e0c4c2 ^
            exp_syn[124];
          I9ac68f228a93bbf4aa4a559b1364e42e <=
            Ifc1da524e7670772834d521a6fc4c96f ^
            Ie2d946edaddd3c87f328e861f3e72c0a ^
            I43c2fab87f70ea883321ab82de85f133 ^
            exp_syn[125];
          I375c5f7eac92d853e85e0606011f3fb0 <=
            I24645082ef16129eed1c574f5fc601ca ^
            Idb1efe99b5d7fd567a7f82cfd52f7eb8 ^
            I1af02ed6cf00d4cb0704b5e44c83bfa3 ^
            exp_syn[126];
          I94f9b1f2e63748c21ec7222c9641366a <=
            Ie8c0fac00a9de74870e59cbf9e87a39b ^
            Ie4827dc0983c1a63053c08de6e36d375 ^
            Ib71611afdd0381cc1884f5ddbbae1acc ^
            exp_syn[127];
          I55500c1d85c4970932be67cc5cd2e023 <=
            Idf8d15c7bd7705b9aafbda09c3a5b46c ^
            I7f720a18542528f0c9bfb14f699ff4da ^
            I70a4926e9e6a05fa9ee51a26988862fe ^
            I38fc49afce0298846ae8ed63ae715e81 ^
            exp_syn[128];
          I36b487cd1a57a3a503e587fdefbb19e4 <=
            Ic6fd9592d2ffcb8f4ca83c6f0bd19975 ^
            Ie4cda4648f6ceb76b8fb74f290ab6439 ^
            I5707d30ca29842b6a96cfaeb44ac6668 ^
            Iddc3e44d83e8253e5129b6cbf5082df7 ^
            exp_syn[129];
          Icb5350e8c55a2adb370078a7575e28f8 <=
            I94009bb7239be96243902ab0f0abea7e ^
            Ic308610ea8bb62ecb6094192e02dbdba ^
            I85654bd3a07b4329aba17d8b27777f4e ^
            I975a87bdda30c5b6be8d2f0e4b107450 ^
            exp_syn[130];
          I8a7a31327c9e4cbd88ce39fea8971caf <=
            I8bd2a9d90074500698b302cb8db7f03a ^
            Ib5ee5a6ffc45ed1fece0822dc4619b57 ^
            I235c3a9fd3e8ea1cee762c10bc8e2c53 ^
            I582bd96afa764ded148202f738b7a1df ^
            exp_syn[131];
          Ied069655ed3775819d0bcb722d6d0488 <=
            I5490039998187a1a2efc3549e3dee7d6 ^
            I0615acb0f7cf79b5f6ae8e91cb525dc9 ^
            I7ec15b73b2811b44e1e50c74a9f921e9 ^
            I6fb88d97bc9ed37a06b729020a1df140 ^
            exp_syn[132];
          I78a5fc80d42e8db1b56cce5f4c97e325 <=
            Ic5cb81c821716a8aabf8cc2283ff73ba ^
            Iffa06a336949f56f4e5a88a06d8b7e60 ^
            Ic68f500938d80460ffdb33a0adc48298 ^
            I1500943c4a550e78fc169437b0a663b7 ^
            exp_syn[133];
          I3ade7e345432319c1a9c91d4068b3ec9 <=
            I22f5bb821a2571d1764978fd76c8f1d0 ^
            Id962beade26396738ba0e97f67d5e261 ^
            I7c965c047d862c973d09a81abe03a845 ^
            I0b83f4ef8ba9badb27e81b32765ec5b6 ^
            exp_syn[134];
          I88aed46f6dad7a81006562a720670654 <=
            I42ae0c42360c977b35429ce290516a6f ^
            Ia03836a4e93d2f36513227d1dfaea0fa ^
            I6d423a7d17e05a3c597ec6ef6c5a7cba ^
            I2c420acf428e44cdd9ca9998e276f258 ^
            exp_syn[135];
          I79e574dc9c7e18b695c9a2619b71b995 <=
            I14bf11ad80890227e47fda26ae1b9c24 ^
            Idd474d80b50992537d6f527faf279800 ^
            I2eed3d32a27d51036e17c4a21382b4c1 ^
            Ic7b6dae3017b55dd3cd27423d5f1b0ec ^
            exp_syn[136];
          I800ef583bec1d46d3d4ffdea6b312ef9 <=
            Iae7b72abf4d3c536330a229e3836b441 ^
            Idc5e98f6958786ccf95d39b922b42ea9 ^
            I2a4bbedf880a9a7b4e1bf946f9f96c0e ^
            I4a91a7c9b2a0f3552b8f2ef4e2398be2 ^
            exp_syn[137];
          I56cc5cd6d0a5a4e4601fd48e838fdaf3 <=
            I3b8cdfb1440732ce98cd1676e05a2af1 ^
            I3fbd40faa4c3b78b547b8348c466fd1f ^
            Id6b508145cd21ba088ab8fda34577c35 ^
            I99ff29c7ba68b5d0819f1e1bead51287 ^
            exp_syn[138];
          I21047a3955b8b89bdb9013d571b2bd0d <=
            I2aea17846a53e2eb2968581ee2c48226 ^
            Ibf2a253afde05c905d0b2404c5a808a0 ^
            I24f82a3f2c0e8df486fe495dd95cf8bc ^
            If06b00be0356a2be5074d958ddcdb2f9 ^
            exp_syn[139];
          I56eb529a34b484cd20e29958cd6878eb <=
            Iae5d6faac1f5685cb1d400ee2b1d85e0 ^
            Ia98a6f01e4eb5bc74d50d350e79be426 ^
            Iabb01dc9980b4879a7356712b51df0d6 ^
            I604283449f13c7b225ea03f99f2e296a ^
            exp_syn[140];
          I74588df6399af2c1112e3fa557e89e17 <=
            I68b152a599887c0039dd9d45c528c219 ^
            I24135210c23b2422a42c90ee25594191 ^
            If4308ed204e33952c9931f8fe257aca4 ^
            I2b600e5f5c146ee97c4044c08e1f5ad5 ^
            exp_syn[141];
          Ic8eae1a92f46db040eb22d726c3a0e6d <=
            I852d5295a32984af00c95f6d9389555e ^
            I33ee415d85e2bcd8f975d34b880f6ea7 ^
            Ifb89e7ad8ef661959d82b7c22f187243 ^
            I9fe16403fc21bb1159a5e0305fd1ef69 ^
            exp_syn[142];
          I854a15bc7e9728b01c9a1960f6248dc9 <=
            I207a0f6184a0b3be71766a8b47ea5535 ^
            I86ba73ee348f80e2f9891d2ebc8a02ed ^
            Ib6ae81df8db1dae269437861ee11ec0d ^
            Iabdb9374e5caee281c25b003624b2c4e ^
            exp_syn[143];
          Iae332cfd000fd0529684ab787041b5dc <=
            Ie5d9cc18b2dd300132470f206452ff17 ^
            I1b695aa715615662eff7065c742b0859 ^
            Id0ab747d92288f23cef793567b2363d1 ^
            Ibd12036702fe60b57354b3aac921559d ^
            exp_syn[144];
          I70148fe95244eebf7f0ec953703398de <=
            I671de3d408b5b783541663c7f1e3a6fa ^
            Ibe01835305315fab50269c72ef849b61 ^
            I138fb0c48f2d27e3315e237d9e61d653 ^
            Ib1639811de6eb1c38257800c201fb704 ^
            exp_syn[145];
          I24ee2d953e65fefdc73b3d3c4c0ddd05 <=
            I169d8f2bb5fde5b202b4239b7a7f1ed5 ^
            I2b97a79c90f6578c8b2f321f8d598cc8 ^
            Ieed4c810a5bb69de112522dcf00b16ed ^
            If926d98f659e8fe4bbf36ad2c5c852c5 ^
            exp_syn[146];
          Ie3a5f8eec283fd4f682b5d0f909b051c <=
            I8ca17b6cf35e1b1f8f601604575d3f27 ^
            I9a6923c6368526a53ef70e16471386ef ^
            Iaf82668eb49248709540f2f529f1b3e4 ^
            I211f8d7f97ebb8eb3e50313513abfb1b ^
            exp_syn[147];
          I781d986d7fd6c2fec3a8cf3f29545174 <=
            I0fd2f706e374a4eb57ee26ab50201e15 ^
            I83ecf12f3b38fc14c3b75e47b71ecc09 ^
            I304ac9f96945546cdf1b6f1fa7136731 ^
            exp_syn[148];
          Ib4db8131350f8605e00907234aff901d <=
            If5ae6fbf843fdeee17945bc5ce81aec8 ^
            Ie039ab562e9cf90289047b5425186123 ^
            I7a9800418bd5c195fc47a72370680b56 ^
            exp_syn[149];
          Ie093f0750b60d3aed75705637933f34c <=
            I9b8023f4dced915cd52c91bc9d4ed78f ^
            I49d35ec6369de10afb15be8e0cf135c3 ^
            I5f6a61c9f0c67510e148e596f553a4d6 ^
            exp_syn[150];
          Id2fba7c1b3dc7a75a5e0d90494d56962 <=
            I48e3309c61918c3991852b45d9c72ea5 ^
            Ifa6e3541f5e12bf9677ffc51d0392749 ^
            I8e313ceb21359bcc44114ab217b1c394 ^
            exp_syn[151];
          I9ecee74c445711a376133636ef414666 <=
            I3c0a621dbef864fd1f566bc2e47f32c6 ^
            Ie61f299252b8fecfd3e8634b64df5a90 ^
            I33ddee677715877c11a1df45cbfb01ac ^
            I4c9518755c33d725221ad79ee6badba9 ^
            exp_syn[152];
          Ifb3cf6b88835d27220df837682c4dc93 <=
            I5cac08dabbb6de3b01c821d4db93a8e3 ^
            I1e96d5af3d0e3fdce39530dfd0131a7d ^
            I373841aa2bcbad8232d54ac9035a3ef9 ^
            I3c3cffec9f47c9979cb9503f222f370c ^
            exp_syn[153];
          I386fbb3bd550891d682e137044e8773a <=
            Ib62b02ddf0f57bee49838d19783ef6c3 ^
            I182b43872d50de6f7afb700f178b160e ^
            Iddcfab4a7022e0f12fd20cb34e9b9d02 ^
            I68d6769541fdc3df321e192f645c667f ^
            exp_syn[154];
          I7ede7d2e1c2730b3b71340b11e880f5b <=
            Id051f1d5454802e0eb37e22248efe8ca ^
            Ib08897f9216599042f7b97b137e07fe1 ^
            Id1dce2b9eafc35fa71df33ada4aac539 ^
            Ided55428cbb77f454c2607ac783d7548 ^
            exp_syn[155];
          I64c65fad4a7d958d625c783626808175 <=
            I275cd09649a750edb8ae8313e4e1e279 ^
            If533578cacb685a95afbb8e1c05d3c07 ^
            I8879df010bbdf6e5fc9370e2fb3289b4 ^
            Ifd3d4f3e2a388b3c70e7704d6351e0ba ^
            exp_syn[156];
          Ib2e0cd0a2b51c3a265bdd20834c0ed2d <=
            I7c791c854d0bc28e8dd787545f8fbda0 ^
            I90b3708abdf742370f06cc513ee307e1 ^
            I9a403c511fe2d44472ab319a9477199c ^
            I17d32f292758416fe02527dfd938fa0d ^
            exp_syn[157];
          I67be0b66c8d0680eb23290a4b3885af3 <=
            I446857735e680cae93a24dccb59b1924 ^
            Ie536879e6fa9be65376d7f00e0fc40d0 ^
            I3ade5535a79ce83857481ac771cd8618 ^
            I9ce3942aba354c1fd7d6b9a39c994d7b ^
            exp_syn[158];
          I01148401f7d058614dc1ae6ed3c8bd94 <=
            I40a223380fb4414a3f26a08cb90025ec ^
            Id0b1c46fa4caa63a4c63a44ba3c5ef8a ^
            I88a89b2d938552458dab9bc34728959b ^
            I2c6c6041c9c69c84f4d64af6458955f5 ^
            exp_syn[159];
          I3394319c370daf6102be00d938d55769 <=
            I0c616f736879c28a5222de3d6f49a587 ^
            I44f170d02bae7fe044456e125a98451d ^
            Iefbdf686d9452a62cb99cf023a4d9fe7 ^
            I830a4fffe1244e071eb82c28ddc4a308 ^
            exp_syn[160];
          I24d6a334dd15ccdea558f32cd029e6d1 <=
            I620b8ecdcaccc1ec80ebcf9fa6af0017 ^
            I94460b6ce7b776bcc5eca149eab80c26 ^
            Ic3ba4531855366e9a060cec1c7694844 ^
            Ifad8e46fc3844bbfaf434a14f6b5869d ^
            exp_syn[161];
          I3a41f68bca2d7edd1f5738c4fda8e73c <=
            Iec91b3ca3b54010755d57f8b8ea4a544 ^
            Idc6b6357741c9887a9db1037ccc2d922 ^
            I21e72a7e5870151c3247d15121e5fb4f ^
            I10a6c6a8fdb0003de1f360c148777d0f ^
            exp_syn[162];
          I9ef1784d165492f3482d14f475732451 <=
            Id806a2df1c4519bbbe811791cb4072f9 ^
            I472352e7027b9df2fa957d9fd68443ff ^
            I74cbc0ec3bb682e0f927890eef8d7a58 ^
            I4cde586fc28f8d03fc9934d56f7ff7b8 ^
            exp_syn[163];
          I9d9378337a77515a4e8d04fb88938808 <=
            Ibd59d0e5a062f149bd0e91ba76985a13 ^
            I51e14ece9ab6607f83e6ba27f3f046a9 ^
            I433dd5092cf1851cd196feade3cfa6d8 ^
            Ib83a067fb08e118dcf794902beef9405 ^
            exp_syn[164];
          If0e20ef9aa69b77ae0e58ca3dfc9998f <=
            Ic4c6f707f461cebbc4c93f2ba664ae7b ^
            Icc67656ad2dd3fffae4e5abe02f8fff9 ^
            Ib6124faff821158c6a2c9a9c454ab68c ^
            I358cf9609272a4562423a85f9b2f56bf ^
            exp_syn[165];
          Iec2cb48bb1b58f268bf164d5e8a8120f <=
            Ic04828ba2db8239b093043c27476d345 ^
            I38352b363fa37f6f822fbc1a39100968 ^
            I759409e242eaeb144a53e630a8cfd514 ^
            Ic1e9d9113150ad57954c0e369259dc62 ^
            exp_syn[166];
          Ia4ae7c98720d43a604f28dfc5dd67d50 <=
            Ibe6b8c57d7ff47b6fdad5fadf1f6b841 ^
            Ic9b72b2a91d951cf08cf54ed215ecaa8 ^
            Ied19cb51636bfb029ba8a2c390f97105 ^
            If7fe3f5ccbb5b279e41fd183c8ff3974 ^
            exp_syn[167];



          I5033323484d90d6bfbe03749019fc6dd <=
            I1a632a3e06ad738d5865acc77e204f48 +
            I71b93abe4b20e6a17ff17e0f33ac2ca5 +
            I9184110e3e9b8614460fc0abe5fff2d9 +
            I535cad8c919a4330257eb5b4bed61b3a +
            I7ea8fe50c45e213f3257060e2813240b +
            Ifec9abca21cf476b70e0befa3926b46a +
            I7c191c2c2be09886d0f31e4368797afd +
            Idd01d014f0469f893305057ae3f4cb2e +
            {MAX_SUM_WDTH_L{1'h0}};
          If5dad13ac41b3034bdb034bc86c9b348 <=
            I3f59174b3764a0b0741462024be9fb92 +
            I0e112f1d4e9c934a118f79f3856744a9 +
            I65708fb59e90bb79b8107da619fe63eb +
            I0fc42ce9cc31d781ea3013318c25a571 +
            I8bc3210e86a523accdbeefe7e72ee4fc +
            I597c3f5c14e235f90dc8c796bc3e931d +
            I07d68462362d8453e83570cc793c55db +
            Ife6be241bc50560a14f97650e5cc2959 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iac428f9f798618e1ef495c626c41892b <=
            Ie04ce30f26a4ef1ee5b34474368dbac7 +
            I546657528d591e8bb44c32fed7707af5 +
            I0ace1d51fdee91f8f3826a945c4e66a4 +
            I8dbe6497a8deabcc60783bfe7548d0fb +
            I9a57f2f03cf8a154c3a7d48ec089306d +
            Icda9a86a25dbe516a93b46fe487029e3 +
            I64ae3cd6f36b8bde29cd3e1fcba7bade +
            Idc4171a40dd2470e852af37a461013c7 +
            {MAX_SUM_WDTH_L{1'h0}};
          I5a6427c8f18b36d2ea18fe60a0831ef1 <=
            I43864225be03ea8e9379eb28dfa6c599 +
            I70e68beb262fbdeba621b3794adf9f84 +
            I656852be6f5b3542862e0f68d48be518 +
            I041f9455435bfa375395eb330a34993d +
            Iac48d2ccf6c6e0c555e874ae77123f2e +
            Ib76e892d1a1271844338042381b5690b +
            I45b64b2b963963d2d0a8318133941f1d +
            I8435e69bc1ff06e7edfabbee7b9aa49e +
            {MAX_SUM_WDTH_L{1'h0}};
          Icc29441eac6ca7a138d45743d37505e3 <=
            Ibfee0b4ad5cdf16e88fcf469c5e031e9 +
            Ib2afdf9534deaae465d99b7e377788bb +
            Ib6cdbbb765694d822639b7c8fbfc50c4 +
            I8dddcade21ad3bb330c1c25970c32b73 +
            Ib63574478126e6ee30a388d9648cb548 +
            Ia1aedd38250e76763aaee3de2f832b3c +
            Id5ddf5331aba567aaf5b7eb88b31a52e +
            Icb158c031d434cb419c15e0510511231 +
            I79444eef1875b6ad1a0675b66392ff9d +
            Ib88c884e54d6e6ecf5ac015bc304e4f3 +
            {MAX_SUM_WDTH_L{1'h0}};
          I0e7754dcbc04a4850e052ae4a2fbe328 <=
            I31cb0c699cffcd2fedfbed0e1b86490e +
            I4363ca6b3d9ca9863f70958aa7c23777 +
            I25eb943ea517a4827efb1e797bfdc4f5 +
            I490996026af34eba5bcd8d553af818eb +
            I9d8f8c1792427975a9e7024041f59be9 +
            I452ba61d5fb5c7ead1824dade4bd7801 +
            I7e36dcae438a712fca2320117b7e3356 +
            Ifc527b6af9486df7f52d7eb9637c671f +
            I1062442edb2bff727ca6283c8270bf28 +
            I2959f2dc554e599d675eb6912757e413 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia30c019ed8ce395556494a92e7b42a92 <=
            I4d4ec5540257040d10182ed478a71918 +
            Ifef870b405335975988b58b2273d4e1a +
            I9e0a36d0be66b4c02b03e5b75b686226 +
            If404a00ab81d6ebbc0dbdf4aecdce389 +
            Ic6f40833f5f6284c9015304fd3fc00f0 +
            Ib8664a2abe9d6326d6e45bb2a7ad59d0 +
            I36ed1a0d0d618f90443fbea17b7c97ec +
            I397a69dab323c7148b620dd6fe0b0c51 +
            Ifae488cb68d95ea517376319eb11f1bf +
            I10f045edf47784a91a5599494c2d3de2 +
            {MAX_SUM_WDTH_L{1'h0}};
          I9799695ea8244992a6694eaf5c8ae64d <=
            If0c2d002c315b21e11ae776bb48c9338 +
            Ifbe29365e7035c78af9f42902b0d303e +
            I6922b510e432e06d209095bcc6297e7e +
            I31bf4597a3b776962f5c820378254065 +
            Ic3e6e38a2986c7f14fd0db2246367a1c +
            Ia1d9dee7a9821283498d17de0cfacb32 +
            Ibac0851ce1a3c23f18b072d263afff36 +
            I53971b75cbd7ebc74b579776a6ea4778 +
            Ibeff607ba15fd8ef504224a9c1d102fc +
            I4ae2f2330a8ee7d5626499f2a030c7a5 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4524cd664b4cb41f642c675fa484c84b <=
            I8da7e01f56dc9a70eb6b3f110dc005c2 +
            I005e8b590924f9486cb23191d35c9797 +
            Ic1f6842b4f246d624d91daa6ada10ca9 +
            Ief90f8a8efca2b06eff0d4cba1cbb342 +
            I0f46a17f14ab18e6338aa3d06678b0a5 +
            Ia3bfd86e26efbef2cf6bb72be7ac1453 +
            If6f5efee5e1f9709d86bf28cfb741955 +
            I60520c850a95b893528569c4069bd677 +
            {MAX_SUM_WDTH_L{1'h0}};
          I64e959d80af111ed2fcd54a5407d21bf <=
            I18e548b082364c75686f2b7ad2ef46ab +
            I6e4ae763dc4e8aa8afc4599de96c75d3 +
            Ic8759e2f58848b33082bd1b02acc9c0b +
            Ibdaa6d215d34aa0cc27d5234da6fd991 +
            I0f9bc36c9d40290f83489aac3d674924 +
            I9a2bba3f62de5f750dc8161a488dc331 +
            I898d1b59aab3d5d4adce8ec3c0e14a0d +
            Ic92ab3dac1a151d6ff0b4e0c21003eb0 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3e0da4bcbab4804b5397fb3aa2c94f51 <=
            I3a4a965f22487553dec2a3e8e7836264 +
            Ie7bf11bab3d601fd0a6e3eb415e263c8 +
            I6eaffd980e4d77fdbda5e63bad9489d7 +
            Iac4b8906947fc90bfe76cee2f1d4c4ab +
            I612a41511db375f10f3c2b10d13edb24 +
            Ia6a78664c080829664158f53ba330312 +
            I6a81b4485598387e4656c35e83866209 +
            Ifb09b84f9681c7bc28ffd562b633ffd9 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3740b30d31f3c61d93a14a46e3199c4d <=
            Ibed5004d869a01005768ba694c2234d6 +
            I91c2f3cdd7cc98a60090ec6e46d52ae7 +
            Ic902e09b33db1b919c102f7971cdef7b +
            I1eef40a71c8d1e2da9802929a5347e90 +
            Id58474582f209a3859f65a447fe99191 +
            I1939152ddbede923cde577984e0aa743 +
            I4aa98503fc71292d42dba1cab6db952f +
            I8ce945d9f70bb317064a8d2d4eafd2d3 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibf0a30abfec9031737eada436ac1a0d4 <=
            Ica3d4ebff001fb6ee69a66eb898eb5bd +
            I99ff3922e018c409dc8ce5f3503e3c56 +
            I58a490344f87b4d5bb319e3e85ba9278 +
            I58361fb97f1b5aff0a2751d35c8da672 +
            I581eb136fdd08302e02c1fafb5d5c90b +
            I91893028c4409cfeceeb7976815b2d31 +
            I19032091a26dfdfffff60818041ec79e +
            I563802213afb6abe2f6e8c6f4d1e5b08 +
            I4ae59dd2f57bda295e11b077e8668f1a +
            If525ac3dc97e3187e036d70e9984939d +
            {MAX_SUM_WDTH_L{1'h0}};
          Id36e8953a02400a5ab1f4dfdb0422e6d <=
            I4254f2987cd014ed703ae18e9963e585 +
            Id6551b6b053952162b90792ab73a1a49 +
            Ied41909cd443432dafadba42672151c1 +
            I74a7b85ddacad06ab1c6b0db9b084bd3 +
            Ic4501a8a1fb34c30a97e18a0ab189e3a +
            Idd8643af2515f65fd9a1dfe66494ccf2 +
            Ic9e06a355beabfacc053ec48f17f49de +
            I31d94aae2e3721045fe850d84dd2225a +
            I71da7e172b2b967040b6e6d02ef9949e +
            I3da241c7f221413abfbf1b4384bfca5a +
            {MAX_SUM_WDTH_L{1'h0}};
          Ica71108a53bfcfd1892b4d03ef68110c <=
            I8c5f98353b5b082dc3cf056469945a08 +
            If8865fee7dbf593b34ea54692d947f10 +
            Ib5334df42ee8f1574e41cb30b903fae9 +
            Icbc12ab47f586b12402ae5d4361c967d +
            Ie8644d7edbadf19937c399cf275946e5 +
            I2087576fbc15119bf5d9e8afa2603b69 +
            If1ec4241fd12255369f72b3f3310b6e7 +
            I401ab1ad994f5018061a3f57d3a51ad1 +
            I2ba16a10a82c20d54c776a9804ee50e4 +
            Ib55b0e4c45ebbdb605f0ba9d62bff21c +
            {MAX_SUM_WDTH_L{1'h0}};
          I7c97629ec6e594f9b2160815ddd133cc <=
            Id8c36004ae8e550569a491f6b514945a +
            I840a1a7c0bf49f4f42499b33f32fa02d +
            Id769d4a92f5f6da262ce0521e5509368 +
            I19875f52f79482b477f1febaa7e97090 +
            I3f2507530dd648814af0964f7da11d35 +
            I8b5d10c412daccdcb07645bf239d61bd +
            I3a09554ca009781e28ef1b3ea70d39ad +
            I37e5c3118e8536e37bd797aeaa92476c +
            Ifbcebda2bb0ce58a0e1764c392a816df +
            Iaed105b99eae5b078521e3a94d8a79b7 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4823c8239ace86dc399e906c1b5a0d74 <=
            I2a2d014f94d7a3b9fb3024a3e9107a73 +
            I9aa11f30712f1779339b985212a7979c +
            Id15c3bdce785df234c68432ccec8f959 +
            Ia0e77e9544481aa0f56dfdb6eb253137 +
            {MAX_SUM_WDTH_L{1'h0}};
          I10ad572ca72c2ea991487c39f7eabd7b <=
            Ia4b2db3d48f946b0bfd0be0e32d7518d +
            I111ac0aadbdd3e4479ca0786491a7b08 +
            I7caf8c7496dd96c1ed08e98b415f5775 +
            Iec0d7ea31e0f1a75b15121090dcf1e11 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie9f3fd3a6d16316e55addbe0e336519f <=
            Icc5d7bcbd7fcdb5092e6d8e18f6de6ec +
            I27951ef3d612004abdc639662807426b +
            I6c9ae8b8191507f908c27bbde53bf2d5 +
            Ia98bb3648ce3719b1c31ce0f41121c63 +
            {MAX_SUM_WDTH_L{1'h0}};
          I07965bca84276dd56da1af98e64b0adc <=
            I5e0d6b44474a226ab2ce916a6d46072a +
            I9068cca0de6ecff56ca542d0998fcab2 +
            I9cab38b69794ab661e12750cf69c822c +
            Id9c8055ef530f2cb8096cb7bb2af55a4 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ic2ade31b8bcf68c4dcc1a371ff14074b <=
            I5bab5ae46114c487f67b8e779d7461df +
            Ib3ec015a3d43d46e0b7142b21a81cfee +
            Iee0e45914c52a357e1e32922299d6937 +
            I1684820afb9d9cec38cfdfcd6ca8b36a +
            I25888aa2135fc403ca9eac4df634549a +
            Ib9081d438413a627f5b16f68c2eabb80 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ic0edcf240048fbfde4e938c3e4c5e281 <=
            I4d908bbe633c193cd9fc93dd33c60bd2 +
            I65928407b1d5447dbc815cd2d2e7b37d +
            Ic7855ca956651bd368cbdde7ec93ba6d +
            I7a6ab9e700bd94208ab6528af413f3a9 +
            I7fc6e2aecff5bd691872d1e10a39103b +
            I9c5bf5451736358f8c84e150004fa5a9 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8b42e89ff5f780d4ef8cd1cd5c99ef61 <=
            I83cec264bd378f1dc23f87e439e7310e +
            Ib83242b57ab050b0e5f9bdf91fa118fb +
            I8ab7efc436a0f2cc3efbc299a0ddf914 +
            I9b1390839ee2b9ba591e3873e967c8e2 +
            Iec936eeebd1f8c95307bd8705e6def81 +
            I377933518c3807edb71f648c65ad5c85 +
            {MAX_SUM_WDTH_L{1'h0}};
          I70b1b8521b36920707e95fc9418eb8a9 <=
            I0c53d8d6a5b92960e29fc31cf456c23b +
            Ice4f4ba8bb3381c8846941d5d5fe4534 +
            I2b0b168ce4fe8aa4a2e7cb69fe532aa3 +
            I2e14fb1e667e967ab4c116e0c7438aec +
            I24180fba17c21bacefa8a4514e4b685c +
            Icec98d794a64752081fadfa74308fad3 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4fb1c32a62cbbaeb585c6564a3c938f9 <=
            I45373bff54eccf8137da2931d841934e +
            I3934ed7170967ff3852944cc39ba1de9 +
            I17e818b67440efaba9a5d19e7467bf85 +
            Ia5b779ef95333736b08f63770900e275 +
            I83bbe6fa947f9f909e1a6785ab31901f +
            I7bbe4d0a7d61d3f7da346de71b9a3a5f +
            {MAX_SUM_WDTH_L{1'h0}};
          Iefc37daeec14e14ef2fe0716f73109dc <=
            Ib14733d3585dbf7f196cfc068e9508f0 +
            I3e8d26ea83937cae01aadf1092c59bdf +
            I0fb60c4f56f6d7b4007cf0dae39f4573 +
            If3bdbb4c20efca0c5af78614b4271ed1 +
            I632ffd09a9091335b3aa91ab2a8f1cce +
            I197c05f74bf7fb8d44124d40bd7c6563 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibd15f164f6d2ac9e5721a21464bc2c5c <=
            Ied7e494fb288f78d110ed06662f1926a +
            Iefe423653d454e21324a6857b52f98ac +
            Ice8a82bdd966719098a8d5f2a826f73d +
            I3a47540f34ce47bcfa1da66cc4e6e088 +
            I49321308413cb4dbe5e6c01ba5b9023c +
            I92acc55d81ec6e02880337b0a451ae21 +
            {MAX_SUM_WDTH_L{1'h0}};
          I951dfff9507bb70214d48e03a0ebb3a7 <=
            Ib16c6096ce80e2f15a5ccea145e28510 +
            Ic57a2627a194099105a2908a41feddfb +
            I4481555c402ba99bee05658ba6017984 +
            I9c68bfa3b888b6a6d41e38e674578284 +
            I6332af145d560e3f22a4a88106749f98 +
            I35c0ca76b28cd2f9355276b5d2f29ad4 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie78e30b2a2eda75d0df7d10fd67b5e36 <=
            I8cb171677016e4309034dc5d83981a48 +
            I4d1ba6ee8fb9505ba3b58b2b7553245b +
            Ib849494e5087777f646ee0947b4f634a +
            I283331db80e6d0891b13dc55e6a7d76c +
            I0c1e4d400520935c5c78b792a9d554ba +
            I29da0e5661f29bd8493c19885c998582 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia0b83a372dd4115dc4d61eb8ff0811b9 <=
            If5b3850da967f6f3d7a71d680341ad1c +
            Ic690477b1672dea4905a5e1c92b47366 +
            Ifa67d343acc6f3ec50c2b01fc26b4374 +
            Id27560fb44b4f2fda98d47e9f20d6898 +
            I0807a826e91f92ef279ccf0b6512a428 +
            I9426c8c1b4d988d5cd7d89a7aed4f8fc +
            {MAX_SUM_WDTH_L{1'h0}};
          If5c5bcbbea01aa22f242b913f0d01929 <=
            I7be8b2f8a9fe8e13001c2a1fce4a8a3f +
            I90a4190941651d885d04deb86a163365 +
            I24b4c998d19ae97f7178e37f75c77d06 +
            I0c121fa3e9e6e0e2e8291a594d6b4ceb +
            I4319fa23d59f4e690e31fb7e3a823d17 +
            Ibd010f15e36194cbd2ce9f01c98a2b6f +
            {MAX_SUM_WDTH_L{1'h0}};
          Iccba58cd3519fb4cc75a61b50da1d562 <=
            I223151b6414d9979d71023053dd3f5e2 +
            I6d6a242cdfadfc97fe656510bef73adc +
            I338400586daa58006c0a3dcd82ea8f4a +
            I202c385beeccee309104b66f8f096b2c +
            I05a812cd935867d1e417c64c26ea0952 +
            I7e86ab53e6d9647b230a94e076831ba2 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibc0999e4d0b3cc2650f9348b8c204b14 <=
            I0e7ca2d6470b9bfc6a1ca6143b468507 +
            I0aa5522190c741b7df4c4d7d34e46987 +
            Icf7630b6002db2f9b59d5323d6cc8105 +
            Ia0ecfaedbc1d546d484978fd50096d10 +
            {MAX_SUM_WDTH_L{1'h0}};
          I2aeff1fb4b839a581acaf26f90f9113c <=
            Ib9322ec1d3866ba3cb42e96b5ff5cfb2 +
            If4d030e5858f325debc6f37abf4a7d6c +
            Ic35d5ac4dac46d47b2796bbac6452161 +
            I27098cbe2d4fdd634385d771cc290c2b +
            {MAX_SUM_WDTH_L{1'h0}};
          I7d60d53f883f8187700c4e78b4c22f1c <=
            Idfcf7f3240d92bfc87d44833bc00ff9d +
            I73d2731c1b1ae5ef73ce0eb9c8995912 +
            Ia0caf6693d441ac622f416a86b665166 +
            I5d7a0739e447775e00115799c52b11dd +
            {MAX_SUM_WDTH_L{1'h0}};
          Id6fcf4b7af4a37c854a12e2ae80851fa <=
            Idd5b362dab4f93bba0c39af78c4c5981 +
            I2a4b3573ae7c3b38ec34591f20c1d076 +
            Ibb6e54edb9d277242c06d386a9a75a26 +
            Ie95793e09085b6de1383a37cc7fc41ac +
            {MAX_SUM_WDTH_L{1'h0}};
          Ifa5e5f7d753964f14f0f16dbe552fd85 <=
            I627e4bdc8061c69e3fcac17535b9f1e0 +
            I28ea268c5b51ac1d9249e96599bb6b0d +
            Ib97b2670a6cd88b2327f07f62d887900 +
            I134a734d93e62f6ac6635015fe3a2096 +
            Ib24b68cb35da39a743e1d90bba3f0836 +
            {MAX_SUM_WDTH_L{1'h0}};
          I900d471b087cf5a436c2ad66a84d8280 <=
            I5ca15c7da1f49580ddedd9ff8ba822c0 +
            I6aba8ca0e4b20a6355b43a70f19d9d8c +
            Ie9a316de516ec4fb828a614c67e38b2a +
            I745187336b8a5ae4eac66e90539752cf +
            Id4cdd72193e90dddd211af73d7f3634a +
            {MAX_SUM_WDTH_L{1'h0}};
          I6d1434907f0292ea2ee47cbc5b52bfb9 <=
            I276c2ce5d3a1b7551c2790971071b094 +
            I77fd8001d879fc9e9117464fba27902d +
            I6d0d098e6d47dea04d6d7be67b648a0d +
            Ic3c59a5167cb83fd76ec6236572b1f3d +
            Iccab4c19a9190689f90a42160e2379de +
            {MAX_SUM_WDTH_L{1'h0}};
          I938bef7ba7ae1739d8e6a6a7c117a1b1 <=
            Iff777b2c4a3939e330c4cbb36cbe1ac5 +
            Iedf37dac8b3a5331277ae4f0176968aa +
            I3f6fad8bb0fba790fcdb1612b6fa7712 +
            Idc549661d6694035874a3366704801c7 +
            I275ea08a3dc0600d8ccb6300eb7f2a6b +
            {MAX_SUM_WDTH_L{1'h0}};
          I6384a9416b2d1da01df1b2d7b16c5390 <=
            I0a9cb91319cc0d0c1c4d0020cce321d7 +
            I9dff504e40aaddefedbb7b0f822c844a +
            Id9edc6ac95a260bf5af3de25f00e9e9c +
            If0676ef300628c4097565b13ef2d8854 +
            I1b53098a7240d2b5dc1f5c5c3b4bcc11 +
            {MAX_SUM_WDTH_L{1'h0}};
          I5097a79e7cf7a30d38ba198d1407119c <=
            I1cff7306aaf303bb3342ea3d72048908 +
            I2d839c10960739097d449efab58b9fd4 +
            I080832c25509f7003ed50d71210bc7f7 +
            Idb73eba1bd4ce25a6109e296f51e7dc4 +
            I278659ca1a0b093fc883d01987989dc0 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib113c26c8dcf49c972c41a938059a787 <=
            Id033e7adfcfb0420cc592a1fb6c297b6 +
            Ia443284a35e0873de59b3ae55b7f809d +
            I2b807c16cfc6d65cb2a7f28ffa837974 +
            Ie467c5fde1d123da4e9587b5a56748a0 +
            If92e66cba66732798dd19f968a5ef8ce +
            {MAX_SUM_WDTH_L{1'h0}};
          I970c4a25a8bce82a9d2846679029fcab <=
            I4ba05e74c2f63e2f4c59268775d549aa +
            I8289bfc08a5d8979ec26825bcb6e3d18 +
            I2b32537c9178028493af165398a60875 +
            I18d0dd7a10d6533f721a2392d4ad2d02 +
            I784c4e9fb75c314f271477e0621aaf7c +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibe2af096ad2db26e54d8b4b3bb05175c <=
            I299b37fd45c6ee2031fb2c74caac73be +
            Ib8603cb82ceb97c2f35bf8209306a457 +
            I18916d0023ca275d84c52af07dcc5ca2 +
            Ic7d5fe6c4b1dcb97d10ba3de2f95d1df +
            I3d3aafdd4d9d3e9fdab1f487c48a0ea9 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie48569c467fba0c1291f71d6080ebedc <=
            I26bdcc44692db066911c8d5b0a1aae0c +
            I8d26e73fafa909f1e26e329828cf4888 +
            I2c72d6c5fa6968dffa6517cf81219875 +
            I05aabdf73200996b7bea8db700fa8930 +
            Idb4c722992139f39914af7085378c6cc +
            {MAX_SUM_WDTH_L{1'h0}};
          I90e7ded06617b49cdb8b5301fe9c6a20 <=
            Iaee91a5e94c3f174682f72a1ebfd0021 +
            Ibc1a16427d8dfa5ee20dac15327a53ea +
            Ic1120eb027841908cd64fe5c7274da14 +
            I4ee3f608cc8f8df27345949f1a3713a7 +
            I63c9deb7e6a4b400e0aff6887a09e647 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4920014f5d017f4e840dc3b88526955f <=
            Iaed26e1c4a2578d16b111d15d31339d2 +
            Ifc52604a4f9f9de392a35f2f9fe885b8 +
            I4037f1b207aa101f354e59eddd7c9eb4 +
            Ic0a580f94f3d03f72e3a487f84bf6612 +
            Ie6f67c6e4c5e2b8357c0a902979e8722 +
            {MAX_SUM_WDTH_L{1'h0}};
          I03b70553f1c501609400574ae7cd73f5 <=
            Ibafedcf9f2990ed9c1efa973a0b1d81d +
            Icf4405d4a4063448a2be8ad0354ab1a8 +
            I778fbaea65beeb6de599490daf3b7e3c +
            I1d7a4f99e3975fd01bfe5a9a1da84765 +
            {MAX_SUM_WDTH_L{1'h0}};
          I63c9bf68b43ed66c51b0f4c0ed92e9ab <=
            Ie3c88bc240576aa220f0f110b13bfdd3 +
            Ibc8679379ddc43ee4bc508a1f577eb2c +
            Id66798f8ea67e74a67f264fe6b4503a3 +
            I059d847e09f5aa3f6a8147062f4b13bf +
            {MAX_SUM_WDTH_L{1'h0}};
          If408dfead07757878cc878131bc7d6a3 <=
            I4ed5da534afbfe9ecbc10ef4cc649a55 +
            Ie2e3d64640c339dc51512979dbd6a173 +
            I772e844c41387e7079259875e0ba3fa0 +
            I48e5256ade4d061a3b5ba08a53252bc3 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia0857d63d309807789b6ff4f6028f1b3 <=
            Ice8765807beffd3acf59fa137ee0baac +
            I6e4786234b286b12c83e06e93c628534 +
            I3e8e280553edaa5c8555ace81ecc10e0 +
            I635fb29c55e0fb5cff0b6f443c2e3de5 +
            {MAX_SUM_WDTH_L{1'h0}};
          I53921b825c5e434b63bee0e1ecb7a517 <=
            Ic2f450f7ab60ba57dfc1406c92c0f077 +
            I529eaa7e5eeb6d0a1aba78df5d5a2fa0 +
            I839895c8614ff28df83314c44824900b +
            Iede5d56e52612e083407888da49470e5 +
            I088c5b971a2def57248769a33b7d2a2d +
            {MAX_SUM_WDTH_L{1'h0}};
          I5e68f84e123c37f19a03c13892c77e19 <=
            Id144785da9b171f1e2d0e9182d693e31 +
            I439c7c302b535bfd7db655c3c607d71f +
            I2a0dc4ed573a544cb13544e049514903 +
            I39d9044227c161f0163e58dd82aadc90 +
            Ide22394fce1658f9e7002bdb30d03c2f +
            {MAX_SUM_WDTH_L{1'h0}};
          Id5270b57c6fb4b18db3bbd0a523e467e <=
            I0cd8a6e719305ee3fbe8228081993957 +
            I583c6d23506c7d7b84403bfe977ec1ec +
            Ia422fbdf8f318ff3ddc049d1374e7939 +
            I8efad9622c05177563ab8a2747879044 +
            I9ff276a14d3205b98174a8a736f79774 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3c18a84617eb21472d53e598700d7f4c <=
            Ic566fe27ccaf2220101cbc49fc187a6b +
            I618363a8ac413dd0ee52eb658940eaed +
            I1d648ed8f07f0743a6d616584270c513 +
            I03038b940be8bd21bd26b150b28754a6 +
            I123255637493b9c7924e3a72d1b86ee9 +
            {MAX_SUM_WDTH_L{1'h0}};
          Id36663e7a01fff3170833ecfecac1321 <=
            I2133d362ba45ceb3dceaa84e95ace1e6 +
            Ib43383830037df764b48c637a28ab6b5 +
            If2ce7b8d2573494564393f7d426fa47f +
            Ied4ddedaf801fbd7238d8a55c17c8090 +
            I87e6ef84894cfc86b94e19c9d3065bc6 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8d3be15109c7007a79fecaac0d891626 <=
            I768afe193d9d79b136736abc6846d945 +
            I0aa93075086164fdbab3814d60633141 +
            I32c35da92922c5b477f8aba837fa6d92 +
            Ibf547f8a5e1059ffaabeb3f447904dcf +
            I4c32900878260a261bc5403e8abd6258 +
            {MAX_SUM_WDTH_L{1'h0}};
          I92169cc57291f20d336a479e392ec271 <=
            I54166b387c02e12374d6febc425bfb7a +
            If06a1563b9d7348de03a98d31bd85b06 +
            I3e466d40a4447a23953d96d2e6d61d47 +
            I3b2739319710681986b9d3f8cd04f619 +
            Ifc100357ae3f754fb0e3863334bcc764 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6178b220b469b40dac39168057023a1c <=
            Icb2805685607d5fedd0300c9d800f863 +
            I28fa295ebd90c2b7255d48ca9ffcfcf3 +
            I4fd45670f88265e5d7aa6582f3ad3ff8 +
            I5f607bdc9b276fdf07a17a11a20a6720 +
            Iefe9e5376010997c0ee52eeb28e57a25 +
            {MAX_SUM_WDTH_L{1'h0}};
          I55342938216a0ea0889f96c2f6c05ce5 <=
            Ieca5b21b91e150c9d509964bdcea500d +
            Icaeb9a2ec8ec5822658fa85b88cca04b +
            I76e4c55148effeba62a4837cd19c5e51 +
            Ie6060acdcb16b6fa6aeeb649ed621053 +
            {MAX_SUM_WDTH_L{1'h0}};
          Idf28431c76a84a48dd895979d2b11a63 <=
            I6b7a8ba12de5b44817ec99faebe54617 +
            I58416287b268462d28f55c6c2705e613 +
            I2d636a246d815a4d12c478794860dd40 +
            I46c2b923860b0d1c01b9475f4467f280 +
            {MAX_SUM_WDTH_L{1'h0}};
          I1ef61124c8d62e8f6a82a729fb091694 <=
            I9b8cfdb69b76453a3ac687a1e098417f +
            Ib2963b82260024e1853d297798d88d3c +
            Id59cf860d9f4aff11b205b8970d93df3 +
            I38b4eceb159ecb0dda3920290a21a02a +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib8bb96f0372323e6a8072ca56fb9396d <=
            Ibf9f6d7baed9e761b69fb41442761ac6 +
            Ie945349d77442536992d9ad52ce84218 +
            I3bc01b072987a0c980615abbc2251e5f +
            Ic45561ffe1837c3d5bb42c695a377f82 +
            {MAX_SUM_WDTH_L{1'h0}};
          I432f74dda4f6b1cebdf5ad59c659080b <=
            I67534b68fee8f76ac0c5e64cd02aba42 +
            Ic79072d9e42dbc9974231f1d642b3f12 +
            If08adda7d796da7c7849e472a73282a3 +
            I3db0adb3457cb22c755f5d29a8fe7ed8 +
            I3e76abc721bf7ed186f4d0f8f4bbf4e3 +
            {MAX_SUM_WDTH_L{1'h0}};
          Idc689442305acd00f0f32416d8fb3773 <=
            I277d7065150714e33d8ba64875d18190 +
            I9bb4d58b1fe80549451b00c4ed2b3885 +
            Ie335e68643fd2b0a53351f4bd45c3475 +
            I32679702c19eab37b46d13bb372967ea +
            I1afb4061458e9d2f5799afa1f2373bd2 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ida03738adc101c03c2229756bed2469d <=
            I0b6cdfa1dbfa774fc9a12d856e61cddb +
            I5160de2c5ce4782d8f8be10dc740694b +
            I3319313fe1d2b4ec2626711b187b4a5a +
            I85dd6a9634284c22027b4241551ea628 +
            I18bb9a781a4c314fe6bd990e4c275f67 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4d14c75f28f3e516c259ea288996131b <=
            Idadf072247b351cf51d718f797c3b375 +
            If4d63635a5f99c4dc9e5b57712830c20 +
            I75aaeab4f372e28a8e51453540f9c6b2 +
            I51b1cd475d0e389326b182cbe680a402 +
            I49d7342f105c4502377abd23db973752 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6e6cbbf430d57f347a0d70558af143d8 <=
            I6fcb3b133a6a654b69f41468a713d922 +
            I5eaa11e26f19b94dcb7eaee7f09d24b4 +
            I586aaa5c55efd37996b01febd3bc60a4 +
            Id5cedaa397ebfc2567efcc2f8a648db5 +
            Ieeb12d463444ca36af1ecf2e09504c06 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib7487df45118e44acec6b9d07bbd5969 <=
            I8613cac4ccd4f956e8a0ae7b627f5be2 +
            I7d85b73e85379bf3a480e954c05516f3 +
            I2266afbacf1ba750ce18f296aba1181d +
            If12366160fdc899bd71cb0de5bcfd84d +
            I17525df1798fa2c1c4bbc4a1ddcdd0a5 +
            {MAX_SUM_WDTH_L{1'h0}};
          I492f382fea500462b3d0866240fb91b2 <=
            Ia5c77c9be26d62b026f24ee5a5e25fb8 +
            Ib5c8d91204a2d313c9c23110a53cd0cf +
            Ife3bb8945e14d8746c82b66886293997 +
            I887911fd9466f4d4fa7f50642d610d88 +
            I90c44c31fa7903a81826c1c568597362 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3fb3ebddaf28efb56092d19a1b4695de <=
            Ic4af6c9097257c9b22a57ce4b79b40fe +
            Ieb7b388ff89e352dd239e0ccbe7b9ecc +
            I89f75107ea95f207b9e664a1f4f0746a +
            I6a86b03402bd2e35208d3fc74601f9cf +
            I3997cf122743b612f49cd5dd125a9201 +
            {MAX_SUM_WDTH_L{1'h0}};
          I22a26b7f0b1c8c16b00597732ce2ab23 <=
            I4a403449a9ba75243369032e1cca1a0d +
            I886750aaf8d2040c3f12ff113294f658 +
            I0e52c25aa840402d944cbd81f73c1ffe +
            I1112c4267582ddb8148ee40d9529beee +
            {MAX_SUM_WDTH_L{1'h0}};
          I2ac08a2d8c917ecb37fbaf5325cb0473 <=
            Ic2159627df2efa5e677fa6f4498bdd31 +
            I58a7c7b05b84d292cd06d68e96ecb9f8 +
            I20c4e393929b875521e5316f4d8e2d42 +
            I21c207af859b94634d3750482b42a2ca +
            {MAX_SUM_WDTH_L{1'h0}};
          I50ff8f51e75fb9ce3db983c2a0f57196 <=
            Id5b4ee69444e5b499476c05a7f1d6e60 +
            Ia308e09137af1cb50167562efb5da628 +
            I2418ae211f327ed45cc70c42078180dc +
            I2ff2421bd86bf9ec110724460f1171e9 +
            {MAX_SUM_WDTH_L{1'h0}};
          I444bc340ffb7ef7b72d4d2e761d58872 <=
            I48b39ee498563e23c3a4be079b6100d8 +
            Iddf65ccb4396288264a400ba37cbb655 +
            If29fcea810adbdb1c4d8a4ace1d8081b +
            I6ba5c453b17e4b33c61caf5d70041c4a +
            {MAX_SUM_WDTH_L{1'h0}};
          I039c6cac5830759529595a958b7f65c9 <=
            Iac8cb32c2d86b975f51a2ed605002e51 +
            I88a325547ccfe4eabf90792abd60e356 +
            I0722ec4e9d400f8eaeacd060e42de79c +
            I08318099725fbe033ab8d5427eb8b278 +
            {MAX_SUM_WDTH_L{1'h0}};
          I0584de7d919236ab138e288a27d08ff1 <=
            If85d9a95c1c02ce2da1dc3486b53eb81 +
            Iae21bdea20a6266d3f69aa680b6b2817 +
            Ic6a7a82d16e6106071934ba79d3698cd +
            If36cb462cdf20b0b1758cd6417e524fa +
            {MAX_SUM_WDTH_L{1'h0}};
          I086402c82ec67ae09a9e6360c58904b4 <=
            I59fba74472ded0a985cb237104ac127f +
            I77e1f5f504a794edbb89c66cf1ffcf66 +
            I3cc30aaba3dcd3eda262a19e85e53117 +
            I40e8463645b1122b7cb224770fa00447 +
            {MAX_SUM_WDTH_L{1'h0}};
          I1cefdc831c146187c77f861b3e2d1af0 <=
            Id6105518ade80c89d4f20222a2382efb +
            I8493e2dac01f009db1d2d5504b49d135 +
            I106d0e71b7378d110b0a624e5cbf0d6e +
            Ide386e751e06dd5df0c042cd76f0f800 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ida9c16ae57d17b6faee8a54838860447 <=
            I185085cbf8da6df921ba32442b28bcca +
            Iaf3a0b5ea5d9eda47fcced9260922bc6 +
            Ic8f0049e1298b14b4e039075dc0d5f74 +
            If63bb4681bf1116c0d1db3aa21bf52ac +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia3b9fb112f39dd0ccbf7555659369efb <=
            I5c278aad08b7c4b0237d68f88fcb3f3a +
            I9222c4c0eb2b110fd80547d46ba17036 +
            I95ccc219b5f5038641b38dff6db0b222 +
            I566c72342c69969892480fae41232c37 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib1bfcdc0c972aafc99116ed8c0511445 <=
            I21842d06e25948ef461d1fd03485f86c +
            Ib2c1636a66f6479d6123a038cbc668d5 +
            I69c2b063e61e14f5d49b907095ece00f +
            Ia0f7deea6b1ce1050dcf97fa99de9178 +
            {MAX_SUM_WDTH_L{1'h0}};
          I7adff505c50450a04f1717cac1adebe7 <=
            I37e360420c7dd061de93a6647513676d +
            I535b29f7177b4fc009ee998f1f4f7d7f +
            I45ef0ac486fe043f57e8a46aa91461a3 +
            I992b9876530d53c1b62d98511bf41942 +
            {MAX_SUM_WDTH_L{1'h0}};
          I699feb4382974a02b21cb387c13f7f3f <=
            I8e470b68bf35c647af42b6e46201e570 +
            I8cbafa797ef136d7e50c909dc160deb1 +
            I850c257a0412bd9bd6001817bd9d0ee1 +
            Ib8861f627f6273c0a031bf43e7812a5d +
            {MAX_SUM_WDTH_L{1'h0}};
          Idc99c3b23e49aca3c98f0685ea34441c <=
            Ia526539cc0f844b802d412b7a17cb6a6 +
            I71bc7271cc432bb3c5d0b7a416cdfc60 +
            I12e8b8cf609c2fbdc72efce9bb5dabee +
            Ieb5bac4ef0f5e4e0b826cdc43ae71471 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib67318fa6954ec8f3247927d34e74f8c <=
            I26cf25e680483bf4e556d74efec35ee7 +
            I9cbe73d708c561d43d05945552d32dde +
            Ieb9720b6beb2363d651346ef0233cd49 +
            I3cd0883d9f0ba7475f474f1e318ef023 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8774ce3f11362915c4331d1026e452dd <=
            Ic989dc794ce4356856b3916ab1889589 +
            I82a225237aeb1ceb31e8cd18b1e45c6f +
            I2ea27544ba4cc14d0f7ccf7158a27a2f +
            I5f8a41ab83a9257e534973e981e28e9b +
            {MAX_SUM_WDTH_L{1'h0}};
          I2392b2d17ffed6073875fbe8e92534cf <=
            Ibcb80df5bed66f8498561e3f3ffa4ec4 +
            Ib7fde6a2ec1ff0a3af10bccf3012e63f +
            I0e420136675d5f0d1aa027d589ee8741 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3a4f0d3e32596ef05477f494768d4266 <=
            Iba75ff0f3b67c7e28cf627706733d528 +
            I4854ff71aa885da3d07acaaa24740d7c +
            I4aab6ff52e3fba90bb7417cb50766125 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icd08ff59cf6be3ba97698dd55703339e <=
            Id65f22fa8fc9c47bfd00c796b63c9fa4 +
            If7543e2f5a158b1f3f3a4078ec54cab5 +
            I1ba7f209cb735471073e8051026a148c +
            {MAX_SUM_WDTH_L{1'h0}};
          I985fb7ed22a8476ea322c9e3c2b3851c <=
            Ia81c31ea4f4786136b539c9766987596 +
            I6a3824a6598bbaa138e1e763ad85f5f7 +
            I711c5cf9fd8c5161bac36060b3443503 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ib985709316b1b0a9d3fa3c1eaf6c641f <=
            Ie380b37a78242e6d45b659d568887457 +
            I72108531a608f6d5e51a481c68d7b271 +
            Ic9740baafb1c92e3a25f0a1e7bc46486 +
            Ie3591b22e0e127f04658da68d4846be9 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4be898887dff6e2cebe53f135ece131b <=
            I484ec87270fcc959a486ebce40a9a03c +
            Ibdd9957b7f1a319b797c021933ff75d7 +
            Ib1461f456ebc14f449eee77e386a4c69 +
            I409129c0bf5d361e9916b6dc98e69a7d +
            {MAX_SUM_WDTH_L{1'h0}};
          I004db04f61fb57aba81e15cc015442b3 <=
            I5d80b7c7d102d2c2bfa73a68c73376be +
            Ib2c327648cce481482eaf0467e9227d4 +
            Iaf1d3be13e6441a7a9ab3f286a7dc21b +
            Ie4f4faa470f572da2081b63b6df6e392 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8f7e3dfb2f728d4cd1e79b82b62b0406 <=
            I8636f5c91b567780d3324e4b8a320fc2 +
            Idcc745602c4b7b34df9c3d68f9a9d76d +
            Id5c9a9b9c34c8f9d56df0aa8d780c9d3 +
            I5011dfbbb0eccfebcff255e4a2c5e64c +
            {MAX_SUM_WDTH_L{1'h0}};
          I991054370345e61638ddaf81785505bd <=
            I2cf5304a672431888916e08b3c15f0c7 +
            I989091b3586964ab598f166a89279d16 +
            I5f7b6e6a30348ae86057f7e56f625846 +
            Ie32ca6b91d1c55883be8f63acca78764 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ifa1f503965270d10e7a5c9a15576069b <=
            I9164fa2a9a33da6612ea692cf3fa7d2f +
            Ie8befb003fe83e774e8d1d01d4e2f4ad +
            I1f1f2fefd3381ee48ab0ec9c9301754b +
            I6c7965d39dc839a9df56e628c77a5457 +
            {MAX_SUM_WDTH_L{1'h0}};
          I24f773842a4742fb58d09cae45717b2f <=
            I288ff69a7395e74f7de8da5a6a7f9062 +
            I98a2aa729628adde0b6047869bd12743 +
            I1140fa91b5e22ba0c094c03295781e5a +
            Ieac9cea5f36bd82f87105b530e8fb614 +
            {MAX_SUM_WDTH_L{1'h0}};
          I5bac7e0d778a547a0ae764fe259b6f7a <=
            I5a4f0749acdc34fd0786e4b3d062f88b +
            I283107989a436e2c720123b8d9e335c2 +
            Ic488e78b5c73251b673301e84c4b5b0b +
            I79657595561eac53237215fb4110f09d +
            {MAX_SUM_WDTH_L{1'h0}};
          I255577ebee6768871df0224fc1db2db3 <=
            I079932780612fbce79cbe9b58bb6c2b5 +
            I61f5ebea2bbe443b644c95ee559c2234 +
            I9b46463a6c54c3668e76190d942b7b38 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia7fb4af3d3529a32f902a52cf5598474 <=
            Ia92defa0ca87c7c30fbe901da40a575e +
            I21255a0ad20a9668c958faf68d53b2bc +
            I3ff883ad434cd5153b67186b6b21418d +
            {MAX_SUM_WDTH_L{1'h0}};
          I2c98806141f064c9e92935b23a84ede1 <=
            I914bef0326cf82d350344317eb1359be +
            I6f69796a6fe6da57066319ec8210c1a3 +
            I92abaae6fb89206885616877cca1e25a +
            {MAX_SUM_WDTH_L{1'h0}};
          I5680847bc8d224fa4ed93b2fc0d841e1 <=
            Ie43a7f8082f91c2955076a6373028b55 +
            I8786eb767f02164cdc32f14f41b5d0e1 +
            I33668b0ef7defef974b7a4c0f87689c0 +
            {MAX_SUM_WDTH_L{1'h0}};
          I365254279ebb10dd7ba0b3482d5e34cd <=
            Ibfb57f2b507c27759a3556759f23977b +
            I064499f0315fbeec7b6cb50583388a07 +
            Ica0a119af1728ae253c16cc3eb93f802 +
            Ib7875bf9d30d071e62a474c50d88ba06 +
            I338daeacf82ad288b14c6b5bd4099870 +
            {MAX_SUM_WDTH_L{1'h0}};
          I57bf4ad773cc058ae1bb7b1911dc3174 <=
            I7b12345fe53174cadef6811fb8869b42 +
            I6521c9167261db6eb37f50b66159ddb7 +
            I44e5ce0cdf812c5b73e6e638da36e414 +
            I6fdccefd034e8b4b86cfa997502512ae +
            Ibe085a39ecb07a8dca62002afa38df93 +
            {MAX_SUM_WDTH_L{1'h0}};
          I57072dfb29c4a3d2e2b40e46e62f0d95 <=
            I9785922874bba479ce4a9bf1759e2933 +
            I0e3286fca6cd040758950259ab663df7 +
            I9ae284c0089ae462a1bb9d168bde2fd0 +
            I202aa0814e7e28a6bd21db116b652b4d +
            I1f88dddf05f255942e2749891a7733da +
            {MAX_SUM_WDTH_L{1'h0}};
          Id8cafb6f76321bdaba9711133be7be99 <=
            Ie7e196fbb66ba6bee51ef0064ca519c2 +
            Id7619819e1297844d92c8bf3a1d61926 +
            If8a259e0c4f1839e852abec6e1b904ee +
            Ib2f34922b0d5346500de093275bebc94 +
            If1d0be4e9b995ec98c346e8392b9518a +
            {MAX_SUM_WDTH_L{1'h0}};
          I6344e71ca2b0fd39d36caedd889c3085 <=
            Ibb157b97546cb19fa7c1c0a7c79b1d38 +
            I3fdec80112b3fc543b217d1c253406da +
            I56a4443759b3d786bc9a34a0dc32abf0 +
            {MAX_SUM_WDTH_L{1'h0}};
          I0c99a68e0bed90afce18807acf7d55bb <=
            I8fb1602dcdcd2912ea8aec42e2b7848f +
            I5aa85d9503b0e4ff46bbd63e873053ca +
            Ic826d371f2cfc503f5d9e43dc17481e1 +
            {MAX_SUM_WDTH_L{1'h0}};
          I1c95650979c86310ae2a949961c9db11 <=
            I7de222bc26e38b8b6543819701740302 +
            Ia7673d73f0535906a99d6cb467892104 +
            I5502f383dff392ef1be4cbbf9dbc3c2f +
            {MAX_SUM_WDTH_L{1'h0}};
          I04eaefa5d133e53494fc270b07be7043 <=
            Iea765ae5e9c65b3186445b15c56f69e5 +
            I103ec7cf279f527fc6e3648a19a12a8a +
            I96e6f1dc0cd451da6ac9170d5f83976d +
            {MAX_SUM_WDTH_L{1'h0}};
          I4a64fa2412eb8058c2dfd9351d7b297d <=
            Icf266f710358631b7119ef526acb301c +
            Ib20dec1346f227042c749ec1abfa4d39 +
            Id6fa8ec5d1062fc3e09bdac65ff79f45 +
            I10cd840a369d3e25556a41beede2be27 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie8bb2fcb752c6a33254963d1ebb4130d <=
            I0f3c4fb63ef1e88168b4d28175a0b68c +
            Iac6fcccf3a0cfe04edc0d998b60c2681 +
            I1fbcaf2f6be01b129ebc24dee8a65396 +
            Id85c2285fcc45211f0fa6963b74a663a +
            {MAX_SUM_WDTH_L{1'h0}};
          Iac05b7e3ae18f948b72c356ccfb8000f <=
            I2ba94ef71f97b9ba731b306d4a5fd02c +
            Ifbaae8b3da03911a4c96d4efdb9283c5 +
            Ifba1584d599da13b98a3b76b4db10974 +
            Ie0bdfac78159144aa65090028931a3bf +
            {MAX_SUM_WDTH_L{1'h0}};
          I27da3f75cca6c49e55db90306aa68e94 <=
            I5529d6db17b6184c45cc4487e5a2c24a +
            I685699f60c76b00df87c9c53e9a8e448 +
            Idb862697f62a6c678072de760e176096 +
            I28fa30cd1f3b476fa6a354863108cbcf +
            {MAX_SUM_WDTH_L{1'h0}};
          Idc7fed723190098341225fe01ba65ced <=
            Ie3361a270ebc41698ef4651bb3548a49 +
            Id0842da8068ee88d99af7acea50e7b77 +
            I7a927f4f266cc5253ec30f5c127bb17a +
            {MAX_SUM_WDTH_L{1'h0}};
          Ife9065805598960919ee4f14c3cc6fd4 <=
            I74b55d2f94073ba8f948e4b02386867c +
            I03a8a458ee0942c35001cbfe8e589222 +
            I7571c7c306861230de71a75fca79c5dc +
            {MAX_SUM_WDTH_L{1'h0}};
          I717c5c2d6a2be61593492ae5f17a112f <=
            I45cb51c25c426c296f97a5d23a08c063 +
            Ic1af7410a9d11c5324f3ee5b2e0e9dac +
            Ic79811a48840357d0b6303e7b19413dc +
            {MAX_SUM_WDTH_L{1'h0}};
          I4c31fa8e6eb648439cdae1de1afe0d6f <=
            I0cedca0e2c589104d6f3318505910594 +
            Ica02d19b129c8b1d491ea4747a55113e +
            I0f29300446f020dd23cf847d3e3d3530 +
            {MAX_SUM_WDTH_L{1'h0}};
          Iead549a9af27f1fced7d9c36e7b5c3f5 <=
            I77a54091bc2c3d9006ecb3471b94d8c8 +
            I1c0df8c2c64b688ae417a238263f33db +
            I696db0b98e27dcc4657dc7feb23a881b +
            I9de41d0b279b84366640880dbd18c502 +
            I802bd5b13c183c37e842f7e9278f35a9 +
            {MAX_SUM_WDTH_L{1'h0}};
          I10422eb79364e7d0e21e1643d9060331 <=
            Ib6c0e635e659f54724737f0cffd1b0fc +
            Iad0f4602ec545dc6ef12aa34add00ed3 +
            Idfa432a87877e1ce103e56891745b62a +
            Iba52b84e6e215842e0ca8e72c42ebce7 +
            I0297905b35f06697625420b7fc2434f7 +
            {MAX_SUM_WDTH_L{1'h0}};
          I914cb87eba8baa40cd515334e59f26b2 <=
            Ifba318d4faf308168c5eac8fe92395b4 +
            I06e05a1ed002175a75d02b8b76f52c50 +
            I894ef04bfa1b7b39ef51b7c82f7686eb +
            Id2989aaee3930698cd374e6c9feedf82 +
            I8487a819dcb61016798cde56f9662fcf +
            {MAX_SUM_WDTH_L{1'h0}};
          I32ed679af4ab759901aee43c9d93eb67 <=
            Ic9678deca4bf44a7b99f853334f6a05c +
            I83b77ad1a40dc102f28153f692516eb4 +
            I920f95bb52cdc9b07f93afc3a6b5c009 +
            I8d07beccef519ab4ce4024d911ac2346 +
            Ia2904a5d5db43a209bd4b358ace68c6a +
            {MAX_SUM_WDTH_L{1'h0}};
          Id376dfa5141402f4d41a8858180ed87e <=
            Ia209e5b03deaf4fcb8ae12b731a49e0a +
            Id2e223005a932987b6f60663773187f8 +
            Ia8b29ca047a643f47bd3a0ffb50bf8cb +
            {MAX_SUM_WDTH_L{1'h0}};
          I98a384bc62ee03f5ad7df20ef2d9af95 <=
            I99d236d41be79090ca7ba1fb6faaec4c +
            Ia92b76ee5b7d82a992a1b58147c0c0be +
            Ic45d0537b94bc30713c0a0ee07b1ec40 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icfed259ca2bb2732d8e0c26ef67cd4cf <=
            I26ae9e570a101c6f8237d7941285b924 +
            Idcd5283cf7b42d403ee0e4404b5b311b +
            I337231f0dc7eb85f7d950262e0adb724 +
            {MAX_SUM_WDTH_L{1'h0}};
          I20861535c450d6e6bf11c45dac120454 <=
            Iabe5aea929c668c9b9728d073ffb00c8 +
            Id201f81bbd80a70006a10866b8efeeff +
            I530cf1f747d1df44b913f49eee90c079 +
            {MAX_SUM_WDTH_L{1'h0}};
          I013929385ad819ddfcfcc59c22902ee3 <=
            I1240c9410b897a4d0504affca5ba139e +
            I4f169c2c8c0768f2725ed655a03acfc2 +
            I342a563de39175fe4a6eb7e3e1ccac9a +
            Ief52461e4a5ddb128be5e439edf34862 +
            {MAX_SUM_WDTH_L{1'h0}};
          I34fffcb07fe82f11fe142f7c37f39155 <=
            I015630502f5cb4eb27b2a673e810f1dc +
            I8bb46c3eb9f54c5d1b28dc6aa0154358 +
            I938dd59e4cdf3434086f60d000113430 +
            I46d86bfa6de26f3cfef9d802549ef2ad +
            {MAX_SUM_WDTH_L{1'h0}};
          I61ca60fde05ed88cce714dcd8c13b827 <=
            Iff1d4b06901796098f91e87a3c30f7a5 +
            I1e110e27162231650875dd1152d96e64 +
            Ie7274a7ffa053ced4f12a67986d3c81b +
            If6a3bd6f002d91e0773c4ab9caaaa01e +
            {MAX_SUM_WDTH_L{1'h0}};
          I4907dd45c158dc7e0041c64f1fb388f6 <=
            I54c260db5c1b2c76527c8fc1cee229fe +
            I55e54359961ef6e5a63f1c2eb0ad4aa1 +
            I4f38c3d620b72f21cf6d54c7df4ba816 +
            Ib33e1c6d57e5e6fc465dc9c9a7cf29fa +
            {MAX_SUM_WDTH_L{1'h0}};
          I2c8f6a9b9f655b317bb0af4d60fdbc4b <=
            I3a8bcfdab631a268d21c87b98e9d1c49 +
            Iad0ecc5208263d239e4a62c5563f52ab +
            Ic0b2f9717b8aacb34325fd5aaf03a366 +
            Id92a319da408be46970faf524513fdd8 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ic7dff631559304ec59f0696c66436d62 <=
            I95b923444062b4a98918c685c65996d0 +
            I06c0921675f464807a63c7965796f0d0 +
            I59adad4fd84c1fc233dc58f70a12779d +
            Iae182ffae6cea89363f0ccc8b5679561 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6a239d3e55b4a9a3be9989a85bbec545 <=
            Ie40c90fdb38b3e4046ba89295ed77d7c +
            I13b9e098622d90a1074f636d8f351aca +
            I1972375d51767f0cffa5395a354b3493 +
            Idfe6aecb694385ce8c3c1544a4992a20 +
            {MAX_SUM_WDTH_L{1'h0}};
          I630f905e55f08e7d1569a08e937ad216 <=
            I9859b94cda465ceaaa5674eb19e94824 +
            I8d6927b0bcbbb318cf52987c121a07b5 +
            Ide40b1bf9c0b642c49a5685a62af1c93 +
            Idfbc5726963cfa31bb4324143ffd08c7 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8d13eb3669785c4279c685763d4f3fad <=
            I5085f161323433d8d38be2e4511b0c46 +
            Ib66b897398ea0702b74bdd03774f3ae4 +
            Ic227f42a20219c6638ee3343ca445acf +
            I205d5fdeae55fae7be2f06f11c949244 +
            {MAX_SUM_WDTH_L{1'h0}};
          I25a6f3de9a9a01cbbdd32ed848561aa4 <=
            I16db9cab1981451a02dab21e2ca221b4 +
            Idc758f8e6fabb6b31b0a7d9c0c590310 +
            I3188d354c2ba494ffe210dcd89c00620 +
            Ie667e1755ae1561a2eefae9b63845dec +
            {MAX_SUM_WDTH_L{1'h0}};
          Iba3dd4b2c2c85c4cfe770d9b52ef4634 <=
            I3d700e050cb7f22b0e381f3c72a20124 +
            Idc198bd5732ca5760d1a700a25273ce3 +
            I2253b32e46200a23dba243819fce02f0 +
            If7348fdbe0400aab92e8fd6a7cf6c267 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie1b744387b5200a504e4874e14d2f282 <=
            If17b4f86674bc5fb212a1f7751fb043a +
            Ife7985db888089ea618413810611bfca +
            Ia020344403aad35e050765a4b0cc42b7 +
            I143b91852fddcdcc30bf1041332c4ed7 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icf76cb69aedf4db01cd3444f4c4ba471 <=
            I4fb3fe065daa2708e55c812e57c19fb6 +
            I96f65790e2cacf7b529ce5b88598da00 +
            If077c67a062095cfe69f2260cee82833 +
            Iee5e74945ba15220f0f707c9c1927ba1 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4857b5b50556c8e7fff4b2d3e08e4b28 <=
            Iffb7fe9c74dfc01a43e99a099c4e7e04 +
            Ic09b4671e867144fe9f54a09e74c5519 +
            Ic0ae1191869e636f9e4391efe93309ae +
            I4d1c47569b0bc8c651c897ac8e88bd1f +
            {MAX_SUM_WDTH_L{1'h0}};
          I0a1e9cf99f1d4725327615f50fcc3ad0 <=
            I487b9b236d118786e475ccc5e4e56a6d +
            Ic46357bb77f6183329946f7e28294365 +
            I382153cec6f7d6258574e7c532186473 +
            Ib9d6c5be487a434fbafcda25ca9351dc +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie844f4c446983ce381b0bc4c0e8ef7d7 <=
            Icb92c7c10f0bfc5d287228f98d8a235c +
            I90001da8c360ccff128f637cd672ad42 +
            I5001118df37d08bd19d322aca8ff3996 +
            Ib0d033ba28e8c606ed92207049c76884 +
            {MAX_SUM_WDTH_L{1'h0}};
          I6067f47cccceea96ac46ff0d457b25f2 <=
            I72756ea6a4997bc4afd4bfde1dfb2d26 +
            Iea4a7766d3b9d5d030ade1739859ef0d +
            I78e1205de9119fac3ae8f43c72ac71f4 +
            I300d9f403e33d860ff5dde9f91bae11b +
            {MAX_SUM_WDTH_L{1'h0}};
          Ifd6fd1f3cbf8884ca7f64bc42278e4fa <=
            I63c0c8bef1dea4e499a16ce01e781951 +
            I5a7746e9fbb8c009f83ae57423296cdf +
            Ie0ce2826fd13b0e0b23c91e97787691f +
            Iebfe0fa45e4b34e142e82ddaa15243cf +
            {MAX_SUM_WDTH_L{1'h0}};
          Iaec9fd9e79371676bfa8ff14b4feae52 <=
            I275f6334127640b2de3f0f87f54fd74c +
            I3faeba79f7af7a006ab5cd256352e2db +
            I0c0be3347a7df9cc39997208b013f17b +
            Ieb778442bc855e93e11c9b13f1a7ae06 +
            {MAX_SUM_WDTH_L{1'h0}};
          I500757c4eda5d3d899aee47b87da585b <=
            Ie9fd8f7dc0c3849c0437a2a3d8607b4c +
            I45a6ef43e6e42594444adcbda26700ab +
            If36016df78d833c80e1355151c038225 +
            I57a393cc9cc9e1abc7962aa2cc840a7c +
            {MAX_SUM_WDTH_L{1'h0}};
          I47bf091b0fa74ad511a760bad9d2506c <=
            I002869e450d79649d27441ce00bfb575 +
            Id11fd3a31b70da0e64138e71840cfb83 +
            I0ffb8b65525af38861280645ac310e3d +
            {MAX_SUM_WDTH_L{1'h0}};
          Ia4c3d0cd9957f678880de5775de76e0d <=
            I8e01532a1ab9534b8de0474549d41a2e +
            I507e9bd0265d9ca6cd21a46fa21ba084 +
            I30fb41a57460a0b1f21065b4b97ddd42 +
            {MAX_SUM_WDTH_L{1'h0}};
          If5f957fa2f055b1c2c28e8d7cfe3e9ad <=
            Ifb19d75cfa0051107b5fba57bfc002b5 +
            I09faa07bf38acd96c4e29afd8a5167e8 +
            Ie8298c5c8ff538a3e37af46798f6d753 +
            {MAX_SUM_WDTH_L{1'h0}};
          I3608378a5da8c66bef58528d56192530 <=
            I79280400a4c9bed015106e5d006de757 +
            I1b01cadaac7d3d15007f0afe5c0ab0f2 +
            Ie7dc322fee8ca0b6b9659e5183e0d6d6 +
            {MAX_SUM_WDTH_L{1'h0}};
          Ie6dead855e00ea0a8e6a9b7503aaebb8 <=
            I6cb09ac924c3b3b44443263e08c3315c +
            I8741c5cc763512d16cb1186fa3323f45 +
            I22c15857572603cc24d8a87cb47c33b0 +
            I91bbec0523f77fc52a88ebcc49267e9c +
            {MAX_SUM_WDTH_L{1'h0}};
          I3bae5e6862e003a8b9a476f72cc6858b <=
            Iba4972a3b71a3101ab23190ed905dc17 +
            Ib38a46dc131d635b81fb7c196110fc4b +
            Ibc03a9b6115d0941ce9233df7ef2fa57 +
            I38ae79956762380fadc94f8126dc1c90 +
            {MAX_SUM_WDTH_L{1'h0}};
          I4431adecba8be9e5f21bc6b3e1f8cb10 <=
            I4bd98e902e805426fdd4606fcb5a5214 +
            I6b5720d71a0b4cd10ea34affa6631a25 +
            Id92d779518ae724b5fef5221372f8f26 +
            Id55a1ab9d158ea509e5f57286a3d1b67 +
            {MAX_SUM_WDTH_L{1'h0}};
          I21c7a2885126d532d00484376588a469 <=
            I43f52bcba1bd2e8ee5fac03320e4f19f +
            I391a2f354262558ff17d7d80b8c39e8c +
            I351dc309e916f282cc1e19303eee4112 +
            Ice615e7e18356ae4c3f615dd997be943 +
            {MAX_SUM_WDTH_L{1'h0}};
          I2c4d7339ff2fe68d060dd8d961dcab8c <=
            I9306d9ef7934ffe5902306b9783c351e +
            I70dc03a46e1ac0da826388abd3bdc503 +
            I72b4ef48363856af7faacc85eafbaf2f +
            I57b40c72004f2c3072cbdefbeef72b7c +
            {MAX_SUM_WDTH_L{1'h0}};
          Iee518b15b067eec58cccfa37f7432ea5 <=
            I2882ae2eb6d79a5b96d1ed937dcfd8bf +
            I0dbf900b4f430b4c1106aa86b640bb37 +
            I9dfdffbfdb83572cc3205f674e5db753 +
            Ie38351e19bdc4f2ce9caf75fc3937dd4 +
            {MAX_SUM_WDTH_L{1'h0}};
          I42145be9c2a80288ba4a2edd91f661a3 <=
            Ia8abcb8cf8d9ecc17c27ff015aa0b71f +
            I5bbbc4eedb7c61516769f429a8498ea7 +
            If49068db99aa9d09302eda27ab51fcb7 +
            Ibba6269b560db9d4913e1e515ed8270d +
            {MAX_SUM_WDTH_L{1'h0}};
          I9dc297ad41fafcda77f5347f331cfc25 <=
            Iec844d10736440b96f9d6c651e604efd +
            I7dbd1aeba00bb8b257990b7bb294211f +
            I0b3a936c3f7e0391111e696b2445803b +
            Ie392719059587a201c0148138ba2a2d4 +
            {MAX_SUM_WDTH_L{1'h0}};
          I846700c79f30ca954cc2933fc94d355b <=
            I02e672436ade3ee620c72c0d9ceee664 +
            Ie4d20df6b1e7a42f0df9a3cc26b12ac1 +
            Ie04e44d8e0756cdf34cf9ad53da76e47 +
            I4852d6bacfd82fef6fab4502d61e9a37 +
            {MAX_SUM_WDTH_L{1'h0}};
          I8af96a91457316e49e3f7dd5e57c82da <=
            I508cea40d87bec2672f980d145c89b55 +
            I80af3dcb716f3474a7257700aef89b81 +
            I6d4867d03d9187e95e27e99f7aecddec +
            I9200526d94c38e638370e9a2d7fed75c +
            {MAX_SUM_WDTH_L{1'h0}};
          I7d1c247500d7d32e406b2a5f7e2b745b <=
            I844b9a89ffb7a5e48979fdea546e244a +
            I9d05dc0e39e85c23b62f343a8de12e64 +
            Ie96877deef8b1676138f814c4a720800 +
            I15b8aa7d973edcf3b2365040f5570d82 +
            {MAX_SUM_WDTH_L{1'h0}};
          I66d85c030a8864505298919046056305 <=
            Ibddcc2e26fba20dfe2a2d399be2bc45b +
            Ic6e3847f035738243f4c5f71f296da57 +
            Ie9c5e7c98281cd1deb6acc51590c9d9a +
            Ic3f8e77259ee3eb5be80e11b607818bd +
            {MAX_SUM_WDTH_L{1'h0}};
          I4841257ae596d9d3e4eb1e6f886956b0 <=
            Ia5e26c2417aba1005971749f4ab2f367 +
            If6b40a030cb120fe017bf9d39e1a35d1 +
            Ifdcd91f925b63e0817798aa6e9200e50 +
            Iabf228f57ac154c417389f6711af1950 +
            {MAX_SUM_WDTH_L{1'h0}};
          Icd6f7ec117f9ab4eda8c5eba41386ffa <=
            I9fdfe73e77c384d33196c0f2d2a2fde2 +
            I30b5c7aadb5312ce96e833704bb3a320 +
            Ia18bdb8d2f02b50281f0acd4a45ac973 +
            If37de611ce4fa330c4fc9dcb87d4d95c +
            {MAX_SUM_WDTH_L{1'h0}};
          Ibc0498839d1d9b6dc853b8e5d7a88fa3 <=
            Id924dafd31fd0af0b28c7e6b7e95ec37 +
            I926c049036f53f0a0a6ad369de116c57 +
            Id0762ac7710c93249bc11c6ce4ae51a0 +
            If3c44eb85217da3b6bddb5aed97a9bb7 +
            {MAX_SUM_WDTH_L{1'h0}};
          I142ebca7f155e287e38ddf45423ab0fd <=
            I33703f538ec70268e6c00ad6eef6c4e0 +
            Ifc7eec6765af08463751db128f8818b3 +
            I9de5e90485b3f22e9003dc8a7b22a79b +
            I8c36318c45dabe6bf540381373f09fe5 +
            {MAX_SUM_WDTH_L{1'h0}};
       end
   end







always_comb begin

            I5deafec6e5f32da1bcf8f7018cf794d8= I5033323484d90d6bfbe03749019fc6dd + I8cab6f6faf0758f26d1a8851fae43896;
            Ifeb14203f4daf31c7701a6a742be57cc    = I5a11c8e7d2b7d4c0253df9015b7f3ab5;

            I35b3fb2670f3a60d165c1fd10f02c00c= I5033323484d90d6bfbe03749019fc6dd + Ia3f7f07ddb09ea33218afe14281ac3c6;
            Ib581c19864deecf01268595049268b19    = Ib0740d8c9ab158e682432a0e3ec89798;

            I68925439e233444a4da44871f31de94a= I5033323484d90d6bfbe03749019fc6dd + Ie23ed3ee61f468f59f2baf661cb7f85d;
            I661d84af541e30828bcbd962d72baba3    = Ibb6505392d5b3be76542bb0303d46876;

            I3108702b5ca506422c1ba6174619f193= I5033323484d90d6bfbe03749019fc6dd + I79458089b042e181e37cc44c06d08681;
            I1c6928cccb4bf7ea7dfd74e425b9624d    = If23edf1bc3801016b24252fbc3d33508;

            Icc8e8f6446ac64350a05f5e1e0541bb9= I5033323484d90d6bfbe03749019fc6dd + I856eada207c5006beb8f83f01d5d74c9;
            I6eabc5c074fb1e2183a5f1ecee87a518    = I47478ccbfc4c3b944d130a192fb4fb5a;

            Iadebaf3f6cca1ba78feab50ce70c8aef= I5033323484d90d6bfbe03749019fc6dd + I1ddfd31bbf062aa5c3c71d61e492e3a2;
            I0107769bbd7c239685b4818731334437    = I40b126fdab110e58eac80ea13bcc699d;

            I8681cf376dbeceab29279a7637249e7d= I5033323484d90d6bfbe03749019fc6dd + Ic5e0a84cf1a2ef907b2456559ea26c75;
            If723180430080198d18a08d6775ab208    = Ib12b389fb2603e428b72d1e712975e40;

            Ie850a07565bed90389bb125ddcd39658= I5033323484d90d6bfbe03749019fc6dd + If367d63311c96726517240de13bd2a4b;
            I44abc734d6acf92a8e8209186d7a1676    = I22b0cc5517631526be6455fc60dd5323;

            I97b77743c2311ec629ea24c933b60053= If5dad13ac41b3034bdb034bc86c9b348 + If49f97cc0c42b23ce393b534015559a0;
            I72aa55988d58c664f3291b5786fc8ceb    = Ib8aba28214fb9ee1693cafe9175831e1;

            I07a0a8d41ed8176e92380f2c89c2afdd= If5dad13ac41b3034bdb034bc86c9b348 + I6c4ba0863ab4c8d1a56324a4d89ccbeb;
            Ie69528583db8155917ab3d32a446de04    = Ia03282a7ed4a337981d4f5b01f564a1d;

            I021842328f948a94159b32903c8bcb68= If5dad13ac41b3034bdb034bc86c9b348 + I5a3297f48e1045273db6522744582b05;
            Ib22b47d95b72871e74069fe80a191680    = Icf75bf863d8867b0fe354017921aeae1;

            Icaf3bd685005a05c8fb334266ea4e4b9= If5dad13ac41b3034bdb034bc86c9b348 + I326660e98f61bb2ced4c23c7bcc9324a;
            Id9451e945bd26b8dcb4cb83ab4ade73b    = Ia65c174738acf41b82f75be972e9022e;

            I92d9e1d7dcf45a4d738c546e959687c3= If5dad13ac41b3034bdb034bc86c9b348 + Icdb143a4ce96029c2441758bf2edd7b0;
            Iba4627d3d3ef91f168068ed128c04113    = I587a0e70cecf4d054cc0ab53150876e0;

            I39ca3a8ca714a9726114326ae6bfab0a= If5dad13ac41b3034bdb034bc86c9b348 + I3c6fb0df5846a19228a4e6cf9f9106ac;
            I39bef4d462b0a3f88ce1485a58d66da0    = I7dc71f64f9b3940721569574db6e18d0;

            Ie9ae20ed5b2a0cad2c37c5bb2ea05ff4= If5dad13ac41b3034bdb034bc86c9b348 + I6a3854ed571e8c262aa3ec377c247778;
            Ib95e457d5ae9fc89e197c249414abbcd    = I935ba9f8f6e9c68f75a7cb576655cab5;

            I8f131eb6138c23fdcb35195703131e64= If5dad13ac41b3034bdb034bc86c9b348 + If19dc22d45cc4664c85a043ec4c00617;
            I2be28be47a38e9ca9d3b9167327d3d59    = Ibdc981a062c989ada978f733ddff0f71;

            Iff77e08da4bcbb85b95fa277b69653a9= Iac428f9f798618e1ef495c626c41892b + Ia7f53f0cd86055da72c13ac474f052a1;
            I2ee6154b613d0d86c2354604e93a9a57    = Ibcbc5e2720516c24359870ac790373f4;

            I703e0a4879a39b3b8b0a49de86ca4ff4= Iac428f9f798618e1ef495c626c41892b + I0cbdfae6f75a639eb591d9c0022f5838;
            Ia7479d4940b575cf918cb8421f041e44    = I11fdefe51f8f028fba7698870d198df6;

            I3da217f6f2d0f515bb9036673d753a88= Iac428f9f798618e1ef495c626c41892b + I1d0f031e8ae9c0335d501d1565118220;
            I3c5b1cddd608ad869e0182ad68bd0494    = I10f17104471f87c53a589926534fc9fe;

            Ifcc06d5a010e01a781ae8a9e9e2b31a0= Iac428f9f798618e1ef495c626c41892b + I4b66c202450986ef0df05e979cc8bc7f;
            Ic4425ae997c479e05e12347a803213dd    = I8fdaa3f282af2d5f053d77216c659146;

            I42fd611fec087113ba6e35f281bced9c= Iac428f9f798618e1ef495c626c41892b + I972bee4216f8e532e8fa4bd25fbb9c57;
            I3a0518d0d382758ae579acd7e6cd634a    = I167ee185ac7beee082544897898b27fa;

            I5bb626e7347bb9ae4219cc72244b38f8= Iac428f9f798618e1ef495c626c41892b + I1182655739d7ab5bbe4a6546a5ca36fd;
            Ifd28c1cd286b7a483891bdd094b70db1    = I5264a25f96edda24a763298d92cdf8c1;

            I47e2dac0068652338f94ddffd2dbe88a= Iac428f9f798618e1ef495c626c41892b + I195c3a82123142d509886ee37dc6fc98;
            Iadf7734be049c645819d9d023b58c4dc    = If7d5260450e23711760a6f9e5f7aa820;

            I59a3f06de2984078a4d4c430a2980fe3= Iac428f9f798618e1ef495c626c41892b + I96ef4b631a7f63e19f67f3920685f0e6;
            I5f23af0d0853ea6de084ccf77702b78d    = Id1265b30a8ed85169b1837aa1b656aa2;

            I857b7fd58279b1063a06a4f33b880ba6= I5a6427c8f18b36d2ea18fe60a0831ef1 + I5f68368511b59d2e365cc91b806b334e;
            Ic5c99c42e9ebe5dded369ac78a1bedb5    = I84e6c5099aaef8094f4c2bbc82989c4c;

            I3901bbda029cd0a41640001c1efd400f= I5a6427c8f18b36d2ea18fe60a0831ef1 + Ia6255a136d5f36ea6cba654bd5823850;
            I4f2498bec0e96802b82f0419d97c527f    = Ibf4bfa16424f7051e80b2947ff7f5533;

            Ifceeccf10f1d85a32f70c04654a1a1b4= I5a6427c8f18b36d2ea18fe60a0831ef1 + I21594c8b0169efd7c2aa6cbc31f4a901;
            Icaf86e0abee612aa972388c0b6f90763    = I0e138642d8ed7e30cc254d4e259e3d51;

            I2d810c1d1304658edff74921e8d0f388= I5a6427c8f18b36d2ea18fe60a0831ef1 + Ife123bf57fe693dabe6aeaa236c4e058;
            I478c4f13c05651605a2045bb5fd6b60d    = If1c79ab7bbf50d343ba3f758a31d6786;

            I575b0201be445388607ab83465eab8d6= I5a6427c8f18b36d2ea18fe60a0831ef1 + I518a2736384c14c02f27bfa3d8ea7aff;
            Ide67911b52687d67ef0c25f2aadf14c5    = Ic2d209d919c7e43f467c3f2d093c9a8c;

            I7928c5ce0f821df1cb6271d15e19fa22= I5a6427c8f18b36d2ea18fe60a0831ef1 + I2dcc0d17b9fcac35693bf32b5c5540fd;
            Ie9e7630af25f39a0e820181918edd029    = I6c59651ae65c67edfa963ce797b98234;

            I12695a21c942d02a432cf6382d7d7452= I5a6427c8f18b36d2ea18fe60a0831ef1 + Ic0819ccefe784a6379716b3633ae0196;
            I0e1f07f30cfe36f189e9dcb4e713b5c8    = If4b95101c6d8670411a018ed1ae697d3;

            I00d03f0f71b008dad8035bbf251f41bf= I5a6427c8f18b36d2ea18fe60a0831ef1 + Ia540866403683bc30504bace19bdda7b;
            I31cee5e2a93635987776b0ea477e6211    = Ib1e406a5bb0569ac2c25e7021ec58edb;

            I41afedcbc0f492e3243436cbefdaf609= Icc29441eac6ca7a138d45743d37505e3 + I915054f2fbb8b93516d8748a3e3e29e2;
            I84721f2bc5ae10db78d2e7e07cc28d94    = I8198f75286b8c817d3b69cf7537b1c38;

            I638c4c2708e437a050ed7cbbac516a59= Icc29441eac6ca7a138d45743d37505e3 + I42460fae0acff25fa2b829e39ddcc4fd;
            I6c6d057e910da53aa47441566f95153e    = I9431b10311eda8240d91bed96a969523;

            I6877d3306b1f08c236b5d1b59f0de259= Icc29441eac6ca7a138d45743d37505e3 + I77a94cd9186ca546ca9664942ea3537f;
            Iecbf70768fbaaab8da98eaa9a2b956ee    = Ib623d99c3d272f39c518b6a41dd03e8d;

            Ib3e66aa460f39d32110ea6f115785b3d= Icc29441eac6ca7a138d45743d37505e3 + I9a5388f8aa6e9924a309aa8db4c1983b;
            I71b8492d70b423e95938995c07395def    = I388b66a7b7e9225f7aef4699521e9250;

            I5e603e8392a5322951b3225b65b19446= Icc29441eac6ca7a138d45743d37505e3 + I3a76f70ca3bfbcacc6f3342aa71f1912;
            Iae469bcbba9598bb46aa7ccf9fa06a37    = I532db075ab1b0a5a37a2085ecd0611c3;

            If5da7fa1a615e1122445460e33487772= Icc29441eac6ca7a138d45743d37505e3 + I46e9c76b19ed1ff21f102efe6ee5c732;
            Ie2e854376f4b6509ec41507401173269    = I357c21c29061134ed6e5c872836f4759;

            Ic4153dafafaf7d047478c5d81109437f= Icc29441eac6ca7a138d45743d37505e3 + I3096d11098113da669ee0a94686e600d;
            I7b1401c3c2c389d9bf05658c88ff6b40    = I5a1d671b8b8877192d2c129be7f149c0;

            I7b5476007f04e81afc0125e6a8930303= Icc29441eac6ca7a138d45743d37505e3 + Ie6764a631310e312ba5c2c1e601d828f;
            I88ee95aeb6c744eca0e127e8497b5dc9    = I4d1c830053fedd74930d9992732e9542;

            I3521a18022925249caddb8e37d2c1262= Icc29441eac6ca7a138d45743d37505e3 + Icc6d895d943e14f2801c22e79ce190e8;
            I5573e18ade3430ef3eff5e6d960e44eb    = Ie53c31ded4a5c8977f956e968dd5a9a7;

            Ifd0f52d4f814e2bb4c3bd34c1e09bda7= Icc29441eac6ca7a138d45743d37505e3 + I9b09b800a9dcd8ac36f25cb0324e748d;
            Id6260fa8a9be077673e82344c736b1c4    = Id5355c3ed75d1aed52250f6f0d00b1a0;

            I8945f6d420c8b373225451defcd2c805= I0e7754dcbc04a4850e052ae4a2fbe328 + I71e4d98dca37256fcc84248a26d703e2;
            Ic052eadb342350c52d89e73d5fea80bb    = Ib43ca9d864e41a89bec5344ece17fd10;

            Ieec6cb6518cc0d9300de0c4f2d32487d= I0e7754dcbc04a4850e052ae4a2fbe328 + Ic6fa98631d742b27f252fe7c95caef55;
            I98b8d024432fc54ebf2f15d99968f2e0    = I6c7b0be00e8302794aa3a79fb2acf100;

            Ic62eb7e90d703ef994e68587345a4293= I0e7754dcbc04a4850e052ae4a2fbe328 + I20c65000bbc10299168af7390776a03c;
            I98f54ab8454940141a484332f2a05369    = I144843095a5e8952e26bb5c9943f0cad;

            Id3efd8419da986aa89b8ad8e75848cfa= I0e7754dcbc04a4850e052ae4a2fbe328 + I66a304016a9adfd85a2abb6f8fd39afc;
            I9d94ad2da06ac1fef4da7dcc56abffca    = I0b6cd5372e2cc6a72c1c8f984279cb69;

            I40803f10b7c4dc9ae4969739349b0265= I0e7754dcbc04a4850e052ae4a2fbe328 + Ib303ea0240e7ab5f000dd10e975b2274;
            I51262e3abe460148e3c2d2b74989c2b8    = Icd143823913eb777c0cba42d8a5802e9;

            I7d961743fdeaf1e72e4b25c12a1d4c46= I0e7754dcbc04a4850e052ae4a2fbe328 + I5dfc71255cba279420b7545df4d35c40;
            I560583680bb2f5a0b5ede42ceaafcf8b    = I02a575305a6112f734bc3ebf6b883b90;

            Ifea156f33eb61fece272efe379327f6e= I0e7754dcbc04a4850e052ae4a2fbe328 + I02330ade2eed926076cc071e45eed82c;
            I389f83346ffaffe8186fb0074d71f43c    = I20f0ea42718bdd84caf3da4a1b32c5a1;

            Ifc99169b3399f3d14121c1a9bce3fc21= I0e7754dcbc04a4850e052ae4a2fbe328 + Iae9e023628eb6686708b2656f15616cc;
            Ie89c2a1b3943d12197bb972bd12595b0    = I11489ad40e6ff10933319784981fe59f;

            I6536144383cbda6f3b3c564391866906= I0e7754dcbc04a4850e052ae4a2fbe328 + Ibf482db0f5058be72061267c42ebc292;
            Ic7be56919976a2d1088114c21c3c1ffb    = I10fe1f517735fad803f3d5d75fa3d406;

            Ic21bf9a8a4cd85ec123d7fe142ed49c0= I0e7754dcbc04a4850e052ae4a2fbe328 + Iebdf938a28594624f4d4a337356485cb;
            Icb5dab0df062ab46bd3d1a73e85ef4c2    = Ifed41503f4acb3625530d3c74b5ccb52;

            I1f31fe6a0ca8510bcadbc2069403150b= Ia30c019ed8ce395556494a92e7b42a92 + I6ecf7249e6151477fe74a79d0b126b21;
            I27a568cfc2df13cf689d366a25e5d05f    = Ic9550361e9ae769b5095df4857041e60;

            I0e40933d00f4a7d9b53b2764aa0da700= Ia30c019ed8ce395556494a92e7b42a92 + I737daf208eccf95feb3192897586cdce;
            Ia6688964078f1ea87b742352877aac45    = I29cedb22eb565264529effcf107e167f;

            Ic41a6e00bc84bfc1b8194d15bb899c93= Ia30c019ed8ce395556494a92e7b42a92 + Icfc1c6d96a3598af73e99a350c387d72;
            I180deab4fe0d03104cf2ee035f6a9b8c    = I229b8819c94a612ca986936c96ffa9a9;

            I2832571f2b0a7fbb41d2e8ca7f64e003= Ia30c019ed8ce395556494a92e7b42a92 + Ie3e0c0e40c7a67ce7f957e74bd2a895d;
            Iff6cd034bb64d13c21910c11bd92266e    = I62c0db0621c1a71960770d14c332dc0d;

            I9593c853e41952e408a809cb24efa4fd= Ia30c019ed8ce395556494a92e7b42a92 + I847cf7ff866f8a666872c12d6b67b1b1;
            I7c34057a77f2bdda93c422506959818d    = Id94e17f3fb5b4fe7a5fbe8e25d02ec27;

            I6edffbf4136e193dca0fcec3a74e8e9c= Ia30c019ed8ce395556494a92e7b42a92 + I954ff0f9ee871a31774a3d786128fa13;
            I7ff7d3fd63fa67cd72d1591c1a373180    = I10cb83fe0a939bf2784eb93ca1d7b3c5;

            Ibaed50cc2e36ae58945887d11a6ec9e4= Ia30c019ed8ce395556494a92e7b42a92 + If8b0b96a659183e3651c691a2848b86b;
            If910e75bf10cf02a5b414cbb4fad1304    = I8f8b2e93ca65e789d13d66ecea733894;

            Ie4570cac44f59e6ff46f73a703026479= Ia30c019ed8ce395556494a92e7b42a92 + I7168b0efdd2fae57292379c9d15c62eb;
            I266697a6eca2b73a76fd375a0ad72a05    = I2527b288272a0ee2127436252a47a6aa;

            Ibaa136d37936687e9dbe4222749d19c3= Ia30c019ed8ce395556494a92e7b42a92 + I9e2de71442b8f504358e582087a6d19f;
            Iba188abd7715fcbdad3b1f3d985c6fc3    = I743dd733d1c20868da7a802ea99b23bb;

            If85de3225f45478827b43b89089cd29e= Ia30c019ed8ce395556494a92e7b42a92 + I3e265a7dcf29687248b9275df49771fb;
            Ic60c640562e3e45c89a1de78af509b6a    = I5dacf7fba8d457b393930fcc76135b39;

            I0344b86a6e9c036e103a9c1f3651175f= I9799695ea8244992a6694eaf5c8ae64d + Ie932a22a7f1fa37087cbc9e8d73efef4;
            I0456494b33e4ec852c123cb3003b9886    = Ic50ab0fdec011923b02c0c0d717befa5;

            I5463d13575e0b9fb8a0f6cc8b35d0ce9= I9799695ea8244992a6694eaf5c8ae64d + I0c0d844fe3b7d35c1ed6bd7cc4e0dc24;
            I2ed7c217fe3e21fcb27e04f68b95dd6b    = I3afc7e76861fb1fa36291ac8d5508483;

            I8a3c63ef122001a29e5abe93c4e1a48f= I9799695ea8244992a6694eaf5c8ae64d + Idc77c7d5123717fc2596a51d904c6d82;
            Ifda5780b42bf451a7ce834f17b3fdd20    = I7c06d7efe631bc01f98ca137df06876e;

            I6a79108484fcb192f6d93bfb98e271c4= I9799695ea8244992a6694eaf5c8ae64d + I07048dc5cbe24ff72d24902d572face0;
            Iadca92fd39d1fd6032feb8415ca5246f    = Ifd5f5f8f7ac4238cdb3a5fb2e86eecad;

            I9001e95b71457a2bd09a9846af370b16= I9799695ea8244992a6694eaf5c8ae64d + I79a46279070c53678a5af54f661c5821;
            I613453382f19dd7eb9bdf51e945a33b0    = I17e9d58c80d0da6e6093836deecfa743;

            I51620de618db6327358a5cac97e1e97f= I9799695ea8244992a6694eaf5c8ae64d + I5e8ecdbb018402b2fbc0049ee44bae8c;
            Ideafa683e6a3a38848fb8bee22eba11b    = Icd18edbcc227111c037023bf2b57ee5a;

            Ib9c58818059af5c5a03e77a5dcef4654= I9799695ea8244992a6694eaf5c8ae64d + I9aab16e89f1b64117caece8ca8af5940;
            Ie4226e7e17c7971f07aaf0cfaeae495a    = Id22f8eb74ec1e8499e150278e438359d;

            I8081c71aa01a8d575bfea6ea7f2f595f= I9799695ea8244992a6694eaf5c8ae64d + I8110a5a62607093b21b7cd088b1d9ee0;
            Ifbbfa268bd4c31c7eed45cd43fe6a405    = Id10ed140128d500e98d984a15b479fb4;

            Iad999607ad8d7da0f3b341f83ea030a6= I9799695ea8244992a6694eaf5c8ae64d + I05fb1982415bd3fa78dd9a00af7a3d4a;
            Ib2d99d95f7a31e4745211c5ff96f851c    = If89f8e436166d9beeca9937c45b2c7d5;

            Ie7291c914d2cb66f547b0a7717f71311= I9799695ea8244992a6694eaf5c8ae64d + Ia9f375709014a9d553d46cff2799b59f;
            I692c0a91b415b400a3640e2d9a40edad    = Idfd24573e271b5cdd6f051496cb6ba8f;

            Ic01018a5f1bc392bbd267016f6612a83= I4524cd664b4cb41f642c675fa484c84b + I3753b2c4ba8f1bee70def390a96586b0;
            If8c4dc70212e8873167e1cad8e8e5692    = I145c31d89636b936f18a19bf50966bbe;

            Ib11dff839e7e532657b32f29fd9b1651= I4524cd664b4cb41f642c675fa484c84b + I4dbd1bb8f1641f15e3a4f1e309962811;
            Ib2f75e91bf9e1d32a3f170fc85244139    = I15cae93770d041e2ef681a81e8256059;

            I251d7ea16dd5407d22a6846ddcfe12d8= I4524cd664b4cb41f642c675fa484c84b + I29c8133231cfda17668bbe7b692bdfe2;
            I3606dc61f24567cb1ace443cea62a43b    = I6a86457e1b16bfc515084fe599281818;

            I773797f81f73b9b6e844441142a1bb48= I4524cd664b4cb41f642c675fa484c84b + I779da979707d9712c1626d6025f97599;
            Ie402c9f793b7306323efb8fe23533250    = I2453c39e5805313c3a8fd0d074058916;

            I853ecadf30fc10a13dd1ffb1f2dfb5d6= I4524cd664b4cb41f642c675fa484c84b + I09a1d04c307fcb8a0e30925d86df3fe9;
            I54652565023310e2eccfc4cb87c56b43    = I34636cc42b16776295078bd349a76ac6;

            Ibb8b3c91e1d3b890cfe58f32f8ec3ae3= I4524cd664b4cb41f642c675fa484c84b + I2cefbf897bb7f6f67ca500727e85c683;
            I616b7a5987edbc001e0ae1b638f25a39    = I48f8d5589f772fbb4b3923fbd213e7f7;

            I3485d69de942d64e56925da522175b51= I4524cd664b4cb41f642c675fa484c84b + I74ac0327175f50f508a5013df298df02;
            I06604bac478ee906b3fe8ff307cdf046    = I83e4b71b0a0a3a82fc0a9fb56f803fa9;

            Iae42f12bc0475c8b58341d80027a57cb= I4524cd664b4cb41f642c675fa484c84b + Ifebfa58419ecd22a334ed4b67f5c3581;
            I135dd8a85aca863db660f2ad4f80ca2e    = I2abd0942d4d5e3aff2d24db9656c025f;

            I22fe2af25463f87ee7315a9aac32854e= I64e959d80af111ed2fcd54a5407d21bf + I2956687a5fc2fba7149889624ef85647;
            I8715d73b58270dfa33b903e9cfb50be8    = I0fa19f52fef5a583890e3096eb23f1db;

            Idf44ad78c338c39699721ce511691dfd= I64e959d80af111ed2fcd54a5407d21bf + I088898ee932a96c14f2f0f568f5455b6;
            I7f60cb59895af6d314f5d0f401c80350    = I0e4a9bf26a9df3551a69edced6128e30;

            I984a657f9265d41318c0290e249e9712= I64e959d80af111ed2fcd54a5407d21bf + I2d9632ae6a0f3ba44c3da8f56ba3fedf;
            I3e25e6e9de5ee9242a472ce957056762    = Icd359ef9d3a983f4258cc4441110cc97;

            I915fccfb1d1ada9aa7c8e24c2eebd04c= I64e959d80af111ed2fcd54a5407d21bf + I3c0ddec25c53c166d30eb78d4518840e;
            I4c5f36517aaf872e7f05de2f7f76a6ce    = I31d6000373f248b1dde9fc0108bfd280;

            I2bdf58ecd0974720631be830efb48dc8= I64e959d80af111ed2fcd54a5407d21bf + I296bc392d4223cbdd6f77be6523df819;
            I0e993e6f98616632f17835a2994f45e3    = I445cd3125f69b7e29d582a4803709c8f;

            Ibaedf6246fa43acc8accb5a24d49cc2f= I64e959d80af111ed2fcd54a5407d21bf + I05028975b49ec0c089bd981696f85a8b;
            I281f996740b16568b9d29ca41a3fa50d    = I2a8dcc8d3db0d8b5bb54bc7fae5e6ca7;

            I904d13524dcdf55478a5266d50e53ff7= I64e959d80af111ed2fcd54a5407d21bf + I3fd068d55154441ffd005999ea823fd0;
            I55bbb73d68871d9dbce4d590c029aeab    = Ibbf4549a33d4916489e7e325a811add1;

            I22d8e5d57c1bc082169437a654d22bba= I64e959d80af111ed2fcd54a5407d21bf + I066cd52173ec5dbce9a3f470d73325af;
            Ida491561008f4984480d1b0f09d2fa77    = I9a2d80bf2bbc2101c8e426cfc1c8277b;

            I719cdaa2a2e61a0df7f1fd5efe517426= I3e0da4bcbab4804b5397fb3aa2c94f51 + If257757fa31c2f4cc9ec322e4ecccf83;
            I624e237f248d292c0417ff85056857b0    = I71c9904d29e88f0a5e6d7f8ec88de592;

            I8e92a61eb73c41680652936cfcc614ff= I3e0da4bcbab4804b5397fb3aa2c94f51 + I2b9584392ef9a7828ff57bd4c522a302;
            Ic7c1fd79ba76dbb254c6183017f40b3e    = Ic6c8869890916818213809df90b52856;

            I7ad5af8319f6da469858300f0777b580= I3e0da4bcbab4804b5397fb3aa2c94f51 + Id3670a6f05d40ab69624544de92b9c64;
            I546d683af76dc209a5205c6274abe908    = I3c61b092287e1f2c446aa7346b3dfcfb;

            I32be72eaf04e79120a57ea94296a4e56= I3e0da4bcbab4804b5397fb3aa2c94f51 + Ia840e19ca36795a50ab1a6e6a1729edb;
            I7b4bb785489c5bb22c84d9778192fe44    = I8f94e1fe9df14c5dd75421cdfe8b1efe;

            Ie756f6a87d85adb40479ce7cf3545556= I3e0da4bcbab4804b5397fb3aa2c94f51 + I87d958c00fc6209d901147831b0c951c;
            Ifc6af7d7aeb7162d554b8604a44f3361    = Ie2a432bd8429925297936c8aebf7282f;

            I8794c6ce0a3f2e6697372e2c911ba420= I3e0da4bcbab4804b5397fb3aa2c94f51 + I1abb512ca0383c9e7104418e07281841;
            I5b650c4c3291670b480a7f1095093dfb    = I309c99cc023e0c7804b2574821d63f10;

            Ic82b1a29b5e63bcc3686a0d4bf1f5c24= I3e0da4bcbab4804b5397fb3aa2c94f51 + Iffd94cf3a8a4681ff3327c90bf89bd8b;
            I2f5f88cb5e5e4723bd8a83c5fa80cc4c    = I5806c65240e9ce9f9d0804d063c2674e;

            I253ef976058080beab79646af18e2d5b= I3e0da4bcbab4804b5397fb3aa2c94f51 + Ifb8b3586a5b69b20cf03eabf51344ab6;
            Ic174b361182c98486e65b7f87b073274    = Ib73d05919f3373f122b121be5a038f4b;

            I930dd54c36540d75dc870eef89960163= I3740b30d31f3c61d93a14a46e3199c4d + Ib8380902ac4082f834744ddef6d0cc6a;
            I7ba2f7201745258dbf224de087a25233    = I84136dfec9c8ab98228801deffbe8c19;

            Iaf7554cd4e8b5ea6155ec61a8d589b86= I3740b30d31f3c61d93a14a46e3199c4d + I25aefb53f59a00abe88b9dcf6be6907a;
            I131a4bd335fc23ee10f7ccb1881ab9cd    = I09e9850f90a7f073169e66c9e2339f51;

            I50907c7d1efa0038d81efed82b192891= I3740b30d31f3c61d93a14a46e3199c4d + Iab6d0f72579687407e029c630b107f7d;
            I90cb3e06b42f25956b788a792eef371f    = I1260922a3e6cd464e43f215299d70ef1;

            If3e9486d2960d164d94641d4f1917416= I3740b30d31f3c61d93a14a46e3199c4d + I523e9b6f828ec7f166750112f8a3f676;
            I56302770a8d56932e7bb5dcff56c71e2    = I97cf4612b19722d7f5f4cf9a867a9b22;

            I2bec61db45dd79b98d6ebff6c5a4899e= I3740b30d31f3c61d93a14a46e3199c4d + I343df614f97cf732e57cf2ad3f95dc9e;
            Id3b8c058b3838c388eb5ddcb31dfc799    = I4856ddf90e056e12eb6ec14d66f776b3;

            I7f31647f3ea6ce7bbd211c25cf4828fb= I3740b30d31f3c61d93a14a46e3199c4d + I0c4bbd1827b1859caabb067e864ce4b3;
            I7ca8ce63dfb821d10304958bada71737    = I370986beb4c411ce7154bb1c7045c5d8;

            Ice65387e606faf9c7b884475b489abba= I3740b30d31f3c61d93a14a46e3199c4d + I34d428a56bd0142a9be9f627f1c3c87f;
            I06ad44414b45d262f9542015d2dead8d    = I0b22c5487df5e2b47d2ac3e16ca195b9;

            I63f914927dcf49552e9f3fe0180a30e8= I3740b30d31f3c61d93a14a46e3199c4d + Ice66c108aa66981051df71e226cb0e4d;
            I833ef4acfed17e4699d65cbaa3e7dbd5    = Ic7437fa32ca344b6eaa895d35d335e57;

            I742ff5725e3a18acd03454cf9f313f4b= Ibf0a30abfec9031737eada436ac1a0d4 + I6c1235e88ae444a96ea64fd1bfd04d8f;
            Ia77e3db939408af719e0a8555dcb68ed    = I1dcfffaaabc223ae08cd9d08d6e968d2;

            I84e4b3bc63ec0b0bff7f98f433c1fd67= Ibf0a30abfec9031737eada436ac1a0d4 + Ie2c801b2de066c3218d7312615b7bfda;
            I57ab4999187992eda55a82bf0f09b31f    = I16bb10e8ddda86c2c8a1df7b0ec4c133;

            I78c6a1428a1f211c5e89b8c76b3dc033= Ibf0a30abfec9031737eada436ac1a0d4 + I7d98d1e5f07fccff5f20eaca6363c700;
            I21f7b5402ae8e8954d99931bd5108250    = I50ab3193dde101b550b508744be5a775;

            I9897cbf9d7cab759f99f5f8f4bc125d0= Ibf0a30abfec9031737eada436ac1a0d4 + Iab3876e5107e3a56b1fafe41e16d9482;
            I3627708869b47d460182bc5040092f9a    = I022ed4e5e55e9c3cd418bca5475beb82;

            I9a6c1ff6dde5141849e4aa925140ebb8= Ibf0a30abfec9031737eada436ac1a0d4 + Ica807adc510a2e32580ca77c18ea0b45;
            Ifd88f0f0abd1c037434dc16e34550d2a    = Ie44afe129f71022f34e9f9cb5ac4eb3d;

            Icc1c25b229393361f1245c40f573b423= Ibf0a30abfec9031737eada436ac1a0d4 + I31f6bbfbbbd4c20d0c5c71663da1d4c1;
            I27eec53da48406e7e1202345a0810e08    = I38c8f2c90a4d997e5597b462e7e8c613;

            I53b5a72e41ee53037ee3ae040799f401= Ibf0a30abfec9031737eada436ac1a0d4 + Ie4e4eaf3e5d2f581210af8054df71c6c;
            I682d42afaaf103550ce4fbdba6192c88    = Ib38a5e546fdc5837a97c4ff3a627777d;

            I3cc25fb583118f45babf457fe78d5434= Ibf0a30abfec9031737eada436ac1a0d4 + I220f8e45e5fe6e69f02cded87f12e1e5;
            If225534847db8723768941c3819ed7c0    = Iaebf3465f121a3c054c87227d7e9e167;

            I20c046dd8a1265e12e902275b73417da= Ibf0a30abfec9031737eada436ac1a0d4 + If47be2ca4617a426258c51f8d977ba3f;
            I43a91b2232a47d1f6731bafc15ced5db    = I6fd1108c6ac90f5c69db5aca76055a32;

            I1b184c9a34aeb6eda813d86556e235d9= Ibf0a30abfec9031737eada436ac1a0d4 + I71a28e8525f07dabeabe4b4f45f353d0;
            Ic54026604afd19b0c7c71ea1ac0f1c4e    = If6f92d3b43974c88963a188a26bc3009;

            I70e03db993e1d26d5814ff5fcd38ada1= Id36e8953a02400a5ab1f4dfdb0422e6d + I22c3140a8db02352d2e2a2a11eeba117;
            I218bd69f079aa21f0dda241ae6e387ad    = I19fb6cacc6841dec5653ef273676f18f;

            I119dc168a44950d215af877eb81152fe= Id36e8953a02400a5ab1f4dfdb0422e6d + I15022e1b349eee259d3567837283dbf6;
            Iaaacca4d06ad0f202d839fd7674f1829    = Ia0abbf270f98b4bf4f29b56611db23b6;

            Id717ed42457eb1d3f4e3edbf0dd72c41= Id36e8953a02400a5ab1f4dfdb0422e6d + I79259217f63b2f6263552c434d0e5c93;
            Iecddac410bb2121da0df2d73c2d23cb8    = I38ad3c494c777f3985d61eef7cab8fb6;

            I79d1f852a03bcc11d6121a12d8c5b86d= Id36e8953a02400a5ab1f4dfdb0422e6d + Ief76663994991118b1899ea4ddf4527d;
            I1aabc0c0b7b602297ad592ae48b23452    = Ieb8d87fc8ecfad97cb9840b3739d6ea4;

            I769e650e49f152c0803b06232740691c= Id36e8953a02400a5ab1f4dfdb0422e6d + I9470c7ab9634c01bb832c9e4ff5496bf;
            Ida3aaf7237b1383cfe95eeccf3971a8e    = Ic1087bae156ef4dd5fe218537432b0ed;

            I1ef3c09b8481f14c3526224430a5f4b9= Id36e8953a02400a5ab1f4dfdb0422e6d + I06d859184884c07a14c83d2f06587ad5;
            Idd2a8ed39edf6697b0988ee4eb4f2d95    = I6655118cfe24b706e6557438ffa1711a;

            I2a38d43a7e25050aa672cbf84a409aa8= Id36e8953a02400a5ab1f4dfdb0422e6d + Ie02de90d8eb06b16314946d21299500c;
            I735c660d5232e03dd8fb129e2ca4b445    = Ia12b8e62d6e1d52861589818deb6a851;

            I1c2be5e13c462a8a6b07bca311582ce4= Id36e8953a02400a5ab1f4dfdb0422e6d + If4b100d26126e460c41b8c1bc8fbbb96;
            Ia04d6065987df3f007658614406cbc28    = I59260857d96064096680b8361521b588;

            Ie8fd61caf16aa0e504cc7dc8cec6f0b8= Id36e8953a02400a5ab1f4dfdb0422e6d + Ife732309efcc740cfff5c747aab2e3d6;
            I7aeddde5b60828ac7f8b6c2addaf220b    = Iee39a5d6276b276729abd14472262ed1;

            Icd0fe98ca873ad6dacdf80dfdfc450ec= Id36e8953a02400a5ab1f4dfdb0422e6d + Ic7ad59f6a232a997706d17b4098e0324;
            I150c28296847348d69cce123f20656c3    = I20aa2879f47abd3c368f7494d944222d;

            I94e1ab698dc93ff0764dc5c1e62179fe= Ica71108a53bfcfd1892b4d03ef68110c + I26781ef851ed43c6f88ff1215cddca6b;
            Ib94d38d19b3791fa2d1b42fdfde8435e    = If0192b9580e5fdb8d71b422ccb28666f;

            Ifd48363af9abb390a72991fbdd6f7877= Ica71108a53bfcfd1892b4d03ef68110c + I68e58664be09261e5a80d6f8ecdd1b60;
            I94865622898b2e481e86a244f7aa2759    = I5095a3f4dd1c3bca218d17f5c609b667;

            I44f79397a010088e4ecdcb9669f2efbd= Ica71108a53bfcfd1892b4d03ef68110c + I97aede8502e443f98938487a5a5c072c;
            I1a4a432e735367f515ca747cef7d7d04    = Iea2a2368935757fe57b3d283fdccdb3e;

            I124b0b7d91cfb42b0d9722f3229c2d53= Ica71108a53bfcfd1892b4d03ef68110c + I177be24718c59688752097fe2a4085c4;
            Ib3a2b744d8f38671a63da6f8f8f1a6a1    = I36cd8882960099f242551ff3cbf8e4bd;

            Iadf1875c584adc34f7586a146184a763= Ica71108a53bfcfd1892b4d03ef68110c + I5971253546899e9a82f387d5eabcc7b3;
            I87716ad5a64592abb812ffe041ccc163    = I3ac47b1ac8e31b0082c7acfab65e222c;

            I02d3f9982f02ea85f996bf5b5975b930= Ica71108a53bfcfd1892b4d03ef68110c + Ic75b8bbb1b80001ec188a0cd25623420;
            I71b259faefbea7ce8f47e0ffb556a0be    = I2a4914c71690073767e6f5fe13f26178;

            Ia6e1b39d83ddce053518c5ae9a5ca33e= Ica71108a53bfcfd1892b4d03ef68110c + Idb0a98cea3ee6cd4308bfc2414a003e1;
            I2161b2ff3514dbdbb79d25da87eeec2b    = I99903b3dad6af712c1148c2f43194da0;

            I3308663053f4307d43ac66f43266f706= Ica71108a53bfcfd1892b4d03ef68110c + Ibe502ebbb366f54a8f8fda4e361308e3;
            I860a3c9fca8d240c68ce3825192353b0    = Icccc370bf2f48ce93f479d13fa7075e9;

            I87ad25dff6c0c9ac46b7a129cb575537= Ica71108a53bfcfd1892b4d03ef68110c + I00ff1331b1900bb031ee81d2a58c1bd5;
            Ie4eb18c7e906c9a25c12e9980a9f61cb    = I5b5a0ccc2f5f9a7554d6d55b0dc61d76;

            Ibf5d40b7c46b50866f58f6fa23e1861b= Ica71108a53bfcfd1892b4d03ef68110c + I9ea09f27ce4484f2e7fc3a6b6d6ecb7c;
            I20a24846a74af76fa4470d6350546a9a    = I0cd3d6b7cb85a87bfbebc1982c5fddf7;

            I0e3a9a3b38875156d15f697adaf95410= I7c97629ec6e594f9b2160815ddd133cc + Ide0abde3644a4fafb436aa59768d016e;
            I90d40f6e9721a7d075512b8b81907453    = I38a9b558c3289d954fe0de802b473be4;

            Ie3f87d094e71e4a82f60e8d91cdd768b= I7c97629ec6e594f9b2160815ddd133cc + I9858bb2a3cc458aca5bf7eb077ee55dd;
            Ifc4525a25f38affb399004b057d1318c    = Iacadd2fc2b7446edd7c45341a0670cb7;

            I793f52d174cd09fe000e8d0351753592= I7c97629ec6e594f9b2160815ddd133cc + I98bbe3b75958f10195dee6460cf2aca6;
            Icc93649a2050b9ded1e625be936b411f    = I316810ae743e5626556ad8f3176849bc;

            I89ea3da7db40e7e6705020462b2d1df1= I7c97629ec6e594f9b2160815ddd133cc + I491f2373b2df19a4c22e1787ef034179;
            Ibcc30c960ae0f29c4efb1266c9e490ac    = Ib9d5224a4d0b87aeb65cd6cf030ee52e;

            Ib2af2f1a928dd824f25b99f0b602753f= I7c97629ec6e594f9b2160815ddd133cc + I9e45e3d7117ce48cdbfc5db8c0ccfcf4;
            I3b2ffa79fd2227a24c6468a89f2bd989    = I92246b941db36e725ce7cbb1c9b4a0b5;

            Ie3e887f5f1a64c37a10404d636212b45= I7c97629ec6e594f9b2160815ddd133cc + Ibadcb205c7e9a0f3345cac7eb41b5985;
            Ib489a11dfdd8a2b3ad561c965b3d7d2a    = I62b8229b8e21a4bfd043c23450ff50e5;

            I5c6a004278f155d33d0cc1b576c3b25f= I7c97629ec6e594f9b2160815ddd133cc + I31b0f2fe98cfddbc05dbd14be8be394b;
            Ifa51cf9f9d3d1b91c72387f5daf05c79    = I49266ae645036370bba4d99a1a85bc6f;

            I6a03a4a548a0906d1a3e9ce47f3454c6= I7c97629ec6e594f9b2160815ddd133cc + I8b611f7c12ddd81de403ba74e212857f;
            Ifda20d77c574c8f13816620c56fff950    = I242c35248366a124753da854841595a7;

            I542e525074d049197ac3904e6102f0bd= I7c97629ec6e594f9b2160815ddd133cc + I004c98da87996b77b5761d366210f782;
            I03ce0915d3a170429959221b6c8cd16c    = I347dd57356eb6e025dada067d0f661b9;

            Ie0307a43ce71ba73d4c8e5ad556bd341= I7c97629ec6e594f9b2160815ddd133cc + I645ff0d8c0a87ba7f792fc83f342b958;
            I9c2da511df8277b7e61cf8611d04dd32    = I6bb3031e93da171fac995de3e23c8b71;

            Ib03e1d3a1f27721e4ea32629c2e86f85= I4823c8239ace86dc399e906c1b5a0d74 + If91268e2b84df18785cd6a53e53eb4e9;
            Ib8c628f3d97ffdf8a8b5db0fe90bbfa8    = I88cede4b89eb0f3917530d0ce2468c3a;

            I782f4ab4666c9f550a2cfc943cedbe77= I4823c8239ace86dc399e906c1b5a0d74 + Ia349e1f7c10a63ddccb3f300c73b4572;
            I42e0e42ae26723497a1da5e86e855499    = I3a590077bea5f1023ac006b321083554;

            Ib991e16161d5c8b3b655e3c7c08b93c4= I4823c8239ace86dc399e906c1b5a0d74 + I977864efb0d94149cce7dc4d165f11de;
            Id7e44a94fcaa2ca22ac9eb6756ecb830    = I2bac571cd0d32e8a1bd527245a76f11b;

            I72f8c6bad4bff3b00055aa8824479931= I4823c8239ace86dc399e906c1b5a0d74 + I5f3ff7fa8686f7a380302d71b88cfb4b;
            Ie91db5e628b828dfaa8c1bd7d614d986    = Ic1c911bc20d03275c7d20ab993e9a54d;

            I58e5100cc1e9b809e93125fe5d08a9d8= I10ad572ca72c2ea991487c39f7eabd7b + I9570f8498d95bee230bb3c5e720bb857;
            I683ebfd7677d9e175d7a86479a5b42c6    = Iff207077a60c0196ac33f68e37d7d824;

            I0aa7056fdacd6022f328a3be49048856= I10ad572ca72c2ea991487c39f7eabd7b + I08581dc8d42be712cfb36d744f2786e0;
            I11090ba16ce17a70438618b474837c33    = I0980811a7928bd72e415daf24b41137f;

            Ia2f40b5c49a2284fb6a234bf7472130f= I10ad572ca72c2ea991487c39f7eabd7b + Ieb664ac9be65fba2e25960141f7fb4b6;
            I845dd61995152e9d39cea7f0370b5a4d    = Ie5a8e0e3d35d27fbb680552444f2ae65;

            I8da184aee7953890f2c89e40744402f4= I10ad572ca72c2ea991487c39f7eabd7b + Ic01904f7c518990eff2dc1de127676c4;
            Ia3e4dff8c98b38b6aebec9094ed26421    = I91e4dd08f282857ab4c275bb1441c9d7;

            I613ccfc7dad5627cde02fa1720244d01= Ie9f3fd3a6d16316e55addbe0e336519f + I9b919f3d4ee3f33506b87bcdaf2d43a3;
            Id69a54dc4854348a482f052c64a736ca    = Iea26a1265fd6c48c038993b2038d2747;

            I080fc6c99e506e569b97433f3fdc3e60= Ie9f3fd3a6d16316e55addbe0e336519f + Id09b8242c22851fb960d55222fe733d4;
            I0f56c52253603ac01a22f3b942429262    = I7920256f397f35450287256339769d4b;

            I79aa118ef8ac0d9b13723fb1f5a7e4ad= Ie9f3fd3a6d16316e55addbe0e336519f + I6d2dbb953a58b91dafa7f0d34d41bdc3;
            I718f82404f82fe0e822ee20d33ad20a2    = Ibad06757b56b14755f0e50620a53dc6c;

            I7e6e7601245ca5b3a58b91848e25a6d3= Ie9f3fd3a6d16316e55addbe0e336519f + I43f2ddd9780f86af489f8deae51168ec;
            I6c86073aaa32b64a43d06eb1a2d9fba8    = Id76592cbf9ad537e9cab20469c5e5861;

            I2792edda66743635b837aa3bec0c58b9= I07965bca84276dd56da1af98e64b0adc + Iebf28886bd39c2540c90e808a9c20d3d;
            Ie0c8e27167e6ba97a83dd238086f45e6    = Ibc80d98586cca13a6849ae053b68e5fb;

            I085cc29465c945957d00cbcf804e3ae4= I07965bca84276dd56da1af98e64b0adc + I954dd66f60316803a8f13a39c460a39a;
            I6bb5e8ee16a2bc0c3b77c882cfb659e7    = I257237e7bef8b0e4cb27bc9a3a93aba6;

            I74a8e879666bb216a331fd2ab723e37c= I07965bca84276dd56da1af98e64b0adc + I1fb13d7500f5ac3821c424bd3688cf4e;
            Ieef625ad664ddadc849be46d1c083748    = I1980cdd5ecb000134e55f507f369af66;

            I7a90a43ed71e82862457d9fa40bd005c= I07965bca84276dd56da1af98e64b0adc + I0a013fff6c792363bd7feb03d9691db8;
            Ice91b069200a91b2ad48fbf87bb2e766    = Id0efde1d7f80f8848613c26fa4637c37;

            Ie1e7b4bd6201baa02b8d59cb0f6ffb8e= Ic2ade31b8bcf68c4dcc1a371ff14074b + Ia072f1d679429d3c3180f8eb67fc7dd7;
            I9d4c7c85b4da5f7003ff05ed3a240a2e    = I76952d4ed281844c1c1795290b1ddc05;

            Ib7b7cdc22b22f276b1c021abaa8fb443= Ic2ade31b8bcf68c4dcc1a371ff14074b + I37b3988d699a1ed42923e3fd1584ecc0;
            Ia8f1616f8a65025446a5ab4cc1624f9b    = I7fa89ba905b099ebafe001878c4f0bed;

            Ib58e33f31be36b28997ba05ef1004573= Ic2ade31b8bcf68c4dcc1a371ff14074b + I7e66a42eb7cdb820cd1297c39f0625e8;
            I29848deb21ad480cdf155d849dc7bd48    = Icd841b02588f755a3133b72f8c625897;

            Ibec394e82f499e8d2d5a9524f943d6ac= Ic2ade31b8bcf68c4dcc1a371ff14074b + I79e3e49f57d47231c0fe6aaafdbc57f1;
            I1ae69988f89b200bd0e48f640211321c    = I52945b9d986280c3dab4248e69247005;

            Ie06ad127e475dc131859992bb5f350a0= Ic2ade31b8bcf68c4dcc1a371ff14074b + I9362b615a612599239e3b752a9334e8c;
            I7ddcc3c9f4d21aacc07d8eb285dee83e    = Ia0319e76fc112b3457f20662a7a51603;

            Ic494a58468b6a7dda76923a9475bf173= Ic2ade31b8bcf68c4dcc1a371ff14074b + I7cf8401bf6893eab0b9f33a0f91ddd05;
            I28f7cf50ea7ac81667ff1353e0e121bd    = I7a82bbf1146a3c68f01abf488a2e3c8f;

            Ib82a2db86d03fe8538fa19d06e501dae= Ic0edcf240048fbfde4e938c3e4c5e281 + I55c425102db0a6838012a165c0597680;
            I09b7dd699ae0c4d34a7d1588efc90452    = I05b26dca2316a9d527da24deb63c4756;

            I5b64727fee9d0825a4ea83261992e489= Ic0edcf240048fbfde4e938c3e4c5e281 + I50c4e1d3a3f63b93bc36b5141226fb3c;
            Ic937101cc53e67403e56ac85011aa9ba    = I256d84c23de18bd9a03cb41c0e3e4b8e;

            Ice7e502b9c2b797719448fde8376087a= Ic0edcf240048fbfde4e938c3e4c5e281 + Ief96603d41b4f670d2bbfa3d3875c903;
            Ib42b03d2f76b8939ff3183008b17a969    = I619aafd5767c45229765838152161b71;

            I792b4f73ed7139b8761443cbc0833e39= Ic0edcf240048fbfde4e938c3e4c5e281 + Idc7df6877bdb7e7d392307d78183d31c;
            I4b99f00b1c2cdcee6bf4f1d2e8199ee4    = I4bbb9f6eb1d79d41c7b5d61df854bd16;

            I278d57d1964cbf3339db450926ef4782= Ic0edcf240048fbfde4e938c3e4c5e281 + I66071f20991b414140869a2e3b750471;
            I01e153b020e1349eb66b47de581408df    = I997c88ff27fe957ec35a2b7146dd56f0;

            I9c1a08b61782ef6c72545504693ac54e= Ic0edcf240048fbfde4e938c3e4c5e281 + Ic7ccbeaf4ab94d0660eb7a0533723e24;
            I8ca1a48206ed8f1dc7ca57d77d0331a2    = Ide7fdb7a17f3d99a7840a648e0873bec;

            I363594fb91d01abca7a2b7402e352fd0= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + Ib3be128b6704cc04c61e0fc9814dcf20;
            I40e8430f50206db37e500c22f461b0c7    = I93dc025ca2d2cc3002c62c5d2e13d45b;

            Idd284c75a230f4b97d5acb98a8e38b2d= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + I29fb3830a5fc5922f1ec687a38941e97;
            I521128b7d945e025ded04037494c850a    = I9c656300bb176deba4be8400371f0ef2;

            If040df53a6410b263f5b3dc3090631c4= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + I511a55c2f4d6d3727dff5825597f55a9;
            Ic24dbb1a30bb9a32c1992afcba90d4fb    = I141a53fdaada1994dc38d694fd03b5e3;

            I31df60ffcaea9cee63b920478cb058f1= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + I762b2abb876381eff6de97cef0798405;
            I06cc903106b42e397fa7c4bc6c5edea4    = I1d81174ecfb84b8c906126d13900178e;

            Icdd2f6ce69b389fbf712e45bdc0a0257= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + Ib393146d81d3cf031466543311cee2ad;
            I765dff22de01d419a6626919d23850f2    = I92ab5c30a7bfae4e698a74d2e48cde1a;

            I8971b250393b397b94db38b9fd0fe501= I8b42e89ff5f780d4ef8cd1cd5c99ef61 + I08043393cb7f2558c145a698ea6652c9;
            Ie9538b63a057a50371de2d17898d3ad7    = Ifd41e7ed8ef5fa870c1abf043b5d5f2d;

            I9199e5e8fdc0e2c62ad1d62fc4d873cb= I70b1b8521b36920707e95fc9418eb8a9 + I8d4f3e64c8e3b0710a4a6b30d27c8be8;
            If93a5596528db9017b8783fa0cf1dbc2    = I983825ee77db3cbd86c937e5fe4707fd;

            I6e03f71fdf20db836c5772658a050e9c= I70b1b8521b36920707e95fc9418eb8a9 + Ie355fa27abbc41291eaf08f2cf9a6ff7;
            I68016caaf170fbe2734c5b6aaf089894    = I715efc0ca41f678f8c582aaa3f255767;

            I2ef49f893dbc8581725ca0f6d1c3305c= I70b1b8521b36920707e95fc9418eb8a9 + I6fb63ea54e492bdbc6d1145affc683e9;
            I169b0fac6d01a713986b636bf8dfc3fb    = I764815deb8bceeb1b9929de2dfd46235;

            I8796f168c892ac60c38a0a7f1e18035e= I70b1b8521b36920707e95fc9418eb8a9 + I1898bc3cc6a8b6f71d65c758d1f08366;
            Iddb14d68b464d04fe9e0b4e62789601a    = I1b869d6b94307bc9bea28db11161e61e;

            I64a26e5117c8f3ab95bf0dfa97427243= I70b1b8521b36920707e95fc9418eb8a9 + I2aabda12ff89e708d04b4399472b5203;
            Ie5b71f77beb734a6ab7f7be6c6f9c252    = Idf695c6735d8d8aafa37ad4cbd5a5872;

            Id7946a0299ced3ba00f6c3e6e664931f= I70b1b8521b36920707e95fc9418eb8a9 + I84865c4f872c0845124b78fabf695c2c;
            I59f9fa0b81ca88915c338ece1d1e08d5    = Ib9114ddde15c1908595081b52ba00c48;

            I5243b90640ea4680de83021601c85c39= I4fb1c32a62cbbaeb585c6564a3c938f9 + I91a8168d3b087ab3891cd6d479427b95;
            I4f27922ccb21b65dcfe2dc0fcc97cdf3    = I3d52a609547a0ac3cd6d0481f09d00f2;

            Ic8301fceed328cc031640ecc4ff34803= I4fb1c32a62cbbaeb585c6564a3c938f9 + I2493237a24acdcab8b5bda10e804a5cf;
            Idd7ae55ba748fb36e49684037212936d    = I45abcbcdc3951ebaef039e6cb2562d4d;

            I6e852c94b6105af62ee85f8adf77fa55= I4fb1c32a62cbbaeb585c6564a3c938f9 + Ib3e7633767b6e09e4ee54f6feaddd31e;
            Ib8da505d1572487e814e7b0682e6dfa9    = I5bed8ad020614972a82bf3ad66300f12;

            I7d98c5c2a54832b6368ce60009208eb0= I4fb1c32a62cbbaeb585c6564a3c938f9 + I896cd566a3d078b0f697a788efd223f2;
            Idedb59a6fa2f6ad049f81ac652c645d8    = Ic7ec84d03001998a8504a79afb1f0d5c;

            I7e42f2281518bead81a6d18d2dcbd1a3= I4fb1c32a62cbbaeb585c6564a3c938f9 + I8c733a5d394e6b8d045eede5cc7451f6;
            I7d50b49718ab2007accda67ac77a65d0    = I43cfed51e8dec917304dff4f44a984c6;

            I63c126c978154f2d68b11f08a938dcb4= I4fb1c32a62cbbaeb585c6564a3c938f9 + I57b9dd7a7deea6695dcd03439c9723cf;
            I27e0600689451a7475a36143f0eb1079    = If34baa3a92291d91308582e9c268ccaf;

            I2ff7719c35578b47720cacd9ddfd92eb= Iefc37daeec14e14ef2fe0716f73109dc + Ic970a88c435a85d21ed71c6060b8a8e4;
            Iba6724b61ecb74552b9bb3cab96480c6    = I8c00e1f1c7faa04600505a6f30e32ccc;

            I480599aef36967a670155dd77120a37d= Iefc37daeec14e14ef2fe0716f73109dc + If83ce1cbe3a73472419520c225b288a6;
            I0abb44bd896fbc695e880fee67fb0c42    = I225a03b34b73fee071973985a66f9213;

            Ic000b2c844de484b8f30b7b84dd6234d= Iefc37daeec14e14ef2fe0716f73109dc + If86532f849bd392dbf599eeb2fae0545;
            Ifd714548110aa979e735cc6e13d3ef57    = I4b819b7da7ced2a32e77b3b26682168f;

            If0e25df151db991185f992eab5d5be99= Iefc37daeec14e14ef2fe0716f73109dc + I85a7fede715578be0634d71e9c7951cd;
            Ieeb6c7cdf1379ee3d2933d81bc812dbc    = I3d1050efa384172a3af1fa5f259a3877;

            I2f533699abb7a997160bf4ee4cda3efb= Iefc37daeec14e14ef2fe0716f73109dc + I5d4fb4b5a5ad3dc48beebfa0e0cebbed;
            Id682af5250edce8e3811d418ecf2dd10    = I66de52bc354a661ccda6f4d6d744bfdf;

            If6b33cfc6d34e33fbb18e08fb4d8a5ed= Iefc37daeec14e14ef2fe0716f73109dc + I1cd6b35bcdfd461db69a4c1bdb1d387f;
            I1d02127e28fb2e9aaf352815627960e7    = Ib9a88f5ea722553569167ca7b186fd50;

            I2ea5423dc8726fc0217899e0f406a1e9= Ibd15f164f6d2ac9e5721a21464bc2c5c + If365a3c3ef86dca7c7315b91298c2db8;
            Ibee34260749dc92b8523e83cd64d6a40    = I68904155ce7e8d722b67725f81af7f06;

            Ibf3f4f8a04cbacc9624ca5cc73bf7069= Ibd15f164f6d2ac9e5721a21464bc2c5c + If2021f0735c6c5649ebac0d230fda87c;
            Ie9a2a59c7b3571194198dca0c679c5f6    = I7bc807d9f1b67d68e11c8a064b218963;

            I9ba53c36934ab1c7f498241a79cfbae8= Ibd15f164f6d2ac9e5721a21464bc2c5c + I12c07042202f66db926861c9ce7c2b25;
            Ie4b5a941feb385e88498a98e5f8ddc01    = Id1b5740fd8ce883d3cf724bd7410f27e;

            I106a25f18536f96782927bf3bc2ccd72= Ibd15f164f6d2ac9e5721a21464bc2c5c + Ifce70fefde8f5ea4d2c1857236f66d65;
            I30b2b34a0cecfdbdeecba5f286befccd    = I12c6efa1dbc88f222ebcb8866946eea1;

            Ie5cdad65e918679607cc5f816987b736= Ibd15f164f6d2ac9e5721a21464bc2c5c + Iffeefa89a2ba7d032db5db64cbf05e20;
            I8ce739ddc344cacb2de7f2c88a882170    = I9c9d28abad8610fa2cecb74d18a1c9e3;

            Ica6dc9ded8756fd6f82eec4271e246c3= Ibd15f164f6d2ac9e5721a21464bc2c5c + I40a1ecabded8add5bffe316f2d8beda9;
            I8b00260bb93e928e66e9d4aaeb0d9b55    = I21af49923adfeca8b24188a7bba54b1d;

            Ica42ac6ca5813d0d1a67f14d1248437a= I951dfff9507bb70214d48e03a0ebb3a7 + I16e3f3a6802fd206654bb622fa1393fe;
            I9c1ca916654bad308af37d040b486cf8    = I46c921b6dbb398813ad0d6c06e2eb33a;

            I13dc6cfc75ef846c30e5dc1dc5305d59= I951dfff9507bb70214d48e03a0ebb3a7 + I7a029c27d92754041eb6d605837238dd;
            I05749703a8a131453c563ed2264680a7    = Ifa087dd71378f388142d351fa18806b5;

            I33e784182dfb4af39715788b1ae98af6= I951dfff9507bb70214d48e03a0ebb3a7 + Ib8b95ece5da3877b261a06e6d0571921;
            I4b76fe5f9863a41733b76decf9867d16    = I3f3c345d02438bc96a1f7b162315ea43;

            I9e1a66805348d2e5bbf5e2316187444b= I951dfff9507bb70214d48e03a0ebb3a7 + I84a62a133dbceb5a32a7c907f371663d;
            I2805bb16fd574a64de548b39a532cd8a    = I7577c4409a32ebf50e5a187f71c84b1e;

            Ie9619916a96d218cf5eb5f3a4995d0e7= I951dfff9507bb70214d48e03a0ebb3a7 + I42564ec6a794ea803795f0b5b3523a93;
            Ide6a696c06f17f455d56bb28cad98bd0    = Iec97b82162ff77d0b123feeb5b5904e6;

            I02ce7969c51ad141df227ed7d18e74b1= I951dfff9507bb70214d48e03a0ebb3a7 + I7c52ae4af926267b5e27a530202fcce0;
            I39bce1f71ede4663c187ddfd6501eda1    = I2206f864d477e44a18769ea9cc01d8ee;

            Idd73461af0d75c4d820f7f8f0f419e0f= Ie78e30b2a2eda75d0df7d10fd67b5e36 + If79bc5a35cb55036a367efb88c7d5510;
            Id0e769bee61ae0a90c167fab061f5965    = I9b67c7138cc6e8c9ef36b5cb28932c9e;

            I3df6c2cdccb2a82c58c1d81b00af7786= Ie78e30b2a2eda75d0df7d10fd67b5e36 + I00dad36628d2fa923120fdaa79bf0045;
            I83e03af8657a4a237641a9da7922e502    = Ic295c2717dcc256113776b8d39368802;

            I97f441fc5ffb88efeb5ed66b60f07a7c= Ie78e30b2a2eda75d0df7d10fd67b5e36 + Ic99654bf4833c9132912eeb4c0dc92fa;
            I7565e071282ca6e77bb469afc522f1a2    = I4875abaa409c919efee2cde0c90e1e7d;

            I3194a235eb652c8d0e4307cd056e5e72= Ie78e30b2a2eda75d0df7d10fd67b5e36 + Ifb9b29c43f435452cc761218c509f5df;
            I5d0dc5d40385ab67bc7f540f212b6a97    = I0bcc0953acf369ba9571d11e68511af4;

            Ibc315f6c79ba2bf336ee57f2e5f7d776= Ie78e30b2a2eda75d0df7d10fd67b5e36 + I514830acdad20c4ff3d078477e939b4b;
            I548cac395730b8386670cc4c7a64319a    = I4d92612c245b6ebb246d2f41b3dd4107;

            I937a54f5cda99a7079c7fa46b4ea26f6= Ie78e30b2a2eda75d0df7d10fd67b5e36 + I1a5c6c50817db8bde279d5f0b5095d76;
            Ic6d9bbbfb7890540edd10aa5758b0c4b    = I53a8be01a8f8067f67e0498c48cfa2a8;

            I49c99afecc613656cd1469d8c1e98936= Ia0b83a372dd4115dc4d61eb8ff0811b9 + I12334038c2be8634c47869f397503019;
            I7beb1f915a881a302f93c869d81417d1    = I036d8ab76c1f8c3b52ddcad50c6c8a6c;

            Id76ce0333f43bf7bccf1ce48e25ca69c= Ia0b83a372dd4115dc4d61eb8ff0811b9 + I03829256e357ac17c7ca7cae2f980f41;
            I5fc389bbc1ce31f7b326da719dc576d4    = Idaffa51af26a79990b50e9422da6074c;

            I2c77f9644145219005751f7a4eb71aaa= Ia0b83a372dd4115dc4d61eb8ff0811b9 + I3f193e9c265c1dfaeada63d59db5b79f;
            I922e6f05f7c6e0f6f0b1a5c9548df238    = Ia17748dd92434f8658e49a3f7ed682e8;

            I5cecc266272eef88cda88c1df9bcc37e= Ia0b83a372dd4115dc4d61eb8ff0811b9 + I9ab3cea6ee8d8473221da21bae06066b;
            I8c6bb234a1ca3deba637adf746672194    = I1ecdfded32659bd57c752928f0cc12eb;

            I776a0b1b5c14afa21b7fda3c2cacafed= Ia0b83a372dd4115dc4d61eb8ff0811b9 + Icf8cfc800f0a2aa5140a7f83f035b0cc;
            Ide24ebd7423d4c4f43577b019f2e30e4    = If7bcd20651da485996362af6b633fec3;

            I84860b1f933339e0f90beeb3d666393b= Ia0b83a372dd4115dc4d61eb8ff0811b9 + Idf0c1b85712fcbbbcc12915158ebff62;
            Ifc412122eab7560c9021a17d7f8700c4    = I7a04a2c4768a6703cb98c2adfd53088f;

            Id24581713f1ecb767db39d5154c2f5f4= If5c5bcbbea01aa22f242b913f0d01929 + I715d59fb27e519a9b76bdd8b5139a619;
            Ia5a56ed2c6b98e72002c6c5f946e7264    = Iebc9456956b29940df3df4dddae0619f;

            Idb0eae2f0e1dae1d56251d64e2c51f9f= If5c5bcbbea01aa22f242b913f0d01929 + Id1df78ab32daf524b77c0431c782f2bf;
            Ia888ed8885f66084b777f66e25cef1e7    = Iefb9092502c1c93656c9050bf74e6849;

            I2e3ca4b130e6d3d92385928a28644452= If5c5bcbbea01aa22f242b913f0d01929 + Ia344734d285ac29b53cf401c08a0f987;
            I248229aecef00b87a70ce88920e407f5    = I42edf14a24cb1e19924e0f5531f97ed9;

            I7922d80ae333dcfafde31d294f0eb4d8= If5c5bcbbea01aa22f242b913f0d01929 + I4a0033a180d7edce81fcfef603532e28;
            I3d162a0ec918f220a7d5f4efdf89cb58    = Ia332b7b61c57cee58ef4a1733da2afc6;

            I82de04cd2dfef5616efca4af26d7c561= If5c5bcbbea01aa22f242b913f0d01929 + If0b9225e759438be175c4128c78605ea;
            I1ca0372f60e48f2f803778c9017023c0    = Ib4450f5e900229ff87baede34be883b4;

            I7ce384520525b15d24c2ef6f161213a5= If5c5bcbbea01aa22f242b913f0d01929 + I6b32298e8c61e75d0a38bca3084c0528;
            Ieb9693d54f0808b0ba463fd3c316a80e    = Ie7d8f527db720e17a73a57400a5360a5;

            I56aeea71c7bd19d47620cf36adf3f115= Iccba58cd3519fb4cc75a61b50da1d562 + I566224393f6bb27bfd8b0b0d6b8e53d6;
            I63da03315d7e51fcacb0bc0298e506ed    = I7c420e9724fd4bc31071a57ac1ba5293;

            I138e1a6db0c6649bc023cc36d81d5b47= Iccba58cd3519fb4cc75a61b50da1d562 + Ie1bf5d97b8f679095d2442bbf9f95608;
            I918f5a12e96bb96941f019940f27a5be    = I5a38174a83eaebe2678ca70fe5915c02;

            Ib5e8b1c4dd9b5dad56b59cc11c87a258= Iccba58cd3519fb4cc75a61b50da1d562 + I9d0fdb45b9e86bd409740e538a690320;
            Ib4fb115f442ff544fa3d21b4e9d3f075    = Ib3639c700fe97648415fd4dfc8a6466b;

            I86f785e2d5e8d6c08fad1d334c7d244e= Iccba58cd3519fb4cc75a61b50da1d562 + I4f45dd50d2825ab338b8a2a8264096c0;
            I387403482432a3196109484d1120d584    = I5228b59565a0ae5f56237e5332ddefa1;

            I9a6c8efca218c724da4ee4c1087d58bc= Iccba58cd3519fb4cc75a61b50da1d562 + Ica94017f26e96fb22a47add326ee126e;
            I619af17eaa4a56726d6ab322a74dd0a4    = I87188c070d52012c107a5b37e718a5d4;

            Ia30e8dbc6974ea94b763842e8dffa633= Iccba58cd3519fb4cc75a61b50da1d562 + I5b0d72cedc120406402076148e2d30b0;
            I7a67ed3bb370520d0d25ce407ab8cd8b    = I7d0ebb3f7a7e77362b41f9ec9b98c9af;

            Ifa60f45f4d8848eb0b89f5644ec69668= Ibc0999e4d0b3cc2650f9348b8c204b14 + I4b5713aee09999592256c407d4b8a95a;
            I7629b35ca548190a81021a2c13d8919b    = I1c2e01ba53fb12e4c3e44e4a9ef97888;

            I0aeb4b93cfa6d62ec41b7e6dd0287dd0= Ibc0999e4d0b3cc2650f9348b8c204b14 + I64692d5168554dfd7ce1c7a046aecf72;
            I004851d3828f135ebe4d2e6ab83936bf    = Icf7e609c4a537e6f2a7b86b7035717d3;

            Ifce1fc978fb5b0187593f46f53c3b469= Ibc0999e4d0b3cc2650f9348b8c204b14 + Iea71417e738c6ca54c50aa014cc38627;
            I0e2c382b2e62ed43b76697230e34b719    = I39d74e21fb67539c0d310571b99a3e22;

            If3b6de7c919c5d53a0e191a75bd7e574= Ibc0999e4d0b3cc2650f9348b8c204b14 + Iaf624549f73b0d13c1a73c850b99f810;
            I36dac27d10701db70fb2b5996a3f038f    = I395b85e88acd203dd93e519710aea79b;

            Iecce594e6e99b0c05fc845144a664b07= I2aeff1fb4b839a581acaf26f90f9113c + Id1dce8c1542f1279badb381aca3c9b51;
            I51d62ebd160eb0d073a7efb64d20079a    = I850e5fd50416aaad26283152c4a49ddc;

            I2c8431500ecb25619d2884a2fb4260c0= I2aeff1fb4b839a581acaf26f90f9113c + Ibe6a876a041198a581c95457a7d1fcf8;
            Ib3545a88d68631af1c94ca2cb1f379af    = Ide38f5cac19b1bc82b26bfa12e5f9d8c;

            I217c710f7ef39035546efcbb043f63f3= I2aeff1fb4b839a581acaf26f90f9113c + I57db98eb439d59a895dabe029c6a3a8b;
            I81ad7b044118734f4dc32a1a4e8eba31    = Ib2d8874232a27b78a8c664e0fa2af512;

            I1b4236130cb1879d885653fdd9eeab4e= I2aeff1fb4b839a581acaf26f90f9113c + Iaaf7efeae9f6dc9e8222dc2b10122000;
            I5ad8c235d46349b6d310d0f175f84288    = Id002a482b2a09d2d17b9fa903882e8e0;

            Iae0f7c13f1564d63b4bfdc152ddf4111= I7d60d53f883f8187700c4e78b4c22f1c + Iec8dc328edd6cbaa2d697e05ed222746;
            Ibc00920378e2427df2a63a47dc3eaded    = I359451948e89283ee89d89cebf689445;

            I010592496030d138a3a4245d00069957= I7d60d53f883f8187700c4e78b4c22f1c + I8fcad6e7d5ffc9f79eaaf634f6fe8cda;
            Ic5195bbaa69d95059cca6e152dc9f705    = Ifffc8f779e22eedf06f7d1c24da411cb;

            I9d7f47a6289a16448221d61f301586aa= I7d60d53f883f8187700c4e78b4c22f1c + Ica26f542586d50c56ce0f3c00f36b388;
            Ia01f20e0bcf35c2ee4963e9c392c1004    = I3ccf7fbf7a13aef5daa7905b485d6e3a;

            I7b8ed2953170c4deadaeb33a6ba165d4= I7d60d53f883f8187700c4e78b4c22f1c + Iea1cd2321d2ac9b891b344e2ba2363d3;
            I9f6f48fea88d1cd73ef2b24c7e819964    = I9deead4d27ef61f468a1bac90adfa27e;

            I4efe9eef6a48aeb0a9ba4e0ffd9906c3= Id6fcf4b7af4a37c854a12e2ae80851fa + I83560e8d0f8cd37815cca6336fb2208d;
            I847feea780cc8a06caea2d2ea79ad281    = I6c050a19b5031493dcc7163509b00012;

            I5a8466bbd83c39dfbeaa6399e3fb3337= Id6fcf4b7af4a37c854a12e2ae80851fa + Ideab06dc2448a6950cd1a06a0c90c2c6;
            I7ef6f4aeda7fd6775839c068c681f9bc    = If74b57fb1d88f063bfef26ae6b74ff2d;

            I1ab96ffa948dd09bcc4f748c6c2575d2= Id6fcf4b7af4a37c854a12e2ae80851fa + Ic5ca74b66763c6e5591c7c2bfeeb0663;
            I0645e741da20a4957747188273a655b1    = I9fc7952b3920da1adf39777e9a1cd13f;

            I016f57568eaf00b26f8a22100858c158= Id6fcf4b7af4a37c854a12e2ae80851fa + Ia544fa24b953fe91800978895e3e610e;
            I71125dffdd2d37e44dbb46143c1e8d9a    = Ic013de8383ced83cb6cb368e54cd0f43;

            I1fb995e302f4f1ba493ff85f39938175= Ifa5e5f7d753964f14f0f16dbe552fd85 + Iec078a95a69b081cfb5e987ba9c5a613;
            I50c166f958b22ce866cd40334918274c    = If71eac564bbca0cf2967a8803a24f586;

            Ie643ad235307c60f1ee96dfdcbc8c2a8= Ifa5e5f7d753964f14f0f16dbe552fd85 + Ia71663e8f563041c27cd21a0c9c27a28;
            Icd225144fd331b870847044b4d02bed0    = Ib19bf2920a5486af62d38fa181293a47;

            I8dafdf2c780082d8dfc2961b3447f104= Ifa5e5f7d753964f14f0f16dbe552fd85 + Idcef10a0465614cf38e0d6f503b5174a;
            I5e876482090ce6007c2a2f2101c24654    = I92a94b468b025e5c1d103b2f8c92709e;

            I3a2841a0f5e1b42556f384231ab0717b= Ifa5e5f7d753964f14f0f16dbe552fd85 + If2143db72bf9a02b64eb45b3a4faa39d;
            I026ded06f56d9ca93f47fd85aec4f7ad    = I76fe38786c53eb9f57d6512adb920d5b;

            I2b00d0e6facf01274c0c3446bb0e1599= Ifa5e5f7d753964f14f0f16dbe552fd85 + I7fa710c37f5f96c3cdc35612a702a71c;
            Iec596e94ec168a564bccbbaa7df833c9    = I7878eb8ad885ea4193b8534015a445bb;

            I2c645d25871b70dae5b2c283695d5130= I900d471b087cf5a436c2ad66a84d8280 + I6f0f74dcc830fdcb0af9df75a2b722f7;
            Ib514e01c261e43a725582a10596eed32    = I5b26270d07cd79afa7019dac72898e3c;

            I540a0e8968a6a82aca775a81ef82b520= I900d471b087cf5a436c2ad66a84d8280 + I0b557cf102da41afd26936cbdb64b6e8;
            Ic19a62cdecb2329370f7e11c48d3738d    = I167dccb5e632afc0686602b35f9dea42;

            I5b95bbc82e6d8d87421efe3f17b97ea5= I900d471b087cf5a436c2ad66a84d8280 + If65eb5e743a7b1878fb232ef2fe13cb0;
            Ib2f5691baa59adfbaad62f6ffc71fb05    = I3cb81e29fa5d50fadebe311acca6d090;

            Iad81f5e5e728ffdec6296b2aff668d75= I900d471b087cf5a436c2ad66a84d8280 + I3403ce6e697b523a9f441d8fd5e2d420;
            I9bdfaca6112385deb86e24ad7e45bbaa    = Ia25c11794a51c0937e0600032133a6dd;

            I960a618f63372da74581b8c352f3e618= I900d471b087cf5a436c2ad66a84d8280 + I98fd105696fca11c1075f9bd30013747;
            I0e647bb8351cfe7828423e7099525585    = I95b38f00928726b7b701405baf74f66a;

            I4f5325f1601acde10018d1fd0aff4d35= I6d1434907f0292ea2ee47cbc5b52bfb9 + I1d7d7a68fc53b8be89c4637ac8f29380;
            I185b758fb3e50bcfb1464fe2ab593cfe    = I32c90cfef12eece5e90200ef79c7231f;

            Ib297101fe456520e72cd9d208af44eea= I6d1434907f0292ea2ee47cbc5b52bfb9 + I3353a7916b569f2c0ca122180608dccc;
            Ie25e944f9e3100c39b69bb38dffca177    = I0b27fcbbc4514fa212fe3d023bdb526c;

            I73a21342321a9d81a0fa5308149d72b0= I6d1434907f0292ea2ee47cbc5b52bfb9 + Ia457938da4efe847cb06f645f2a54a52;
            I8e77032a54376578b3d16799e30c97f7    = Ic420c6e4d3748dafd05197706f316f62;

            I2a486524f4f53b3454ee02a8892d4fa3= I6d1434907f0292ea2ee47cbc5b52bfb9 + Ic7a21921e2716fba55aad2e351f4498a;
            I4cd2a7f8f8ec378200b00d03e447ac92    = Ifd760e2ecefe198d6f583146e8cbe9fc;

            Ic6c4e4e6a9ba43a3354f9f3192ab069e= I6d1434907f0292ea2ee47cbc5b52bfb9 + I61345963ceabdaa0f25f8a463fc9fe5d;
            I1b3c55aca0da232cf3f81d6d0914729f    = I8078293bd2540592bffc91383fa5ad38;

            Ie3cdee3560bd06aed84dac5fcd2a259a= I938bef7ba7ae1739d8e6a6a7c117a1b1 + Ia4b438844530fff602ea04e72b07db8d;
            I34c76f1a126120c4474e750e9b51e034    = I1c0777b46bd3a7e2126f614d55703204;

            I584febaa4c440fd9353108af36d3a5c6= I938bef7ba7ae1739d8e6a6a7c117a1b1 + Id4788855f9a503e8b506d012aaeea445;
            I0edb624c344787066a2267757052196b    = I2a719cff60bf0985e451a32aa71c82fe;

            I515e78507d7419ca14d77b6d52f75a78= I938bef7ba7ae1739d8e6a6a7c117a1b1 + I7c68e0ae30efc4ca4d68b6047119c6c3;
            Ia8443f199838742595ac114f35c00143    = Ia1af17b99a087b22fecb7ff79a370363;

            Ie9578453a57d2b3b9c3b98844044b5f0= I938bef7ba7ae1739d8e6a6a7c117a1b1 + Ib45caf6b563d22144be3e9225a99a1cd;
            Ib25b8a538c9d64880e114bf4a80ca42e    = Id75247b073a7993bff1992cfe1874ff6;

            I1e58b3062097a46d8d590232b40278cf= I938bef7ba7ae1739d8e6a6a7c117a1b1 + I9e8375af6af10f4bac3e87e416d430ee;
            I25f6a3d7bb869082e4dbbd0ee8574c95    = I63a6ad22f067ea29cf79e51ebc011f8d;

            I3af126eb28c67797ce625b0d82943833= I6384a9416b2d1da01df1b2d7b16c5390 + I8983f003c30a218543f39f5bbcd9a25c;
            If96057023747a1538d9f06966af48bc2    = Ic3b5918c230369180edc94c5b01046e7;

            I130ee1a8acacf4cae8818cd8320d050d= I6384a9416b2d1da01df1b2d7b16c5390 + Ib34ad1d14978608d1440f59998a31672;
            I199e995390462e06853b1f5cdbd46e0a    = Ifdf2c8ac7eb668b49ed3cf950d08c179;

            Idf92dd09c29ce8e921b2b34089550586= I6384a9416b2d1da01df1b2d7b16c5390 + I380ff8528cdba4026fac3c4eda8b2c52;
            Iec6325d585ddd0a9f86bb5cd0229960d    = I644ff86dfecc5a20a1431f9cc67ee6f9;

            Iba74a64cc1d2ec3c83a4061db298ad37= I6384a9416b2d1da01df1b2d7b16c5390 + Ie72268e979cf069b88f6eadde789e5ab;
            I4be1ccfec148a522fbf5b8375245cbb3    = I56a7bd438035251cd67dfb97b3a345d7;

            I01364c233ca541914d790354515aa5c1= I6384a9416b2d1da01df1b2d7b16c5390 + Ida1cd844022bbf1b8431225e66b2b78f;
            I074386ff6a3d8d644f4b2501c69f26c7    = I00c294596fc87af7f1b8377260232832;

            Ic6a8297308a63ed3113008a3cdc76358= I5097a79e7cf7a30d38ba198d1407119c + I16d2084ccfb102c3bafc701872f5ef2d;
            I83b378e5534c553b57beb22c5178a3ce    = I7af09468b60d8e594a1aa85ad74911d5;

            I6c7ee9d0bd684a7f54bed3d52452219d= I5097a79e7cf7a30d38ba198d1407119c + I9574759e112f27778f3645d5d49126b7;
            I14f79d67f75af6a495d6eb2986210cda    = Ic0ed40d42c2af78809ecb381660ef229;

            I985ea87550ec8a222e6af621589e186d= I5097a79e7cf7a30d38ba198d1407119c + Ia8094903aed8dd0ce8e9ff459a5287b0;
            Iacd805413ec1eb001b3083554f187554    = Ie03547bf9963c8a716e20e4aaef52dc7;

            I6836a7d1e006d7f7556edf8b31aea32e= I5097a79e7cf7a30d38ba198d1407119c + I502a8e382aa0881dc86f3c13e0566ca3;
            I3e61e09fcc81a0011a79f5c5ce77bc46    = I26e996666f3436cfa998f34c3a05f7db;

            Ia7a356a18af18ec131b9df46019f3e58= I5097a79e7cf7a30d38ba198d1407119c + I30e9ab592e97dbc5fb6ab58d2ffbf8d4;
            I6e6cbb7dba8eb3c02b5b4e4469e23cea    = Idfc51f66e038c5ae625e98b615a7beaf;

            If3a7e111247232c47ceccb5e05338312= Ib113c26c8dcf49c972c41a938059a787 + I099441ae3d3dffe49b18bc578af54dc7;
            I8b25822c33f7d506ef69216af3fdab44    = Idedf5a83a99278f57c6c9294b66b69eb;

            I5f38d1665294b2d3c18f9cd888ff60f1= Ib113c26c8dcf49c972c41a938059a787 + I0e8f3f56bce3be1ee4d5f780a2f2a9fe;
            I06fd642cbc8aa2f65197801d7459cfa2    = Idf55d61336e413c5aa3226b3b44f27b1;

            I10290b9576bf3d8caf90583a388226b7= Ib113c26c8dcf49c972c41a938059a787 + I218ee96418a4f5d734d3d71685bc09c7;
            I22202e6c3de9b06c04ce9514af28933e    = I05ce5256e568621df7129058c50e9fa6;

            Ief36236305fc1521c5bb4c60753a676a= Ib113c26c8dcf49c972c41a938059a787 + Id5fd6f25dc3df22a322434ae3c90dea6;
            Ib991cdbb91133cb82e154c575e00a174    = Ib8af108fab1636823714995f78c9d575;

            Ibaa0539fbf5ccc979511c09c061cf494= Ib113c26c8dcf49c972c41a938059a787 + I2ec2a6de2be39b1bc259b0be72e35a0f;
            I5590364df6874420e169aa444ab520b9    = I166d54ee9aa9002c59a0aca2834632f5;

            I95664ffd0ff13c2893421032149f24d2= I970c4a25a8bce82a9d2846679029fcab + Ieb1dbb98d5e5bda5b9ce803857f2ca26;
            I43a9e393037fb4aa84741dca22648459    = Ib5f971498046dd212d853ff440c553cc;

            Ie390153b3b7985dc63d65913de215377= I970c4a25a8bce82a9d2846679029fcab + Idd95fd099dd2b53c46d02f09575b8032;
            Ibb4d8301d90c66fdfac92b3fbc53c019    = I325d401c6a1f445dcb7a83d90d2da75e;

            I704147dda658f4a03627dacc1c91dd48= I970c4a25a8bce82a9d2846679029fcab + I1fc36e6f738fab96df356979e1e3a612;
            Ibae217fa4b808e4accbeb8f4a9a976ab    = I91eeb6252974a1f69908b7e7114b95f5;

            Ifb09672d505898f081aa13c95fcb88b5= I970c4a25a8bce82a9d2846679029fcab + I2461055ef9b1aa2ffca0f5cac3300e71;
            Ia8bd7a3594f7084a57e64da023bf784c    = I898cf70b6c6b57d256490f44d257fd84;

            Ibb5cb89097dd11bf292d5b5a2422175b= I970c4a25a8bce82a9d2846679029fcab + Ic32e349efae2ca419e095ee5e15a501d;
            I3ce4b9d41f5472bf60ed2802a2ab10eb    = I256f73600515ae5c410454c425b66696;

            I4a305956b18d6ad6901d2c17e99f2bab= Ibe2af096ad2db26e54d8b4b3bb05175c + Id1b5c33bc63f75561b7cce6fc0981c69;
            I93ec9bc6fbd056e7e52496546493e727    = I362d1818937fd8d777531b85e86b4145;

            Ibf5bb3b9eb1812383db9634fa9a27ad3= Ibe2af096ad2db26e54d8b4b3bb05175c + I2bc3ffbe5b42b0833206437d3863278e;
            I2374b90dde1cf481baa40af31e1a43e3    = I21dda2280e7aa79b6abd7820829583e1;

            I66b37d055c3735f011095ee4b1ad02ed= Ibe2af096ad2db26e54d8b4b3bb05175c + Ice2c390d296e09b117d60905343e9098;
            I0cee595f488a909ade8a3b4c90dbb0c7    = I94a6499c7bd1d40e4f363a58db1aa114;

            I43e71dd694d97217e242f267248cd594= Ibe2af096ad2db26e54d8b4b3bb05175c + I036342f6be0f2e2f1f4927099a5c4a78;
            Iba4c3d91d492b000ab1de7add9f171a9    = Ifb6f3d60109d87ffd54e72b3958c7e80;

            I4baa925db1ec733bd4bd25d9dc873e23= Ibe2af096ad2db26e54d8b4b3bb05175c + I1befb935ee9cb871c9a7476c1fc0da3f;
            I2b4152aa4c51cc1c1ffabac78cea267c    = Ia3fca25225f6cd049ec92b44cdb57049;

            I547928c9db7acc531af251264d576ffb= Ie48569c467fba0c1291f71d6080ebedc + Id680a9affed622577164b3a8380494f5;
            Ie4c3dd5c191aff00a6d62006223c2b76    = Iefa9788b8791b23ea0ca3d756d7e4019;

            Ie4ce634b2fb62a20781f8a2e8fddc762= Ie48569c467fba0c1291f71d6080ebedc + I5732fdb805258fc13c8ba4aaf56574ca;
            Ie4c0ba9510f9b924999bb5f432137271    = I2b790f210029547ce774150b5390eb12;

            I0e90e96ffa64c2874d79110b622994bf= Ie48569c467fba0c1291f71d6080ebedc + Ia2fc8a1bbc3cb0dd7d89a7f05b04909c;
            I5bad544a17b384973d5672acbe0ac0d5    = I5c474a60ee2779b8f1477d07f4ca88d1;

            I767e37e3c6f4224eb07adeda480ce253= Ie48569c467fba0c1291f71d6080ebedc + I6bfbf7ff79ff0a6facc9ba5031239644;
            I231bfb8e19e1d9c4bbd29a0bd75c1ed3    = Ie542464c6c79a43b078a8314c4def3b6;

            I75fcaf2c65b7e63adac834054850c6d6= Ie48569c467fba0c1291f71d6080ebedc + I01c57f697f2af7d2c6ae904319f10725;
            I1ecf87e33de04d02db9e64590bcaffde    = I0ae4560405030e9485f14f6eca025625;

            I5f1de2dfbd79204ab2db9b686d6a6862= I90e7ded06617b49cdb8b5301fe9c6a20 + I58f89947eead94b5054a0fea3520ae33;
            I60c97bf58193f004e3fcfdbd6a03ce6e    = Ic14dfb6df2b9a62e5c9471684c0cb07f;

            I8d01de6be4091dca2589cef625c05229= I90e7ded06617b49cdb8b5301fe9c6a20 + Ic462cebbfc39190b22d20013259e39eb;
            Ib71065a3fe70d3ab5f05b0c393278631    = Ia744719b1036a2236173a80ce326bb7d;

            Ic09e773899fdd208c0fdd874933b2cec= I90e7ded06617b49cdb8b5301fe9c6a20 + I7caa41076a293edf18c7c4309fdcfc91;
            I984074a5c77445ad266463e20d77899e    = Ic3f0e0640b27dd1a3bd39f6b9507c7fe;

            I24a3f9fd851c4af70ef66bfcee44af65= I90e7ded06617b49cdb8b5301fe9c6a20 + I33d941ad9d4858fcfb77f0f6cf99d2ec;
            I50bb40691aa09c42e0b64a076b50a971    = I82fa0db281b140ed781dcf5c53625117;

            Idd31807ecd603db8c719349a2be1be40= I90e7ded06617b49cdb8b5301fe9c6a20 + Id580f8a2748efff9b6b747c497c16e9c;
            I753bff437b6c563f5fddf19685405504    = I5dfa454e544e731a6254e73c97d79e06;

            Iaf680cae40d1adf7649da12b31a2be0d= I4920014f5d017f4e840dc3b88526955f + Ife1c8d014675240a94f1133a78703ed5;
            I21f2ec69bcc507756e2a5f85d3ead3e8    = I3a57ff68cdc9b93c07bc79f8cea77473;

            I22d948171c1a66f7a28d5e51007700ea= I4920014f5d017f4e840dc3b88526955f + Id812a8ea2a3b4a912d151be582833fcf;
            Iddec4486996054e475499d370016a685    = I2f363d2944c634905ef5ec14c9cedf52;

            I3954318b2392a82f2da71a0ca1504497= I4920014f5d017f4e840dc3b88526955f + I2d7715a3af03d9664729fa6df85034a2;
            I3d3edd06f8907f4369b825062348da87    = Id15ed601c43171647305818c6f30ace5;

            I15c78b909cbd04fe25820d777655d829= I4920014f5d017f4e840dc3b88526955f + Id32e7ad5b1aa825732d9b26d0fa02ca1;
            I72467ef10ecced8395a6870a39525787    = I75bed085cf80c0672fb41df1d6fc4545;

            Ia529c5ec88a9f6c14ceda5cad56b346d= I4920014f5d017f4e840dc3b88526955f + I77b54488bd26318f14b4364035cd1836;
            I9b74b672f55e7bf7560ba4dd2d0c79fd    = Ib7f95eeae4f4565133ae98a0538e56c3;

            I5b73c81f28901705f6ee26d63847db0a= I03b70553f1c501609400574ae7cd73f5 + Ia73cacadbf80c0701a5b5b430c0d5c98;
            I285b012d2fb5e2279a79cf8edca24ac8    = I5a7c45c0b4ce4206080f2b50cb0a169f;

            I1a9bd3f728db23b679639e5657ced179= I03b70553f1c501609400574ae7cd73f5 + I19eae741ef89baa1a64c403fb29f14f4;
            I8faf911a7d1ea8b0abe54f6688068ca0    = I27cba499cffd339eddcdb4e2c846ee69;

            I57ca72784a7c91cecbd694ddd08bcb98= I03b70553f1c501609400574ae7cd73f5 + I9d6730140c690037b5ca58aa30103f5b;
            I3dca974bf2d5631a47ebf8b945efab20    = Ifafce4fed1394ac5fa8849145960f2b5;

            I50f31ecd3f2b498cc7b759efa057f12f= I03b70553f1c501609400574ae7cd73f5 + I786338397f55073dce91e1c8c5f8e298;
            I12141c45d147b058a9e392f3b7d7d06e    = I1d6de59e71e329f79055285b3a50c2b4;

            I8ccaf29848defdd264f522642968fa29= I63c9bf68b43ed66c51b0f4c0ed92e9ab + I0f277bc88d46a4e6e9f1f2c410b503fd;
            Ia527c96e30b782f837bc6206961400e4    = I9265fbbb34a66f13193ea1220ecb0589;

            I808ea92ee1340876cf1d2c47255dc2fe= I63c9bf68b43ed66c51b0f4c0ed92e9ab + Id9d56f09595e80d66c2ac300f7d1d972;
            I6adbdb64422a08be9bf9e538db97463b    = Ifcc01d5d37df8c68972086c44575e8d6;

            I3da806790125328b626be1949f71267a= I63c9bf68b43ed66c51b0f4c0ed92e9ab + Ice780b1695a8e80607a03dee3c426ffe;
            I958cdf5367c7b0bd58b70b763d3af8aa    = I57c25f5b2fecd18092653842e49e8d11;

            I55e59bc1daeb8b2be3d7a1e4b272df93= I63c9bf68b43ed66c51b0f4c0ed92e9ab + I0e5931219d94c8e8e1f4af081404dcab;
            I91b7b8e8887b5dd9853297463c55b78d    = I4b70004412f2ef37ac00fc19592b1f30;

            Ib0ffadc6a0091ceff91ad1fa435413a6= If408dfead07757878cc878131bc7d6a3 + Id081512cd113e4d09df0fb13e443d76b;
            I6162978f0c57958ad0403246fb0530dd    = Ib952f8ef85514b1832324867adc72ce0;

            Ic863f139e6bed2d06789a07c6dedf6f8= If408dfead07757878cc878131bc7d6a3 + I38cc7b117c0bcd5e3060cd370d710d7e;
            I508142e70fd04513977130556aa574ef    = I08494381ebeda641f05b917fa31910a8;

            Id0e8f6ada5060a911090f76cfaa3c6bf= If408dfead07757878cc878131bc7d6a3 + Ia98a70144e466b356d2998948dc4b602;
            I2afab673e4b803ffd888f187de47fa49    = I3f0568074c465ac281150bb70bbd76ec;

            Ibb8c9b8fc9b58f5f8a6ad342934804a8= If408dfead07757878cc878131bc7d6a3 + I8d96b419b010f8076311420d7b9c8a18;
            I7a56f81596920126a9ea2c9fb3a19285    = Ib6b79505990d6499127f78e3186cc2a8;

            I9323a188737ca54c2dd553cd99bd416c= Ia0857d63d309807789b6ff4f6028f1b3 + I2ffb7c2ad09bac694ef13ec41e5de327;
            Ic6252de2c819f2243476ddf82e22d137    = I5404c19d5b4c44dddcca70138fbe79de;

            I2694cef38855f496e7ca12f42dfdb9fc= Ia0857d63d309807789b6ff4f6028f1b3 + I81800fb49855a4fd2737faa07ff15d29;
            Ieea8672b2f23711c6ba893de5c5d8bc2    = I7265ecc942bf501ad034704f517d4e8d;

            I75790b4c0b1f6c7935f5cfbea26407d1= Ia0857d63d309807789b6ff4f6028f1b3 + I9a3f0b4867087790c78f674b719dbf7b;
            I3a4dbdf517b8f9c93b567f91870e6160    = I1c114e8dfd37b1d182028679b3974a1b;

            Ib8b366c47e56a49fc53ea4a9e1ebbd99= Ia0857d63d309807789b6ff4f6028f1b3 + Ife13f962c7a8df3845cde104a959f678;
            I4731ee7a0e08c69e2bd2a8bcea0838c2    = I9fa799fd606c85184ce84138a90f03e1;

            Ie1c86256df2bc6c4dad41237eca41986= I53921b825c5e434b63bee0e1ecb7a517 + I003f95fb8f2027efa41a1936e8b53986;
            I1b6cbbcf01a65cd1c2f1e241f849c904    = Id8b3ba6e7ffd04674b2ae10b928f26f0;

            I7c9e3f97a94f9a078c209a1b84ff916d= I53921b825c5e434b63bee0e1ecb7a517 + Ib190f589f4d663dbc0a3c166a8dcf5fa;
            I663aee79f824c854f57c19e87207529b    = Id4cc4e9883ae7b27bed350ba292d9349;

            Idde839d34403fdbba62671b83801ea8d= I53921b825c5e434b63bee0e1ecb7a517 + I49eb064043f91112c854e31e4eb9b885;
            I34ff7299c9d83affa4512b7da302c199    = I5c3099cb6fc046e62863a69945ae3e04;

            I824e23c3e43434e0a7bf8c8b8e0de597= I53921b825c5e434b63bee0e1ecb7a517 + Ia0868eee7e7e0640ce1a4d3ca9c001cb;
            I70ca6c9d0a5c99e0036479f7b5dd760a    = If48b274e1e1809931eb2be69a565a443;

            I0f83a2c488c229e971030fc66ce212f5= I53921b825c5e434b63bee0e1ecb7a517 + I7f701ff37ad3fc34d2f4efafe5ff5351;
            I835bb7345787eaadc41816858e0a71a1    = I1667cbf3caf9a10527531b6aa69df847;

            I8fdda3dea7a63fd6e57f70365d7b6571= I5e68f84e123c37f19a03c13892c77e19 + Ifcd68be4bea38622d2d57d3a4e6fc5bb;
            I3c7f6fdd0e9cc7426df76027912d1ccb    = I80ddcee29ed7af07148977eddab4bccd;

            Ifa2fc30c14c549339edc65c3670d90a0= I5e68f84e123c37f19a03c13892c77e19 + Ic634d26fc09589a29a160e4efb5613a8;
            I9ff512085174a7720705d0fb37c4ec34    = I32ab257af6a54e78706c6d83b579bcd6;

            If69bb1bfa10ca7dd37ba57485c3429e7= I5e68f84e123c37f19a03c13892c77e19 + Ibfe760474fcac99f1e5ffa2e008fef99;
            I6a69cdf2bae1ea68c9be56dcc4e76a59    = I907f4db1352049380285f358cac2b439;

            I2ab0738fa2d5916d77a81b9da2315376= I5e68f84e123c37f19a03c13892c77e19 + I51b5e641856239367cf43f9b5679b268;
            I855ddead34ac131137ba644afbfea2b7    = I22cd5fb22f122d99e37e6c1ca2666301;

            I50a9ce776ad2ccd8048b56ce101c80d2= I5e68f84e123c37f19a03c13892c77e19 + I43c815a8ce0b2df9744a525328969691;
            Ib1a463388daf270eb0ce698d7b5ded4b    = I892abe227878c5232de3ccd90e8c13e5;

            I9c9d0332ee7ad6a3488b7e39bcb06ca2= Id5270b57c6fb4b18db3bbd0a523e467e + Ibf565bf1803ed43120fa54b80f6f1f29;
            I74e4bb7530c02073f9b15a6389659d4b    = If5086f7447696a697be414fe50ad91fd;

            Idc155814976f0aef9b56b2bb3d52b3a5= Id5270b57c6fb4b18db3bbd0a523e467e + I66b92f1de2cf408c3af53b161a6ffa60;
            I6721b13abeddc76139bdc7380434cc2a    = I9dc20c15b19d9351497997c81511c744;

            I2e02fbd496d08acb3ad3359b49b9f680= Id5270b57c6fb4b18db3bbd0a523e467e + I5b937934e7aae1f916c2848889f12685;
            I84fba239c5705bcd92096e204cc9438c    = I254c64de80d2a159aa0b3f3170042079;

            If0f8b3dfce99a5a75c2105d45ccad985= Id5270b57c6fb4b18db3bbd0a523e467e + Iedb655aa25e5f0e35137ec6c3acdc527;
            I4d46e4d50176768fda897949545e2125    = I4dae38e87f09d78c748974da00f274f8;

            I6790223e6a7cf136a7e2b261ba4fdb0a= Id5270b57c6fb4b18db3bbd0a523e467e + I6c4a1ded9bf39091cf302ebe0103e2f0;
            I57086cfab3b163c3911c3cf7bfb3141a    = Ic8edf24599f1eee2af3576dfb2a6829a;

            I6a9643afea7a6cc9b94806ccc8e84c0f= I3c18a84617eb21472d53e598700d7f4c + I94d9412a7b43fa0bd4b9a6d32d313fc7;
            Ice174debd5dc911fdf5d5756cff8d731    = I144ca4c629cc3134a991414038cfc9cf;

            Id3d19d7c2b941930478a7ab01049e390= I3c18a84617eb21472d53e598700d7f4c + I57a0f8c3710cf8e216d6dc2420f7621c;
            Ie369670edc5b602d305904f3a4a4381f    = I379ed527c944420bb59be58b85ab4704;

            Ib0a25312d51cb6aa1741f7e425bc5cd8= I3c18a84617eb21472d53e598700d7f4c + Ib46b13498ec14ceaa56719f26f18febb;
            I41f66f79339962ef42fab3b88e571170    = Id37ddd7be0621f84793d1600ce915236;

            I44dd1b66f5a9a6b0b976d3d61d6c5cbe= I3c18a84617eb21472d53e598700d7f4c + I78ade92efd265027807c861be44a10af;
            I5cbd2fad4d90bd77ba3d2448a37ac60f    = I20bbdbbee46a2be5c6caa56786345e8b;

            I3ee456f2f0e7f447ae92b7523136adb5= I3c18a84617eb21472d53e598700d7f4c + Icd4ff8d14af2699db2b5168027894ebb;
            Id86a2869148e2885633d9e277f7041c3    = I02199c9dc39a2c8be49a1c96aa89de15;

            Ic110e2a08b550acd3c8bda4a1bc2bbae= Id36663e7a01fff3170833ecfecac1321 + Ie1374cac341cf353b1863dae9f544e8b;
            Ifb7b585189db23efabfb522c9b45bede    = I17b1742efeadf5df716128d6603ebe99;

            I3f87162d2874effd66a82f821aa6c73a= Id36663e7a01fff3170833ecfecac1321 + Ie018f3003c5f124bddd13c359257bf35;
            I7763f0d28d8065d8c94ef8df96b2ab06    = I68da2c2a43373cf8145e6f7072bb5ca9;

            I660ea6d341fcb38f108270c08d82473b= Id36663e7a01fff3170833ecfecac1321 + I90b0296f5ef87dfaa6110fc2e9d6ed9d;
            I115ba88588187c7115977e95bd26ee5a    = I27f3ef61a2ffbd4154a7b683aacd4844;

            Ic128d603fc08affd2f3d0ab3425710e5= Id36663e7a01fff3170833ecfecac1321 + I0c59e8c82a31aacbf5977ff778a7ff49;
            I6e7f2bdd0c8231a3689893ef4877fdba    = I0726f4d2f2b1d495b1b439f998193435;

            Id5372641727970383a59e08f550814b4= Id36663e7a01fff3170833ecfecac1321 + Ia79d52fe2130426c07890fcaa50137db;
            I546c513d5357ac1a6fe669888dfaf717    = I05e3c3e8567ed11012cf9f9d7ecb629a;

            Ie99ad992d66880542dcd330ef6ccee04= I8d3be15109c7007a79fecaac0d891626 + Id28d9545e8d20ac080fbac5e345692da;
            Ib3e12c614471912d0b276cb9f0382b1b    = I210ade98fc479cdb069e2b028f1920d4;

            I9ed0b194f7d210d57c54b289e01c75e6= I8d3be15109c7007a79fecaac0d891626 + I924514226fdb5bac110a2650bcb2e85f;
            I7187a2499e3319da90b6d6fc64411b46    = Ic89a704c9de69cff5b09d1b3bb220fe8;

            I227828831c4ad21b06ed00fb5781b0e3= I8d3be15109c7007a79fecaac0d891626 + Ie4ca0836695d951ee09622892ee35928;
            I9b46582473bb4dd5541a35ac708486f4    = Ic8ba8abf8a87610d08fb5a8174639f99;

            I09d5ad12cb836adfbb4833ee80fad2c9= I8d3be15109c7007a79fecaac0d891626 + I2bc5a10c587d89d10021aa5eaafb490a;
            I929796fe327ee9c8a05e6bb683ae5d7c    = I9c0a1bb49be6604f75611b92d937c124;

            Ifa9c94ee94e4beb2e7c8d2d57150df41= I8d3be15109c7007a79fecaac0d891626 + I308aaa8ac500b5589aa4af533a9062bf;
            Ib6638da8b69373c2026d3f5305825cde    = Iff70fe838ee16e8e35b1034135555acc;

            Icb88e59e194db215382e8e949603a9be= I92169cc57291f20d336a479e392ec271 + Iaa164a078c8cdaad694a053c9c1e0313;
            I28c26bf4cf9693d1807818b2ca7883ac    = Ibb4daaccffcf82b4cb4c431923c71f3f;

            Id4ebd28aaf1076acec266666f88a02ad= I92169cc57291f20d336a479e392ec271 + Ie2d8c84d8c9a4c8f637068a2ae39fdde;
            I291fc4eef4b80d1020c96488b869727e    = I9c1fd2b57c1756bf67bc8cf5ed4a1912;

            Idf0a0bd862167392357501b3233a8d8c= I92169cc57291f20d336a479e392ec271 + I138f008a6206a1067bb0e22ce3d90990;
            I53006ed50f6211439681aa7659647e35    = I71d437815bcfb755e16fc442431b6f68;

            If94cdb867ea0fc2c5578b16aacb1acfc= I92169cc57291f20d336a479e392ec271 + Icb3ab2c67a87b2ee158e0021b72fc186;
            I47fe32973727237ae0cd4c306c7efbfb    = I4e3e1eb8ea6dfb08ea2634a9bab8319b;

            Ib8c066b0700941a4fa739820ff12b948= I92169cc57291f20d336a479e392ec271 + Iac91f4037e542d9fda30fadafe7e79ac;
            Ic3e0c7d71f13a56a9a63e158c7f2cfa8    = I1fa2749e15c3bd7253a023eb01140cc7;

            I11e0f8dc46b286bafb05f901f968e1ad= I6178b220b469b40dac39168057023a1c + I459c59ac61179d74170db53bf45ba89e;
            If383f241447cbea4e18f4f79fcdbf144    = Ie19e8502010d0c178f9f2da8df3fa63d;

            I608537f5639d5e0cd3e80453e21f6f85= I6178b220b469b40dac39168057023a1c + Iee8f9b0654f6f6797f11cae0947e454e;
            Ia05354d3b4f61299d5897832639df2c2    = Ia512ada6f00f86ff495ae12ead6607d3;

            I0e9d8db1bb6347c9507b645132308b3a= I6178b220b469b40dac39168057023a1c + I9df5b63f66c162d517daa69f5d0e6095;
            I9faec40665477e8b3237773d606af2f0    = If7b2398d3426250d73917539ff743c8a;

            I17033b417fa383a2db41d157df33d9de= I6178b220b469b40dac39168057023a1c + I2d1a5645b126761fc7fb70d24e37189a;
            Id231ab3133d4bed02aad7e5f560ee5f0    = I6446a839157f78880fc3fc7d8c378c78;

            Ib7f45dbcad513b4dafee60f33622b0c3= I6178b220b469b40dac39168057023a1c + I8cd5970682bc84881489c12ff073212c;
            I13616c8c7be221cf4d2c13ae87c38bed    = I53504e8899a821cebe69ed590a3fd7fc;

            Ibfbd8e00e00272f32428c7b4a3c53050= I55342938216a0ea0889f96c2f6c05ce5 + Ie16dc913f571ae73ce03d755077345a9;
            I8793bc728a4d423fb96a88c83bb9746f    = If7d5fe39b147f24303884de3a30d669d;

            I27973d1d4e07eaa49608d6f6975d0a93= I55342938216a0ea0889f96c2f6c05ce5 + I7e0474089ebc1c34747be1bc17a81d72;
            I2fb6af0f152232550a3cadd55656df20    = I24c005d076b3c887d45d1285a4fe1bc5;

            If77fcedbcf99f89045de87e5cae45d8a= I55342938216a0ea0889f96c2f6c05ce5 + I48ad9b737892d7c49340ed679f46e034;
            I5144918fcd4ce1a061644240730fc52a    = I18e00688f19c522b305d223ead684fb7;

            Ie8f8691820e7a560db8116f38dae5d49= I55342938216a0ea0889f96c2f6c05ce5 + I1ee27be7e1a38aff0039b21c45f406d1;
            I1821eb21cdf8208ff6c2f28d963f7bd6    = I0258ec63762460afb41bcd6e8869ec69;

            If0b19af59ad851aded19970494514034= Idf28431c76a84a48dd895979d2b11a63 + I16deb9107193a3536979e4b5e5654b9c;
            I80471575b1d4b69ef073056f798394ea    = Id1280129b20bd6389618695aec9efeed;

            I98b8e05818925a4b65082fa57affde83= Idf28431c76a84a48dd895979d2b11a63 + Iccca1936f4c1c9496205e77b588e9985;
            I890bf9b72cc3c71351547178d72796e5    = I907fd3abdcadda1cd7149c7cf01e5751;

            I69317e8c556ed67630829c990f8b74db= Idf28431c76a84a48dd895979d2b11a63 + I1b40adfd6fa6c943dfa8d230d9e65514;
            Icc9d28b84fa91028ae96cc9b8bae7555    = I73f044469c4dbcd5a98c0f83d6d043c4;

            I9147d103cf235310393f9339f1cbb376= Idf28431c76a84a48dd895979d2b11a63 + Idf90f01353ad1057e11fd060442f4e53;
            I0b0d167c415f8c14594bd61907d46d80    = I2934a8783b90254606bcd933c629577f;

            Ibe0b2cab6e2d3f3cc8baf3623ff50988= I1ef61124c8d62e8f6a82a729fb091694 + I619957528c630e7f64924a25127c93fb;
            I9577d49a74520355e53a1818f479db0e    = Id26b2a9c13424769e1627b1549159a7e;

            Idc64f1443dd2497dfaa223cda3fbd682= I1ef61124c8d62e8f6a82a729fb091694 + Ibd4aaf02982068ffbfd1b8b3795d9217;
            Ie6e888d582ba9e600e91b119e2804642    = I2115e45deea528402794afadd17d9fe7;

            I6e37e92b812099985436851da8a6ccb2= I1ef61124c8d62e8f6a82a729fb091694 + Icd37da8ea84a606529e32b2db4eb7f5f;
            Iccfac3d489b4b110d6b6e005a5ba45d8    = I978020f8aaeb98cc1cea9360ec06da22;

            I057df2bf67d5580275654bdc28b40027= I1ef61124c8d62e8f6a82a729fb091694 + Id45f4e0f142b6c3925f24a37dcf7c0ae;
            I69a67481ca8fd01dc5400dbe887b4f83    = Icded30641e4770e30ee34bbf8d2a5721;

            Ie87a151c8b90942a899b8167bcb34afb= Ib8bb96f0372323e6a8072ca56fb9396d + If13e359e530823319046ce20027445dd;
            I1f36f045becec7f0528f4a935d3da2ff    = I02e3cbacce4e97e3088360f0acccee44;

            I735752035af159b48f53d8302bb33c21= Ib8bb96f0372323e6a8072ca56fb9396d + I24ae7de3549a84f4f88f561b6017b7a8;
            I530fe7720e3bcda35e940aa4973a7da4    = Icbdf81888af42710561aec48ce84e3cb;

            I1f26bc7cb30a9659a638e2ab65e1f187= Ib8bb96f0372323e6a8072ca56fb9396d + I485a48b4ff4da08f977425fd10e6d392;
            I03069dda9fa863172d8747408800eeba    = Iea3ce04a4b8cc466e892aab886e63744;

            If39a50e88c4a7c43428c1d15b0bfbbcc= Ib8bb96f0372323e6a8072ca56fb9396d + I52a9bcfbd2d3a763671f19cfeaf7bb8b;
            Ie7f36ee89f2b092555fbf8031d2347d9    = I3ca9464d884ccc7e2f396a74baea5bb9;

            Ibf966c12f049d603361ad32f55b0a2c8= I432f74dda4f6b1cebdf5ad59c659080b + Ia07447985347e9a7f3739bd98867cdfb;
            I18af7980562b28c537be3bea8dc5252b    = I7b8d02aa08cde64a409f3766f940233c;

            Ie1b3ed6d3fdae47669d3c4cb8af8d969= I432f74dda4f6b1cebdf5ad59c659080b + I4b94402a53d981e953c21ef316c709b7;
            I22ec20f9396d28ed39c5fc4bf060c44a    = I86ad427fe92cd4346b32ecf3c99c93c7;

            I4ec6c8d9e87224ecbe7c69d92f9419c8= I432f74dda4f6b1cebdf5ad59c659080b + Ie8c79e6a5378808c0ead5a4b24319ce9;
            I105eac4e38f4661c7c7ca32161e42baa    = I6667614b2fe12d6f63ac7737bf069b42;

            I2acb34de8c3fc53117a7ea4f9ce7dd2b= I432f74dda4f6b1cebdf5ad59c659080b + Ic8df04756f67e6dd29f3374c5f86d451;
            I5030734bfa54065cbef20c1350cd647d    = I909cbd582f015b4eabefd660b2039ccc;

            I7fa4009267e80ea7eb71194843c3b22b= I432f74dda4f6b1cebdf5ad59c659080b + Ia3cc6acf2cae41e560e09993007ffd2b;
            Ieccf25e3abd6bae7dcf08baf815f3439    = Ie3433004b0ea3bba81f0b7502c69c821;

            I6854329daadea2734e52180a41f56bcc= Idc689442305acd00f0f32416d8fb3773 + I4a5cfd6ebd47cda4fa2e06ba9ad6e5b2;
            I600c21fca7901299f8e95e8fa0ea0eb0    = If548fc27869a7e48fedc89bd5c8037f0;

            Ifca16aebaf75b2990188de201e4536fd= Idc689442305acd00f0f32416d8fb3773 + I2a3eb42a4402e873d081f94a14a99c20;
            Ic4363dfd133124dd45ec2211499d0788    = I7cc21b5c21f6bc0603c3d57c86feeb00;

            I46cc26afc8475f2fb290eefc95a542eb= Idc689442305acd00f0f32416d8fb3773 + I04a9c9765fd468a7e841577f09fc287b;
            I7c0bc779c09847e3beb0a139e8826511    = I9ce2b40cd4433999690bb6e5c368e9b8;

            Id746d6515cec9e60e7478898a09787e5= Idc689442305acd00f0f32416d8fb3773 + I9937af6fcf9d834f308bc3683d524981;
            If64db4386bf8f7d07292f14e3b313520    = Ie102c1592ae8606ab75b1f7101b44918;

            I09a3ad636db96e00adac78c3c94bdaaa= Idc689442305acd00f0f32416d8fb3773 + Iba0d2f08788f2208a648ae7b5414195d;
            Ibf51e537b992c4b4c0539dda9948f45c    = I23ef94c5c29e674714d4ea1ad2d3f0e8;

            I28b3baa225a5fd602c9fee9c948ae58b= Ida03738adc101c03c2229756bed2469d + I7eb76b3d17296fdae702d8f820f1428d;
            I9f83063bdc3c352024f702cb9dc71ce8    = I990c1f1dbce95ae4dfc62588c9cc9e1f;

            Ibe12ef0f56d875c7a44030882deb0e29= Ida03738adc101c03c2229756bed2469d + I928a0e4951208aab170656596f456209;
            I72127f6d422ec68dcd47126b87b3d3b1    = I9d2e71f9a6d7eb4221978fef3c10d678;

            I9bd9979e4acc4944227a4bd62b910c1d= Ida03738adc101c03c2229756bed2469d + I0eb3df4d4094e09e6c4b3c788baed61f;
            I0b4a1b48d110b820d8d87f6e94d32988    = I34754a80000aa92f8a7e4997b91f6d07;

            Idcfa802f458499150055dbe4b1ce8146= Ida03738adc101c03c2229756bed2469d + I7c6862830daffc98cb2c1fc121d82c38;
            I2e3aeede695007fabe0d6247a93ed403    = I055273589d8d967bd5e255808051a101;

            Iee010958cc3e9389cb8ecacff84fccee= Ida03738adc101c03c2229756bed2469d + I9f7df6ad60284c812aeb522974578e0b;
            I8c5ea3dc59fdcdea1c5f503dde1e815f    = I5142a2511a55a7ad420618d874b0dddd;

            I3d74b31096917c53757c829a67cf06df= I4d14c75f28f3e516c259ea288996131b + Ie5e432a991aff25577639f1b4ffd594f;
            I873c4dbe95220e40d7388870520261bd    = I5e008272bf3a470d74ca6b5cf39bf28f;

            Ic27031a9654db9459815fe0ca35408db= I4d14c75f28f3e516c259ea288996131b + I571ddcb0a10938e4c0816c965214b4a8;
            I561fa67a9bfbedffcb04e7a4d6b76a64    = I5c31bbaf08a6e8971f585cdae36384f5;

            Idf6ead2c37f75f3cde1d4b40cd73db00= I4d14c75f28f3e516c259ea288996131b + Ie626a24e3680f7d3995dd0c2ce60cbcc;
            Ia55752d6c4f20378ff570a661ab31d9a    = I509af9c5f9d6bf3be233847dbd05e3fa;

            I66a56161cd0ed67f65834b9eb0e94d17= I4d14c75f28f3e516c259ea288996131b + I5ab556386d2973354a5551ba9823e4ba;
            Ia13307be43e9155ed0333df62ccc8bf2    = I3182472e08e707cbc36d60ba54613129;

            If6de990e26ca9e8efc009188f8a5a4d9= I4d14c75f28f3e516c259ea288996131b + Iab1fb7006598181bd8749ed90c519b13;
            I07b3d1451487a55fbbedda48b0cb6c73    = If2455c2d04521a8d8c59965759eb328b;

            I8d866786bb2dea06f5b30f6ea80cff17= I6e6cbbf430d57f347a0d70558af143d8 + I72064a6a84ff956d76a5aa590bbc05a9;
            I9f8cf1a6cd0182fba35a49bd232f062a    = Ib759c72355cd6e146edb26ad106a0418;

            I01ca9a1d4901ec9b2a64300617ce4cd1= I6e6cbbf430d57f347a0d70558af143d8 + Iae32c44b88fe7ddb5d4f19cf8fff3ba6;
            Ie2e488a8589559deeec8598cf6726f1f    = I6826c8a05953c4df79e31a19adfa2693;

            I2dbead35e15afb9affaa6ad4edd3829e= I6e6cbbf430d57f347a0d70558af143d8 + Id6f7923a16cc5adc96a730083153ca6d;
            I9118ee5ff8c9ba9b125e5baa07bf52e0    = I56122ba51d99f9ca67828649860d409e;

            I83c57653e24cc09214075b04b06bad83= I6e6cbbf430d57f347a0d70558af143d8 + Icf19dd665616a8c96146b3ab9f46c741;
            I13b894057e2deae2c00787385de252a8    = I1bcda37ae1a26452a3443142fbee54f9;

            I56b9c1f555b24c2dc197168decfdb8d1= I6e6cbbf430d57f347a0d70558af143d8 + Ieef3b299ec35075c71ef9fb10525bfc4;
            I7797a3ea5b97b514a797243cf9fe890a    = I3f7dda67dc14fdf45bfb9c4e01dd7f38;

            Id5c48111f1b93de2cfe89f92fd182b43= Ib7487df45118e44acec6b9d07bbd5969 + I2121318f589878b4a9260625f97de518;
            I3af78697aacc410108d0be7fd13c686b    = I6fd4da8e1e3cb360964d6e425d174465;

            I32908c3c90ed6488357ce4869e8a1721= Ib7487df45118e44acec6b9d07bbd5969 + Iff142b88493149045fc0de355b767c16;
            I871cb63247618a543b444aa3f888fffe    = I5f7baab0fcf12df1e886e17375732c04;

            I16b4601f2e07e6cecdb5a030178e75c0= Ib7487df45118e44acec6b9d07bbd5969 + Iebee55168fb47664095b11c9f6641124;
            I124404013f8fc6b302661900b9ad8ed8    = I87303a5c7e205b0b1b196ae97a0c994f;

            I0ae08a41ebd0e6b402a4980478087bb5= Ib7487df45118e44acec6b9d07bbd5969 + I64f65df774d29696425ba460dda09b68;
            I8e413271c9d13748a1aa2d1a018ff28f    = I5ebd9eab33e2e8cd6b2f7c1f3bd2e39f;

            Icb57267a66f117943e964dd6420d7a58= Ib7487df45118e44acec6b9d07bbd5969 + I58a7c08adf48d0737c5803e2a818c045;
            I4d799e93b4dfcabd69977ddb25634a69    = I7f4bd63152869ed52c49aa41eea5ea1e;

            Icfa47fb87b74106cd3814adfce909424= I492f382fea500462b3d0866240fb91b2 + I62bda8dc70e0b5eb38abe094bbe92fc6;
            I1487f0027b7d16f4bc85bb00e537cbaf    = Id243e47daf8a5e75fe52a828af95b5aa;

            I63067cef0e1a348a3e6d8cd9bd88b907= I492f382fea500462b3d0866240fb91b2 + I632469889d6bb1c268b45fb805467ebd;
            I1a5cdaa10022adf0ffbbc0f58b3e690a    = I62bd2c30206c591bcb87f31543bda72e;

            I10aa5ba0f53632578c0e1cefa4bf4fde= I492f382fea500462b3d0866240fb91b2 + I9ca81c841a75a9ac242835956509e0fe;
            I98246759d003e9bc6676ceb2d093a06b    = Ic1238f5f1f2011fa1869cdb2f50e6a30;

            I427c0215d0ac047e8402c20610676752= I492f382fea500462b3d0866240fb91b2 + I546122346a22ad64a6ab2b4978cde095;
            Ia3c2dfb3c4a45091be7cfecfad11f3ec    = I7f2885836616ac775eb9406e8f5d5214;

            Icf4efa87688bd1b80437686eb0126057= I492f382fea500462b3d0866240fb91b2 + I30a1c8fcd9a510a6ed559f07dd809b90;
            I74cda651bcb24472a7697ba017f831a4    = If1608747d211db3fdf51ecf7464c494c;

            Ic373f785ddd1bf8eccce263df5a82c87= I3fb3ebddaf28efb56092d19a1b4695de + I00ecb5e329390023b318a2ceba0df231;
            Id7ba55b14ac0f471142011dc2d57cc4b    = Iccd84e19d39b19bec98dad532ea5b3ce;

            I56f8e8d2d7052af26528530d389b6dc1= I3fb3ebddaf28efb56092d19a1b4695de + I3707f68de059df0af5c652fc0478e543;
            I5890643c88c4255a0e5efd45f8af3ee2    = Idf7e508a586310bf4ca23c84f8240691;

            Ifb145bc18d435fb66779e7415417bc0f= I3fb3ebddaf28efb56092d19a1b4695de + I7b929c228c865112f00bc6b4dcc95b52;
            I4f53e4955e9e506a7169ae810da5dde6    = Ic8ef3162d3d0c57faf5dd1bddef1622a;

            I62a6e0c9952d6c6e6095e2364df93078= I3fb3ebddaf28efb56092d19a1b4695de + I463f4f370e1ecad71de44780eff10df4;
            Ifc7c1ea337b122fb720767f1890f1a6a    = I68115420b3b9b8ca8ca584c260e924ec;

            Id6405c2b2b9aea6bc457f1064d5f3ffa= I3fb3ebddaf28efb56092d19a1b4695de + Ic4f5e9d49419e1c57cfa387761ab643d;
            Id40d6f3a8dd09678b25b3e579dd5fb68    = I5bac906cb51bae905ea33717fe015201;

            I079df9611bd81f672f2ae028bf267995= I22a26b7f0b1c8c16b00597732ce2ab23 + I28cac65a4db3f708cc90a1b023bfe894;
            I7002830b0a5f40ba2a2fe7a00c7b6d58    = I9f261cb4883275f5f9187a1a6e8fee08;

            I096b226cc511363946a39307a7d97867= I22a26b7f0b1c8c16b00597732ce2ab23 + Idc57f37015a48393608e2b026bc7065c;
            I3f377e8994959ef8182a08538e393d9a    = Iecfe32305d22e6d91c3f7d4af2ad9d2f;

            I4cc42c5a75ef339510ee0e86fb44e16a= I22a26b7f0b1c8c16b00597732ce2ab23 + I385d03def4cfb49f54867687ebd710ed;
            I71bf29f3519e3238cec112ef97ce0579    = Ib30aa869fd577fb3315608a85947dc7d;

            I680c01c3327cb9372a42c1ec5b4193e3= I22a26b7f0b1c8c16b00597732ce2ab23 + Id3dd71ea0bf0f2996fbe42b8c3318762;
            Iaa4bc2f51984f383479b597e6cd4c873    = I82209dd60aeaffa4b05b38230c27147b;

            I83451a072082194ecb3f9419edd728b3= I2ac08a2d8c917ecb37fbaf5325cb0473 + If3cc31fd16469339470702045fc6d0da;
            I9066a5cf776f80ebf89bdac1f2edb4ac    = Ifa110a9cdb359c2b0567d25d4dba725a;

            I52ad85b6a1c822ca8c2459bde8fbd510= I2ac08a2d8c917ecb37fbaf5325cb0473 + I114c595caa67a3f777f087a634130a6d;
            I7319203d7231bebb6d6e52422cce5ed2    = I1451eec261d2367ec6e7b2d50a20679a;

            I1c44d2ef638825862061a8ee1a0a2f95= I2ac08a2d8c917ecb37fbaf5325cb0473 + Ifd3638d44e1ba2285891fac152dee327;
            I4e8309976fd6011d78728cef935dc3c1    = Id8f178b6565e3a57c5370aaad14f0639;

            I8fa1fd425809cc39cd8e2785773c1d7a= I2ac08a2d8c917ecb37fbaf5325cb0473 + Ib834b91bf81067e8efa9d470023e8b9d;
            I5ed502118c175d5bdb4607973554a3a3    = I67fb672706bbd331c27ab1eb386c24b5;

            Ifa22335f04d35680eb8cfec8f862f357= I50ff8f51e75fb9ce3db983c2a0f57196 + I221777352b48c4e228c6637410113854;
            If457f80b3d29b60b840f886fa928297c    = I112661c3273bde5c91b800dd8ddb08a9;

            I6aff673c27811b81530453906312aa9c= I50ff8f51e75fb9ce3db983c2a0f57196 + Ie3e54a4700d8d0f6478187e06cb6f85d;
            I7e0f785ec7554540c9a4a413a3afa75f    = Ia4979ed96ea3e7332635e1f1a14d9ed4;

            If674ac0540f457a21235664c213d4923= I50ff8f51e75fb9ce3db983c2a0f57196 + Id5e02d4c48fa6c3b0d45a9e66f09448f;
            Id3662bbe1b5191995d1656045fe6b6a6    = I11a094c5fa993419d19f6361157d6ad0;

            Iac223ac498bdcf2cb2514582aeaf76f3= I50ff8f51e75fb9ce3db983c2a0f57196 + Ic6ead78ed741442f17a15a157cd6ef9c;
            Idf922fab93bc2357ac1f66f73f3ead0b    = I38007605c51aa852477e1901bdd292f0;

            I7f40931ab78ededfcb52ccaac9b81282= I444bc340ffb7ef7b72d4d2e761d58872 + I86e53eed5b857c439039238bb486067c;
            I780371393ef898aa144c5bc36e74c654    = Icae30bad38ea69b85fa826ad52e25a51;

            Iab7c8dad0ca20eb0988fbd99f25591a8= I444bc340ffb7ef7b72d4d2e761d58872 + Ice18bceb10fec484ffc96155e14c4974;
            I79696cd10cffa4c0181a2089da6b3262    = I1afd8ef52cb1eef06769b7a27c95fa03;

            I3cb5f890a5bd3daaae34c8dfb6ecfc49= I444bc340ffb7ef7b72d4d2e761d58872 + I3afe987d8f2c93cc19534a3221d1939c;
            I073155ab0359a13b77f730653dcfc08d    = I9c5442889b71c19de290cf33fa393bd9;

            Id80e145586d7e539a6514dd67ebabf6a= I444bc340ffb7ef7b72d4d2e761d58872 + I4e257dbd6f196a02dc0f5a2e5f6047d7;
            I1b44f781d81438654f69bb7fbdb94011    = I772891870fc29b32eeed162f198217e9;

            I01e09bc554768f30dc490041d19b4da2= I039c6cac5830759529595a958b7f65c9 + I89433799cfa534afd66e8d6b9f1b62b9;
            Id68f1a0ec8ff80da3190fe517bd935e3    = If4167812b028552487002b44bdae0caa;

            I0196f7df6f834ae20c4fdd127e66104d= I039c6cac5830759529595a958b7f65c9 + I223b05d94c09b095d1988df121aa5e37;
            I3704464d41956032b779eebe27511815    = I4d470ec03c4967c49989f59671d735bc;

            I4669c4f256c123a0fcceb55c1e72193a= I039c6cac5830759529595a958b7f65c9 + I788c64785b992c675fe348a1fa181525;
            Ie6756ee9631791940ffc6fddb223b4d0    = Ia28efddccf0f15c926e3901002bf6c9f;

            I4a02ffa2a79df824f406909aa189a404= I039c6cac5830759529595a958b7f65c9 + I3dbfbd34d1fdfd4f422d900154123b6b;
            I085151dfc2e773a7a485f5ef1b7cd6bd    = I1f3c6900aaf35b7e0cf71c04d917cb71;

            I3117e5029119e70846dff61d746699e7= I0584de7d919236ab138e288a27d08ff1 + Ie763738b7faf253837e1c45de255cb5e;
            I2654e83fff153df7760c341f59a23396    = I8788a098d0d9b94af7b93f6b5ef0cce2;

            I1e4e705b3bda1451fc384cd934c0bb52= I0584de7d919236ab138e288a27d08ff1 + Iea32ebc385c6cfc9212ff37973a0a05d;
            Iee3eec7a9d7a3a5c22281545ec143e50    = I46a61c4cc712f8ffcf45f93d11f0e146;

            Ib5bea8e0072de3de2c8431ea6a35dd51= I0584de7d919236ab138e288a27d08ff1 + I449c77140475475b138d839a74078337;
            Ied2b9ca07a6d498abada30fb0726df24    = I2a826f08bf1fc30c125cdb9a93bea1b3;

            I7d9d94022ea95ea01cddc237f3df8cb8= I0584de7d919236ab138e288a27d08ff1 + I529b763dace1924613d184c6c70c2708;
            If95315702519e7a08386a870e599aab0    = I2614ad9be5eee336ad67441c050bd366;

            I3f0f9aab07427fa81fc3096c6b6d3d6d= I086402c82ec67ae09a9e6360c58904b4 + I338ccc17dc6158aec0129c8b0c02c429;
            I1091064aef7d915ba8fb6cbded069102    = Iecd35290f27c4375873e964f2db90ba9;

            I12a7983041f9c298d533bad58f41d24b= I086402c82ec67ae09a9e6360c58904b4 + Iea74ecbac92e1b8f2ec7ad68d10b8e7d;
            I40685c7d2c8be12698f734ec6213b5b4    = I9b90edd08194934b456cf88beedf8785;

            I78503880e5c96ec0a03c75266b1226e8= I086402c82ec67ae09a9e6360c58904b4 + Ib0b46b99e61d724ae664d9d1fec1e29f;
            Icc7775fe34c162006b93662530fd4944    = I7db63c5bb5e53cbc83051b5c80c1a19c;

            I8adeae445b33f634977957bb1a2259aa= I086402c82ec67ae09a9e6360c58904b4 + I7a600aeb6cf8c3311c10afa4d82767a1;
            I2e6f1a5695ad23b8ca282b344832ee8e    = Iaec5353d68ad9092c0fb74683f876213;

            I73bd13f381d15e0b0198b60cee44bb42= I1cefdc831c146187c77f861b3e2d1af0 + I1ee46fec2b82cf8e5142f8e2ac5d9d8a;
            I016ce894bebdaa7e56af9deb1ccfb3f5    = Iec7f88e1ed763c1f55c90b39870875c2;

            Ic8b651c2b043a4a6e4cd259774322230= I1cefdc831c146187c77f861b3e2d1af0 + Ibd8424c228f87f85df3da6204edff2b5;
            Iad2dd0815c1107160992e5070632f76c    = I32f96b4803590ac0f86d2178cac9e4a8;

            I76979d7df582f9306e796a03cb540963= I1cefdc831c146187c77f861b3e2d1af0 + I59d4567d3355fdae5660a1364d1b8d00;
            Iefaba2acd282081b9a0a98ed057ca85e    = Idc0fc3de3b05c5beebbf24649662f02e;

            If61d4585986757a525c54589ec93d8c6= I1cefdc831c146187c77f861b3e2d1af0 + I8c7aab31f8cb705ea13a41a5bd349303;
            Id4ef94eb8d5db8810bca4c9d669f0b7f    = I9d54e626fd0b2e435b117ae6b5d5e194;

            I1bc5766a4a3cc2b468ab8ef62eab691c= Ida9c16ae57d17b6faee8a54838860447 + I4f72d0db9fcc358c6fbec9964fbe0bbb;
            I04e845e6a5ed71978b636593dd749b12    = Id5cff86905cde551a008a19305e87f94;

            I21585169e5fceda643bd03fddf8153be= Ida9c16ae57d17b6faee8a54838860447 + If6d436031f68ef587750c5c1dfcfffc2;
            I0b2760b437be2cb79382f8d6a7b8969e    = I3837a2e882da18f37f074b51cf5cbf85;

            Idb2990946f60939136b3bfddbc7b1671= Ida9c16ae57d17b6faee8a54838860447 + I2b54a135e59945901e9c11580a29ee3d;
            I1b0fdaeebe5fee6fbb2e13aac5e233a1    = Ib584dc3e5dd346562062794c0f1c5f9e;

            Icfbf703890f684bfc96decc429deaa04= Ida9c16ae57d17b6faee8a54838860447 + I171149dcaab2c0f0e2a10547ad95084d;
            Iee872d17e4a28075be0ad7086c3acc91    = I20ac1027f7da12ad62120cd3b0603c7e;

            Id5bb42639a1c1c1d67df1c89a14a2bfc= Ia3b9fb112f39dd0ccbf7555659369efb + I8a7fb51566bf215af214cd2fb5209974;
            I87656ddd4ef8f1ae36c7566d5e7892d8    = I8adacef11a4f33ff1ccea285fd1a8b74;

            I55b8ef91d667c1c1d9e58dbc86a2288a= Ia3b9fb112f39dd0ccbf7555659369efb + I97a75b8625ae2a143cf364790ae77753;
            I865cd0535644db7f17db1180c85f1744    = Ie2ad82bbff584541911e13b90a5d15a0;

            I17ff683da41b469c8c8b82ee32a7378a= Ia3b9fb112f39dd0ccbf7555659369efb + Idf8ebc0d747ae143aa61866e33d458c0;
            I71d46741fa94df65e1bdf6abff53d2ba    = If6243c5fc2ec9a15eecf227b234434d1;

            I51f10296c38872338ec7df35ccd520d8= Ia3b9fb112f39dd0ccbf7555659369efb + I23b60ca4da2df0ec40c1df62d058deef;
            Ic223d7941250d739ce9bb0ae5013646e    = I41f34c28805f2653586d89312f73237f;

            Ia59ff33765ddf4aeb17f90a70c01d76c= Ib1bfcdc0c972aafc99116ed8c0511445 + I5f73e5faf1aca83ee0a415c9ac4a1b9a;
            I1ef9b548b943a1f2012b91c7e0b445f2    = Ie2031e8a9632f0b98f617232f7c462e6;

            Ibf97abffb1ec40f2f0e099a814e04ab2= Ib1bfcdc0c972aafc99116ed8c0511445 + Ice6db5ba70d3c7499df6723a2df56bfe;
            I88b6d7894d82ff394e89c7471c80dd5b    = I9d706a29e764935ac3cabdac4e95af1d;

            I3efc3271e18a1e350473dcf3375088aa= Ib1bfcdc0c972aafc99116ed8c0511445 + Ic0954671eb1dc893c3932e456800fadf;
            Ia5fc7e1f991f30042b848888a546534b    = I7a2e1620640d2060cbb0a1bef5eb79c0;

            I1efd1220ea9100f2fb4f169ceaf462a5= Ib1bfcdc0c972aafc99116ed8c0511445 + I7978d2d800b4438d0644ae3df6bcac9c;
            If699df4c8261ebce5c5d1aebe062cd61    = I2795513c5d99dc8e09be4bebb4d12944;

            I9af399f27c8e2b62b7f3fc6481ef9318= I7adff505c50450a04f1717cac1adebe7 + If845af0d620024f04525244753ba5d18;
            I19338369553e96bb2476d80fe84dec3e    = I03cb6aeff54e7e9e2ee809f8bea621bc;

            I171bb4ee9be2f92e4d82997108572426= I7adff505c50450a04f1717cac1adebe7 + Ie7820d1a242bc28c19ec32d2c91e47b7;
            I9844ff02042cbc04dd5f4179908bbb2d    = I78c43fed329002e5ab9a0e429fb3b769;

            Ib13cd76c20fcaf95f26f4914380c4fcf= I7adff505c50450a04f1717cac1adebe7 + Id50f18f642f3b00ffa34986f78a0eae6;
            I89cc6a060b714985b24f724adc782e7b    = I639755c3c20317c18359e96fce8e2f2e;

            Iafb219f1c8c6883e01fbfb4c887c8d6a= I7adff505c50450a04f1717cac1adebe7 + Ibc4eddc0f1768e9ec7e38e951a28ec42;
            I39d94ce7fbe37a74404e0043060441ed    = I68c7cb0d5275b576e4021c8aedda4646;

            I94fc9b0bdd2b0a89a9f6351f1fdd4ff5= I699feb4382974a02b21cb387c13f7f3f + Icfef12499b53cd84f0aae067f30c17d0;
            I0a1c9a8d59dbcffd6847f3a65107c407    = I2bd974f363231ecfaa9ef8d018a02936;

            Ia9ceb45f33402293c162cef4037ba007= I699feb4382974a02b21cb387c13f7f3f + I1039bc43e88eee527d2ed6adb8c7d1ba;
            I2328556c467a9e639f2b6ba1d0cb99b7    = I675d5b900c6a4bbdb8f14db50b873893;

            I0fa4e12e62e8a30b3b8045143b344b4f= I699feb4382974a02b21cb387c13f7f3f + I5b64997d083769666741c794dd92fb7f;
            I5c9d75d6431d69db1abe412e591000a7    = I36b68c4fcf7a2adafce004ec0e231209;

            Icec1c637d24ca277bb2e488257e92a40= I699feb4382974a02b21cb387c13f7f3f + I1c97fd1d21a31af8b5498a79b1a3e7b6;
            I8dc3dcdefc85b6ff8ecfa09cfc7e69fa    = Iea5c378e0635e3bb31343988c4dc6259;

            Ie9aca08b988fad20904545fe070defd5= Idc99c3b23e49aca3c98f0685ea34441c + I83d71a89f35eb73265ee3e54184e1277;
            I69f6c909ea6b207c200b154e00e13a05    = I2edf197a22f055871ed9b54f9e1a874a;

            Ie82304b2c8583f967649475e309e68fa= Idc99c3b23e49aca3c98f0685ea34441c + I3caf1211dcbcdc746a3e4c7fbbdae4a8;
            Id365c9f8f7f97c777bd5da0ce9490511    = Ie80e559352812ffe4d9cf6006af19e85;

            I60da0fb8a2c0669d5f9037ae99b23565= Idc99c3b23e49aca3c98f0685ea34441c + I49f5f87662fbb540d72c94bfd1acd060;
            Idf0206d2ad2bdef7db1d30a2d715cc6a    = Id2f23da93344ae523d495478dd559ded;

            Id8c19a3547c17ed513d2d857adc66885= Idc99c3b23e49aca3c98f0685ea34441c + Ie4f063eeaf7ee3f033e2a01ffaca623e;
            I07d1c54431eed887554a136f15f86d22    = If18e431ab87f137467f6f87e40b9c27e;

            Id74984743844e9495ea0f528a391f4b8= Ib67318fa6954ec8f3247927d34e74f8c + Ie45aaf966aa0a94803050b5f43d69e6c;
            Ic16809a3c82787ed88819fc9e9613f85    = I3f5b5d6b646070d84f2fb963f3824ce1;

            I9edcdd5b927b3f6b3a4c7cacebeb4a82= Ib67318fa6954ec8f3247927d34e74f8c + I9275bb36e58e0f17964e13ee7f027ab7;
            I1613ae89442495e703a52e65b8a0bf9f    = Ie964e5a463904ac52c4529ffb3ebaf65;

            Ic89597a95f50382cd3a2730896735d55= Ib67318fa6954ec8f3247927d34e74f8c + I1b6d20c64b9f23fb6c30f723546aa285;
            I6089da825af433e847c0b1bb9ff7d373    = Ia74858d5df6a76635e6ba60d0b1a63ea;

            Ibb7d203dfc75bf6211b09ab94877f93d= Ib67318fa6954ec8f3247927d34e74f8c + Ibb3d57d510cad00064a331f61f6400a2;
            I6aa7fccf4e225fa70063fd24dab74e6b    = Id9c69999bee621002fa9b387aa809dc5;

            Id2f2e6837c83973cb2173454433acb88= I8774ce3f11362915c4331d1026e452dd + I80f2e8f6743e28e86e4d85b295e2f768;
            Ibe2a5f680405f233256b6fd806b72ae5    = Ie9e8ae352a1699484f85ae1e7b7f9246;

            I1259d5918f8d65b4b22ccfef22fe3afa= I8774ce3f11362915c4331d1026e452dd + I9bc2d5692474b8368c570d92835191b3;
            I662d408ffd8fb9f249e531a167161429    = I5a006c73dcb7807d5943857199cc3535;

            Ib84e8c6e7fd9d7762e6e7e508d5ee40a= I8774ce3f11362915c4331d1026e452dd + I30080cc6c03bbe933165d266558a822c;
            Ie95b8a5c2da6c0877d49c646c194f5b7    = Idfb53869ea5692adddb6f7452d44effa;

            Ia032017912715abde99ffdf5ba732c5f= I8774ce3f11362915c4331d1026e452dd + I9485ae915474a31562ce358666d66245;
            If940f33461f5e297e158db54f6aad610    = I0d11a8980f8fd7aadc8e48e62a653aa6;

            I55c310bfefb635448ef9c25c5d15987e= I2392b2d17ffed6073875fbe8e92534cf + Ifd958901d2ea2284f506e04a058012fa;
            I54aa9d4c6333d94970eae97aeb3603fa    = Ib843721cd2106b7e5cc21812aeb374eb;

            I92c0f229cf7fdb2cc0fe4d84f4d9b11d= I2392b2d17ffed6073875fbe8e92534cf + I1070940dc2ef6e8ee3d1227ec9ff3162;
            Ib82fc62720e6346e1c05cc33d596447e    = I400d30374ae90fa066db0f5a29195e4e;

            I5570eb486d238fd96f9a59b174f5a22a= I2392b2d17ffed6073875fbe8e92534cf + Ia54b6f7044a831020e49f1bf48bc063a;
            I24873624848b61f313865e10e77e35c6    = I49316949f603c233556dfe520b9e1a61;

            If6f01d24acf4a8b38bdbb1b366cd9a47= I3a4f0d3e32596ef05477f494768d4266 + I7c0f872988488ac69815d288885dfd2f;
            Icc3915d8325c22fc172f731553798fef    = I57c335ac00303b6df3bb5bc5a1b1bcb6;

            Iff29fff36064aa4f9d339d4c62956e61= I3a4f0d3e32596ef05477f494768d4266 + Id2808e0f40992c79ead4da7c734e5b79;
            I93b9837e63103431a0fdaf319a465c90    = I177fce9af9d7a8e9e9dfe423c8abe225;

            I818d7cae6f1b80ac452dbfc073ccfe7a= I3a4f0d3e32596ef05477f494768d4266 + Ie71c7babb5d17378d40444b6bbd4e7a6;
            I91237af3aa2af551dbbc626bb701215e    = I335535f77c13df799b6e5f9613607a9b;

            I77ecfe991c6ec778495d7d5e5e442eca= Icd08ff59cf6be3ba97698dd55703339e + I75f9d3a41019dca3044a1c2cf7069662;
            Ib254d9701567f642d3586641edf85128    = Icbe54351ad1360193ea28dc76e073f23;

            Ie7c6a56e8b6f7756bb5a24bdfd6a855e= Icd08ff59cf6be3ba97698dd55703339e + I6e7e27bb176196e4493bf9c45ca19719;
            I25c50067a62d2b3599d15f12f89d384e    = I812a6ce8adb2ef9a2a9eb7e7e8cc96f1;

            I9f9bc8eb8b2978a3dc529c34516fdf75= Icd08ff59cf6be3ba97698dd55703339e + Ia0977b79857bdbf058535c30e338c38a;
            I238be7f0e4a209a6b4201a024c8aed82    = I87a99623e8305e331ca590dc62df5252;

            Ie3c0e5a4b00a92357a5d37e527d59b61= I985fb7ed22a8476ea322c9e3c2b3851c + I08e907b0619bec3ef2cf4cb3779e0794;
            I233f5ddadd45c0df2108ea6c1d634f3c    = I130df8a2e7e3e33055f2f2997e6d5716;

            I9b9a9486420e7d4aa105c48dd50aa74d= I985fb7ed22a8476ea322c9e3c2b3851c + I64c4bb0d40d80ec52aab61ce46954f43;
            I87a320ddaa1478146ff6e519dc65c40a    = I07ee1ac328d24e8fa9862659903fd379;

            Id12199a504f7aa298fffaaedd1aacc99= I985fb7ed22a8476ea322c9e3c2b3851c + I600ea1371a2be66430ac9534583b512b;
            Ibf03d6940c0a38bef038a28b6a7b625d    = Idd74d5e61d5397193aaf3cdb96dbc84b;

            I813691fd8ea36626d32c8d2562163f32= Ib985709316b1b0a9d3fa3c1eaf6c641f + I1391018fb93372ccc2fcc08700e38b65;
            I90942470e2057e50ce4f5745ed68b81c    = Id74f690142fb1e4a04fa3dca841979a6;

            I5fd3aaddc3eb8afeb82768b45e2d53d7= Ib985709316b1b0a9d3fa3c1eaf6c641f + I749b9c345f23aae03c595a2c76126ecb;
            I77fbc3f3b65962b610e39f4b085ecb7e    = I8327851510864c943e64c3d22b456152;

            I1ac281eab6c7459e835fe992142b7857= Ib985709316b1b0a9d3fa3c1eaf6c641f + Ie230ba3c73808e102eee9e5868595e7c;
            I701845efaf1b02aefa381d4f6b45c401    = I4f37cf4b922e288365376a45753c4a38;

            I49e5078c9161e8bee00fb76bc00b5288= Ib985709316b1b0a9d3fa3c1eaf6c641f + Ife5b9afdbb30c122b84d5378f9cb366d;
            Id446ddfd713c6e1592c562cfb123ea8b    = If50168d2535d752dd95301bfe723db9a;

            Ia697adf14616bf50d6e8178596b9fa7e= I4be898887dff6e2cebe53f135ece131b + I0982b8d7f99aceb8871c9c10448f54c5;
            If4f752779d27392e7536565d425bce25    = I6eb5641a21e34b4ced1cf124c3f23646;

            Iff3128a26dabe63b015dc6afc98a85a9= I4be898887dff6e2cebe53f135ece131b + I97e89a2ee18d2688d7c1a640318a1e0d;
            If112169057d6293326a56443ac3cf517    = I94da98c2f9e0c8be8ab8f23a2a10095b;

            Ifc04708ee5a7cc2b3f1850db778fa42e= I4be898887dff6e2cebe53f135ece131b + I94af4b6b9dc11935db54ba872889392d;
            I78f727f8d85b5d7f0ffa57f02538f939    = I339ec0bef37cb2e72e8e8795686da0c4;

            Ia405859c9dff67905b2e91bcbc06259e= I4be898887dff6e2cebe53f135ece131b + I27556d599dd1a27ee8f49e819ccbf29a;
            I01ec629f60c17c2251f977205234cd44    = If7c621d8183ce83092644a1d80d6c77b;

            I2fec8f62b28575e8f3af756db66fa232= I004db04f61fb57aba81e15cc015442b3 + I7362f08ed4e4ae309dfbfda112c56ad6;
            I23f774adb64807c0edaa9941c75651b6    = Icb4d6012447eb0d6bfa8e8b3f88f0ff9;

            I98e97c02477032ead66dc50f3f274e5a= I004db04f61fb57aba81e15cc015442b3 + I793ddbf6a5d026a57ab72984ca19deac;
            I2361ef4fd70e4c05b25289d0845564c4    = If7c3b54bc0cce4eecf8f55fcf4a5a588;

            I9f2dc5add3a4d1e6eb3116c741cd2f82= I004db04f61fb57aba81e15cc015442b3 + I3bdc5ba374f85dc61346e4868c41a6bf;
            Ic3067b434ca17be7bad595e1f9b822c5    = I1ffe02eedf41df8b947a285adc220fea;

            Ie122f7d8a48d7ad29d998b6a14b8e70f= I004db04f61fb57aba81e15cc015442b3 + Icce595233ce089eafcca3eae5e71e5f8;
            I3546ddbae9c9db4517802db56cee35f0    = Icd8c721f78cfbefbf25c2e094927401a;

            Ib5576c996062391f44066d893dd5cb91= I8f7e3dfb2f728d4cd1e79b82b62b0406 + I88aedd7f52399f5fd435c3415f2218ca;
            I35e91092ed503831ed818f36a1ce1537    = Ie139a6a80ab0051c5d951103b1554338;

            If931597aab866a74c3a3ffb1cd429583= I8f7e3dfb2f728d4cd1e79b82b62b0406 + Ibfe325e48511372569e0d98d9c4e70e3;
            I973f185cf29e13193abf0108d4faa9d1    = I993fd34b89fe9b0af3348cdd91ecf025;

            I79878bd69ed53785b8a5f025a2a00a4f= I8f7e3dfb2f728d4cd1e79b82b62b0406 + I28c3818247c7c6de11790f6692882b5a;
            Iee58b0442a6cccf0990ebb551b47fa92    = Ib5d321981c2997b3635fd0b342993d38;

            Iefb0a20652954fc2002154ea874c120a= I8f7e3dfb2f728d4cd1e79b82b62b0406 + Icc3cadf40c09be1a8c2847caf0e3e63c;
            I2cb3207a5c1b25386ac7eb532955f260    = If1660e858bdb3b0c8a4c1f93f4fe037a;

            I646ca66e4e9f24b4fb75b38bf293b4cc= I991054370345e61638ddaf81785505bd + Ie317bbd70b9092b840c0f2713204fb9d;
            Icd4f07bc30c66f7f5b431ed97e7ac7b6    = I7d9ab0daacce00542083a30a35297207;

            I051f0d4c44123e3637b84a32c9a00a75= I991054370345e61638ddaf81785505bd + I8922cc37cde6ba132f632743113e42af;
            Ifec6f3a1e10144acb320d5d502ed1ea3    = I9761f2282bcb9637892cf898b928126c;

            I1876f9ec3f6f637ee40cdad7cc347f6f= I991054370345e61638ddaf81785505bd + Ia3d129fd297905bee180293c0c39d9ef;
            Ic87bff64a597e6d02583041b552328ee    = I25de2ab105b6cdb0e30ca97822109fbd;

            Ic3d6b8dbec6cf92a9b6a17fb2f75dcd4= I991054370345e61638ddaf81785505bd + Ib43886d923b8c683004713ff25b2f90d;
            I489f21ef8243ef8caa1c29f034c3e2ac    = I23c14408deedeecba4753f182549adf7;

            I7d89f1db7b1015d34363ad781374de58= Ifa1f503965270d10e7a5c9a15576069b + I3521b10b97b0e74888ce385cfc772945;
            I773901563077961acada85962209d68a    = Id208387ab734f8ccfaf1567e6b00a4a6;

            Ife217ec4da1f1477bce034cb3545160f= Ifa1f503965270d10e7a5c9a15576069b + Icb2b390266bff241a688961136db0f51;
            Ifbd176fe3e78bc2dc2e0e77ba3ccd2d0    = I54e43b8da49648867403cf839e87a9ec;

            Idc5e5e98508c94b87a760f8eb36fad41= Ifa1f503965270d10e7a5c9a15576069b + I8bf8b0cf27a2654a0e7fdf3255945b67;
            I53f68a4cb81c71ee7bd6f61171b7478d    = I66c8b8649e7997b7e4c9c17f7c0b17b7;

            I9e72b0c823f297535f13a1b3072c2776= Ifa1f503965270d10e7a5c9a15576069b + I132d9671c582876568c0f7f5335f5227;
            I7568ec59f1359bedce86dbc6af50df71    = I9a0093065fb4cf517f1e7b75b3080b1c;

            Ia81da7c58d6636ab70e0cf3e263a12c0= I24f773842a4742fb58d09cae45717b2f + I820fa56328e3919970dd64adb1d4d8e7;
            Id2bf82d6bf0a201f80a58357038a0992    = I72d18b26784448b5514e66251bb19ebd;

            Ibfc69ef08382c79e30cfafd89bfeff69= I24f773842a4742fb58d09cae45717b2f + I4cff1804df738cbf4f940c775236df9c;
            I22442354ca2b77306f25839ce6124699    = Icec022a0de167257d08e0b2beb6ba8f5;

            I2d2afa9165b7121dc8289e9e6cdab5de= I24f773842a4742fb58d09cae45717b2f + I450c0d6ad5d3b1f18bb28e3a432b5442;
            I71a5c2876a07d8edd001ef2d108e59c1    = I3d8a7850f0080b0d6068d58837e3294f;

            I065052693fd8ca87614feb60f7ef37c3= I24f773842a4742fb58d09cae45717b2f + I0859c80b42a8c60dade8f05d58ee3701;
            Iaf333aa6b135927cf1ad1f76298ccd63    = I26b947511e25e51f1bb9728c169e7e64;

            I13344a81551374f665cbc17c7e94296a= I5bac7e0d778a547a0ae764fe259b6f7a + I68e5b12792a86dda0576742831d3b728;
            Ia71cfd8cf9bea4e600ea204e41271c7d    = I8baf26027cc707ae93b6c74e2af5f207;

            If5a1d2de0715fa87d191ee5f48171676= I5bac7e0d778a547a0ae764fe259b6f7a + I512f57a40c7c8cb2f040bdde73e44ca3;
            I164b032929ac2b8cf1a6672859639a30    = I9902253554855a3d12ceaf47f6cc5569;

            I02b256f74ee86b42ff1eba5e3d242737= I5bac7e0d778a547a0ae764fe259b6f7a + I58447d6ae49a6be2d043477a06f83df0;
            I2ef0447f5c64fd5c65e23c16069a62ef    = I81ab0ce0526dd851c51d5d42f807e62d;

            Ic113fc051eefaef846f440e98f2f8913= I5bac7e0d778a547a0ae764fe259b6f7a + Ib3690ec149adde94343d3e617931a287;
            Ide7008ee7f1fba156dc6145b3505e553    = I51dc4acb242b33bb123f8b106aafbc93;

            Iabeab9bdd0bd82dd145218b563b5dac1= I255577ebee6768871df0224fc1db2db3 + I6c661048307c23c699d4b3636564de0f;
            I129a7ced6bc6f48f20fa552e2519925c    = I32ca8b2806bf397557167b133d1411ab;

            If9ce0a09e3a4e816dda002a24319ac0b= I255577ebee6768871df0224fc1db2db3 + I557ef77ce931535467a07a8d70145f55;
            I67123cf825352e52cf0158060ad69a13    = I5c39fac168568808f33fc6be5eec66a7;

            Ib5a7d72c36e41754033a64fbe0718784= I255577ebee6768871df0224fc1db2db3 + I41f2bf9ff00f983ad1298c8c83b041cb;
            I09923d784a9f9625a37221f639537941    = If355236b8b8375ad095cc46a373ad4d6;

            I41df12c7dee8526abf92b8e98965fa06= Ia7fb4af3d3529a32f902a52cf5598474 + I8be4be8471625db0749e6385f87d2dcc;
            I5947be93fdb18bf0ad341fb826c9e6d7    = I31fad95729e24c7724a73285e966684f;

            I83dfbd224e7465a6fd769e407182829a= Ia7fb4af3d3529a32f902a52cf5598474 + Ib451127b69a0a800332a712af77c6d29;
            I08621ee033cd49702ad08af4d31eb999    = I0415d9d3687656d7a07ea2c12ba505d1;

            Ie57bba5092ec318456365b81b36aaa65= Ia7fb4af3d3529a32f902a52cf5598474 + Ib5414585cd6976cfce42e42190cc08d7;
            Id5eca60b22d3835119571fe4b1a03479    = Id54f584cdc590112180e9000e1d015a1;

            Ibcf043d24474ab8c1002d15fde2d7da2= I2c98806141f064c9e92935b23a84ede1 + I7651176b0a74846108fbaabc5cc4900a;
            I7267ba2b9cb511a48a3a7044e854f7da    = If9930e999d72a139c345aeb1c33e51c1;

            I2e3385871c6ed8cf9519f273c8a19fda= I2c98806141f064c9e92935b23a84ede1 + Ie1e9326e4eee006ec07abb6bb7d269a5;
            I5893fa21ec8bbdcea9677cc12fc4057a    = I28e9624edb8f59290eba51c87f2a88cc;

            I664917b9f44515bf556d69ade4ca408c= I2c98806141f064c9e92935b23a84ede1 + I1ca59325ff30db83df5bf0a2cd9706b6;
            I564896fe01ec799a0fbe790473753559    = Ie6c99d8fe1a105832500bf8a722c82c7;

            I28deacdec0fbd0bce49b654c2620ac38= I5680847bc8d224fa4ed93b2fc0d841e1 + I8fd26d47ecd4cdd08294cf6133468d17;
            If279ab7c515c4039c8272b913c2fa107    = I24307c47884babba3b0a16a1791c674f;

            Ibdfc4852c620f573f929584e6b816f35= I5680847bc8d224fa4ed93b2fc0d841e1 + I38e2dbba093928b874d447362d89b291;
            Ib61705ff5820f531eb17c40ed05f6ec3    = I2951bad4b57a2ad6715844998c491ec7;

            I5a69b2bbb63ab919ea2270503cd326f1= I5680847bc8d224fa4ed93b2fc0d841e1 + Ie2f5b03f3b136e651b8aba92a30d298a;
            I50149e5de41ca2998c4e8cc4b19e166b    = Ie0149abcf22aeff58be4cb418f477239;

            I2eccd8d60a19481fa595566f51c7aa4e= I365254279ebb10dd7ba0b3482d5e34cd + I0c1e22375d5e023c24519901b92eceb5;
            Id40cac3272643f3f91b73c6aa1740f3b    = If8ec8dc5888438922c6074ff23eb42c7;

            I49eb4bba42440657fe04b711eedfa67f= I365254279ebb10dd7ba0b3482d5e34cd + Idd1b6014de2f053554ed09c29bf3e640;
            Ic63eee2d700493c41ee2d186ff7111b9    = If969c721b9636b840193a85d8946fc32;

            I9ed8323951af0de78ae89153cbf9e9eb= I365254279ebb10dd7ba0b3482d5e34cd + I97f2813ec39bbf1513faf66b3e38838a;
            I51de42598e0df4a76cf7b02c61ae9550    = Id6dec5f563e485414043770af559ec76;

            I1d00816529836546b514f54b1275d39e= I365254279ebb10dd7ba0b3482d5e34cd + I0a3323aac825506435068f6746aee974;
            Ia89a1a58f6327ee3c105cae860942171    = I79ae237d2105b50c92b8507272bcbd4e;

            Icc58b9a24fb9ef7e8fa5f13a2cc0a0cb= I365254279ebb10dd7ba0b3482d5e34cd + I312ce79a8dd2ce3d37c930d42640509b;
            Ib149a5872e31cd5df77b66298b4aad12    = I9ea4ebd1f6cea81da598f16b5a7c31f4;

            I9339aef608b029175b488e82f5b3f1bb= I57bf4ad773cc058ae1bb7b1911dc3174 + Id60cbf534604e5dba988050ef5abe625;
            Iaa16c14572ad0442eb3c58a97bef5ada    = Id7b8f8df1818623e7a9e897e019a09e7;

            Ibd2f24860b701ab46e0c436d774e43f9= I57bf4ad773cc058ae1bb7b1911dc3174 + I40e99289d5762e77a3766eb8251eef00;
            I88d5d48e05b1c9a6d8060f58917e3834    = Ia5e1a46c7d21e79ef859b788b27ee3d1;

            I37fe66ec8927f27f646b304500400ccf= I57bf4ad773cc058ae1bb7b1911dc3174 + I9e09c25be9f877c1e1aaf79bf12c7943;
            I4269e18c2df4d39c683ffb7d01a08322    = If5b0270fa354f64b8b58e5f02353daa4;

            I4bd6a48f494cf633a857b8ccbd67af68= I57bf4ad773cc058ae1bb7b1911dc3174 + I30253dc91301ca27b5732312c01145e0;
            Ia29017fa9327fdaa7c10b2797f8aa6ec    = Ie800c32198a9d6181225f2274b301d9d;

            Icd7a7566438dc67e77f138ac814844f0= I57bf4ad773cc058ae1bb7b1911dc3174 + I467d5e2554ef25873e0b44e947ee0011;
            Ia142ac799256541fe33f898a6a31dd71    = Id596782860b623f79a8fd0e83712d9d0;

            Ic3d4239413333883dd926c7a42c0a87f= I57072dfb29c4a3d2e2b40e46e62f0d95 + Ia66c399023e500ed67197dcf236f5d42;
            I4c039794243933a9bb7ad6db7eda6a87    = If5a41054200c97e01b9132f7c7ff9793;

            Ib8298d1ead61bc00eb31599b3087d769= I57072dfb29c4a3d2e2b40e46e62f0d95 + Ic66af6c3c0268cfb0e9f0776c4f4e961;
            I0debb3ed4f9540c162cd525588e0ae3f    = I2cf304c8f8efef74593929b1bea0bf91;

            I23dbe33ce46f94d3dff1e6d391305609= I57072dfb29c4a3d2e2b40e46e62f0d95 + Icaae0fb0f460f68d690ab00697355a49;
            I681eed68ee814fb18fd794207d9266e1    = Id0b597aa1dc456b83d4e38147c97a9fb;

            I138286817f424c76e8a4f30540b0530b= I57072dfb29c4a3d2e2b40e46e62f0d95 + I0d66aa55747362354aa81d96057bc4c2;
            Ic260784b8910f5a0483afee9b68efb31    = I318a691d3ffd634a1c5c362d5b3a8c34;

            I30c645a78b900306864a1ab23e923bde= I57072dfb29c4a3d2e2b40e46e62f0d95 + Ice73b514709469fd21cd254bf4ceadd9;
            I22cd2d30a7684002cacca4deae4c95a0    = I881c34f97e2d2f4765cf3cd7cde53c7f;

            Id88681d0fe3ea62530166938503db05a= Id8cafb6f76321bdaba9711133be7be99 + I54cfd68212d97a2cc8241ef429429453;
            I136b4136d582f9fad21f90297cfafea3    = I922d1ac78df6c82308d2028527f8f56c;

            I808008402174fa4edf42783135c0c3a9= Id8cafb6f76321bdaba9711133be7be99 + If8aa3ec1b5a4a3c122da82467be917da;
            Id8d6be9677d3b0ceca26b3b671757c2c    = I49dbef91e0572ad9296838e769edf0c3;

            I3ad4d02ea2e52a49b6fa4f1da9b58149= Id8cafb6f76321bdaba9711133be7be99 + I53309409a6059c3bd39f037c23ec3458;
            I6a93f928c104ea211dcc8a461506327d    = I8819e4519e4930d300f5536af5d62a94;

            I39486eecb7bbfecf26573a7a5876feb9= Id8cafb6f76321bdaba9711133be7be99 + I7e28234bdf66ab5489d36d15678db797;
            I240da147648bec33195a5f5c273fc6f4    = I4779a6c85288e6dba977cedd1cd3cb6b;

            I21e8ea20029fb2cb62103405b81b21b0= Id8cafb6f76321bdaba9711133be7be99 + I45ba06a6d6f00c174b1439a6f226a085;
            I55494d0e8454e3cbb4158559e0d29984    = I934d36f3afd37afdaad46c93f45a044c;

            Id0b67fa451e276889e02779ddb667904= I6344e71ca2b0fd39d36caedd889c3085 + I786dfcaa131b99c254aaff15bd2c2b6d;
            Ied3cc579b3cf126081acf8e1117007cf    = I2667428380ad21221430252aa00402bf;

            Ic328d25a58ec4559b753da3bcff938de= I6344e71ca2b0fd39d36caedd889c3085 + Idad14b6383b9af54eb35e72ff3d10035;
            I76140bdc374dd6031097575fd231b468    = I257185648f29565e2259890a6a70583a;

            I49c44c2f2522e086c2db8a00647ba35c= I6344e71ca2b0fd39d36caedd889c3085 + Ic8a272f82736fd599fb3250e970edf9b;
            I650345d21e5c2e7a9bf1810630161089    = I49a61c916eb52d0bfd08700d087d379a;

            Id4152a04385391294f4b8a18df2cb9ee= I0c99a68e0bed90afce18807acf7d55bb + I3d6a685a1913bd8be01fddbce1edec2e;
            Ie852635f073dc918e7b1075ffad46f24    = If180a1b31f53c672e4f05b2aeca3caba;

            I5b0213a3df61e94fd0b744a8141f7502= I0c99a68e0bed90afce18807acf7d55bb + I8c0069e8756bcff203ce21ae3170aa42;
            I9ec80c14eb5f0f305e1a9e6107a6001e    = I335057378d9ae46b1e1442fd341fabad;

            If0ad11ed403cbbed68614b01e2a3793e= I0c99a68e0bed90afce18807acf7d55bb + I5b9710b16effc8bf0695517c6e651836;
            I80ba56447ab19b33610c23105b0b1637    = I3027f4cba09ab3eee29cf9b34ed27ae4;

            Icfa1170bc73534bee13778bc3b88a2f7= I1c95650979c86310ae2a949961c9db11 + I57ac487adc18165136e9b3c7c50f95ad;
            Ib9132d9fa7180c3fcbacb7c570d6b0f2    = I9ac1c5487994b853d666af93d35c82cc;

            Ife1bd938a0dd06d8d3cf30ff41a303b2= I1c95650979c86310ae2a949961c9db11 + Ib484aa64b795f7e36198b800f302164f;
            I01621f113f636a9caf9b5ca0bb20ef77    = I099f1e1b4eb55718dd73dff7efc16ae9;

            I4a09cb1b99b476fa6fae0bc44c41a041= I1c95650979c86310ae2a949961c9db11 + I038b42a83025f5eaebf45799d1ebe7b0;
            I3eeddb549c6e1f07469c0e0dca68be92    = Ie9ebb06f41fbc042867ee14d8f4090f2;

            Ie08cf323944813e4b9e2d59a680ffe8d= I04eaefa5d133e53494fc270b07be7043 + I7097c9518bb3351818b96f31ed49c6d3;
            Ibe664dd203ed4162abcd36eb8d57bfa6    = I2647305e100a9fb38fbf290f12778d49;

            I85fc307fb52d58550eeecd33bc4207a4= I04eaefa5d133e53494fc270b07be7043 + I41af7e4c97fc04154fe6de66b82499f5;
            Ia66176893fe306ecfb415d948c50486d    = Iae4b5e5348101abc4640c84686ddad69;

            Id00dd13741fe621d0a240bdc92318f55= I04eaefa5d133e53494fc270b07be7043 + I73ddd7cf9272ceab5a663e2244e72d7e;
            I8bd4210dcbfc1956381b460fd9ef789b    = Ibeba1d51f76197f960672ea90dabfb75;

            Idc8e891fd432df75a4eb133ce35ecec4= I4a64fa2412eb8058c2dfd9351d7b297d + I2f9e56d570e72714a06c59aa9e4334c0;
            I1ba6328ea9cb7cebcce47d5407d0eae7    = I83ebb6a41c9d866a8ff3fe3fa0b5321f;

            I2a51cada20cbd14f7d5a289599e68b53= I4a64fa2412eb8058c2dfd9351d7b297d + Ida5b16851dc06534844a0b037d74feb3;
            I9e79c17bd782bb7981b4a3623baf96a1    = Iedc551659ac328435c906b5748c9790f;

            I65a701d1e083e501544bb0fce24f0c4e= I4a64fa2412eb8058c2dfd9351d7b297d + Ia48f0029e9e76386f3dd70aacd9adbfa;
            I7c6f64d73ff9c6e7f2ed69713e056a2b    = I95e1540f2a2eadf6fb80e3519a1d9d5c;

            If3020a9109ac83274b5bafac18d176de= I4a64fa2412eb8058c2dfd9351d7b297d + I16507fab8f9076bfeb419896fa7cdc1d;
            I00b962a9bf04b62244591051d2dfdbbd    = I3587e6334c7c3f23bee5675353bbeaba;

            Iaa6bd55038c2ae911e4df08f707c55f5= Ie8bb2fcb752c6a33254963d1ebb4130d + I58f0b81a46549cab8e74ecbc285df23a;
            I3a660b57588325989319701026f658e6    = I4e71cbc9773ff4abc24804d39a64abf8;

            Id49065cedf20e13abac8971534bb8b0e= Ie8bb2fcb752c6a33254963d1ebb4130d + I37998a91d20db2248ebdd8e661d42f70;
            Ibae27cccf3f64e8653c1e244e940e421    = I884dc79c03a585814e9d058ef7669ed8;

            I0bb64952d77b59803a561e14b950b9b1= Ie8bb2fcb752c6a33254963d1ebb4130d + Ib4695d4389db72c5ac7e31809072c290;
            I27b89a5001312b2aa48fe385d8a52063    = I0b2b9b8f1d6c6d5c6c5a8bd883d3ea5c;

            I01e295a6ab88c6f34b44efcc32a23233= Ie8bb2fcb752c6a33254963d1ebb4130d + I3dd1f28cf199299aba54e47a429c9b11;
            Ic6a7476db711a812d146331c562ca7c9    = I645a63009d5be827b30fa02df646c872;

            I2acf864d587b7681ca0fb6e2e2bea617= Iac05b7e3ae18f948b72c356ccfb8000f + I05eadf11cdc6c2f2b021e33f2438fa49;
            I01ca07fe91b5f1edf87300b3583e77c5    = If4630c847d9890c2b93acbaa6c9bd392;

            Idfd0410b37713e8808f8bea81e2af881= Iac05b7e3ae18f948b72c356ccfb8000f + I1171dc208d5db1024dc3f09a90c78ca0;
            I6da707fd74249175d1f68dccb66390c0    = I49c56ae29a27e764325a9dcacb99f907;

            I02861f333b5adfd4962356cdf5a11f23= Iac05b7e3ae18f948b72c356ccfb8000f + I3d601db540da359ae4d22f960d3d5af8;
            I0ae62aae426b75b06d95c46baf33f08e    = Ie5272faa6aabb6e8d0720cdb7ec98358;

            I4ddbc3daa65b111cb0d45e13d62cc292= Iac05b7e3ae18f948b72c356ccfb8000f + I49d9203dc6f8c17f17383e8f7e01f005;
            Iec512b5870f295a50921e7e0289a7d35    = I92779ca466dbced9070a774d84439921;

            Id363d158feb8fec19b5f3d73d84f0068= I27da3f75cca6c49e55db90306aa68e94 + I72db05084d30d7c59ba1cb06d3b09400;
            I3aac84acd9d78070472b1cbc745c80a7    = I037e8ab38d779544d25ca5a4bfadeade;

            I8ec9b7a6e65e727abbed336ce240a4cf= I27da3f75cca6c49e55db90306aa68e94 + I8d4e3962525c424786ae822a6981a5e6;
            Ibbb900f56de318bf6e65b49791835ef4    = I3001e26d13b0cca9bc53d24324ac44d4;

            I128fa1e99b7eb9b6905c2cfd26b95ab4= I27da3f75cca6c49e55db90306aa68e94 + Ica4ec1647bdb5a3aad6db6b447bd7995;
            I2c2ac1e722fba72c759f1d37b88a9a10    = I933465899e56523ce1c470cad8dbd229;

            I93d459b6da42a205c91c48622f0c5032= I27da3f75cca6c49e55db90306aa68e94 + Ibeec86c75d950ee00dd63a2930f08a24;
            Ida0a18f1b79aff4ddf0e8f7e27794674    = Id8b135f08d0464f9e308e25b8df2eb1d;

            I1243cc8d5dddf7dd65b40c0b3b958b9e= Idc7fed723190098341225fe01ba65ced + Ic95668328a2121027436f682bac50b9c;
            I9f2029db42c5a968b370587c958c8929    = I938596dee81ba14870ee4acfabce5e7b;

            I238df7e09d42bc93a972da349a00f511= Idc7fed723190098341225fe01ba65ced + I82a14e1ee4723e7d9a13c1f2b8b13691;
            If5755f4f61a89d91a91188c17ff5dc5a    = I61599f00ae7d6964dd40c96edefd6f67;

            Ic658b2afdc7331653fc84d6372d47418= Idc7fed723190098341225fe01ba65ced + I47b2438c3680b2d816168df37d7c491c;
            I4419d97c3174ee4610eb6ee9c06cb256    = Ic847a85de8e8ba2df520b737ea004374;

            If39be111eb101c9c983fe0baa9a1cb18= Ife9065805598960919ee4f14c3cc6fd4 + Id683d693cd50645c3d6d657aa1c8bdb2;
            Ia964f83676273055e20a2f63c8fffa0d    = Ifb0f088bf5bbf1884e1f27ed9808c273;

            I9d19d5b7d8b256c1707de97a4549c458= Ife9065805598960919ee4f14c3cc6fd4 + I461398638cb8280f1779915298540b00;
            Iab4fbc811e87df1d1f5821ea732b6a93    = I8705aa11e5ada7ec6e5431292d83fc54;

            I6c2fffe204091f7f64aea16b0ac98769= Ife9065805598960919ee4f14c3cc6fd4 + I5983bf2c6c90b872ee6cf58b5e520311;
            I4fbefbb10724b0844c95e85495d4a87f    = Ieaa7babedd5bfa1c8e1eb50d62ad9682;

            Ic4ba4d2e5c12d9f1dd233d64929f1072= I717c5c2d6a2be61593492ae5f17a112f + I2b49d74cb130542f2ca99534e2c513b1;
            I717217d0b5a526f04c7f5ab0835dd5c7    = I9eb9f7a6fe5932b574084bb18ce44e78;

            Ia9dec5831998d472d11429e5a7e60ed8= I717c5c2d6a2be61593492ae5f17a112f + Idbea892c8109117f90b453efe8ae25af;
            I235937b643e8f2848116dc76c43f47a7    = Ic4b80e5673ad931188a2edfa1119e139;

            Ieaaf52c1e663f260292bc1529718d681= I717c5c2d6a2be61593492ae5f17a112f + I6745cacecb7ee86cf3c7ad7eeee6048f;
            I7481f17d659cce5b4c72a68a9f6be67f    = I5cdaf1ff24d7fb2bb4411b63a0a4488a;

            I37061896a09588a73445deed73d3746c= I4c31fa8e6eb648439cdae1de1afe0d6f + Ifd77e040c5f82790b1d5636a42fca602;
            I5715c21c80992a61bff8aabc3f80415b    = I7db6dcc03117fef703f20919a3c2ee89;

            I02f25b80945b6f58193fb37add3da2d8= I4c31fa8e6eb648439cdae1de1afe0d6f + I28aa517220bf597cf898660f698ef19d;
            I434e3216a615eb46be5c26ef914b9cd2    = I3d2a8a166ccade50e320baaa68b40954;

            I19045602bb77f12666ebd44f813db2c5= I4c31fa8e6eb648439cdae1de1afe0d6f + Ib9672d20643d856ff31905ab14c0ac87;
            I918326ac0a744d234d74e2c08cf41eb4    = I3356737fddf6440f36fde442d29bb860;

            I4abdc8d5318d2922696a8aaee46ffa59= Iead549a9af27f1fced7d9c36e7b5c3f5 + Ic28b148967a5b3d05409976fa9001ac8;
            I966706d314f4c0a7ec842dd699d34926    = I13d6fc4a99a3a9989e655c417552fdb1;

            Ie139f2048f346d82623c8fc6d40c9acc= Iead549a9af27f1fced7d9c36e7b5c3f5 + Ie81315a3a14a5ef879d8e3f405936365;
            I5a7d246d88ef12e999f4bdee40e5a585    = I8a508ec5f2c2aaa05b632f422e67394f;

            I8d99c96e203fafc81d13ce5aee925d75= Iead549a9af27f1fced7d9c36e7b5c3f5 + Ia605d14205926b3edc6d1c2f69f70ac0;
            Ic2dfaf65c4e17a8dcd55f766c314d6ef    = I451fd82336efc778a51debf10f7cf325;

            I37b0bdeb3cc54d6a97720c4912c67832= Iead549a9af27f1fced7d9c36e7b5c3f5 + Id555c88cf7f0904db74d45cc75c8f5d6;
            I151831ba6bd0e162275c84815e3c0f12    = I76637de9be7c2c0dd0c324b4327a6184;

            I08257e9e6c74c60448e22fb9855f0825= Iead549a9af27f1fced7d9c36e7b5c3f5 + Ib9dfea1f34a120eda30d5bd919365a6a;
            I5a8f1675234ebed14d719344b530bbd7    = I6e6d24ccb985ade6f058ce459592dfb0;

            I32188cca2fc715698fc05b0fc6506434= I10422eb79364e7d0e21e1643d9060331 + I1a5f22b4e326d1684c0a8c7a7e754ab4;
            I95dce76a8d0e729d40fb3f573cfc06ad    = If379a7696fdd0afebcb8ca169bb8f34a;

            I88f1cbab9b8fa3802345f745d024931c= I10422eb79364e7d0e21e1643d9060331 + I2c1f2476efe593829ade470fe8ec2526;
            I6c26c7918254426c18f2e747c91438c5    = Idbd1062a6090858034185f1d5d503adf;

            Idf548c0e78bd221bf9f612f27002fae0= I10422eb79364e7d0e21e1643d9060331 + I8daf79a0a2ee1bac7f055af441539fa4;
            I0414ead2472e42da8a271cb0bd1debf4    = Iea3c638b692d2540c1c8c81a6308673d;

            Iedfd2e04f5740d283388639dde3ecdb5= I10422eb79364e7d0e21e1643d9060331 + I63f82f075d53205b5b556c0054f1a0b8;
            Ic6a6f5090470a76ddb7315c022ddc104    = Icd9e1d048d56d5d8557f80329bc6ffcc;

            I7088c83eacff6f1dfb134f79d469c8f1= I10422eb79364e7d0e21e1643d9060331 + Ia7bf82c9e5ca4467b5e50beeaeb975e9;
            I2a00ee56a5aa639f45eb3b1bdcffe81c    = I6f0de2d570fa0245666c834b823e545b;

            I6f8431671331f4ca7ea19656e0677cd4= I914cb87eba8baa40cd515334e59f26b2 + Iac3cb5b4481687fcf430c8bf52cfb74d;
            Ibceb2b824cd4bc10bb06ee8adc693bd1    = Ief41e2502056d029a0c8bea8c052700c;

            I1e31259e267e04920cbbd16bd7aa18bc= I914cb87eba8baa40cd515334e59f26b2 + Ia17295aec0a40c2b46a595dacfede2d5;
            Ia8b9f373fe68ac4cbca35e04376e3cca    = I7cd5df0d2845c7ed9f336a7940c7256e;

            If54d9f8088e67e44cfa3026f5a520fd7= I914cb87eba8baa40cd515334e59f26b2 + I0d96336eb4d5071d7e1d350e86513b25;
            I5d1a89e85f6609b469e73e15aeffcbc4    = I5471bcc8bf4f4d0fab46d549b43113ef;

            I6fd2c0746407b23aec5dff1e083f5fca= I914cb87eba8baa40cd515334e59f26b2 + I2587a5800a5a9ffeabc4dca503e3d964;
            I677fe06bad241bc8dd6a65a97f6db520    = I599b8e0677efc1541283c2d7bf84809f;

            Ib2147a19b44d361da628a628fbfaa988= I914cb87eba8baa40cd515334e59f26b2 + I327c9acb8934729b4ea5486787afa2e8;
            If3c0f892fd71eb0ed8d1f70b4b33450b    = I4e4829b24a42e96e5c8399156aa61786;

            Ie804d1f4b241a2de3e9d9c7c876d914a= I32ed679af4ab759901aee43c9d93eb67 + Ib65ff82aff398f6ff7ba711a36f41ee4;
            Ic65f0f75f56bf85122a89cdf07e98152    = I1cda8d902f71f780775c85f38f9e799e;

            I6cd1e6db57e06d8f5e60a31f48ae4809= I32ed679af4ab759901aee43c9d93eb67 + Ic2b20168744fafbe15037ed7fa83da72;
            I41d22bafaf58e4a6de04640864653a16    = Ic0b2c3e49d55853bc705021e5c0a2b06;

            I3e0e8832d5338423284ac4b2a0c5f3f5= I32ed679af4ab759901aee43c9d93eb67 + I20beb3fdbe91936f74a200cd8ec9817b;
            I06a46b86f6edede0f5f72658a19910b7    = I6235ba2f129cfbcff36b368a39312bd7;

            I6ac006d79e95e222cdc66754b67a08ed= I32ed679af4ab759901aee43c9d93eb67 + I83292bcda4645233d8e8a1dfe8e5f60b;
            I8591d0399594adacfeb006c5195c2c71    = I6804a691f5de298ab553ee66c3e9610c;

            I29087dda1a527842aeb3d35d66c853cb= I32ed679af4ab759901aee43c9d93eb67 + Ieddef08050c38d07e5d38f5bb7b099c0;
            Id90588b5f82cd32e801fbea04d24e4a5    = I973825f628679f8bbaf0650136e7259b;

            Ia67e5920bbac700dfee52cd96b15963e= Id376dfa5141402f4d41a8858180ed87e + I5b53fd45210b92703cb10d583f471ab9;
            Ib642d757fae818cd6d713ffb6ce18fc1    = Ibfa3babbd7909dfada58a7f579281b8c;

            I1f6ecd894d90547f661e7a3888d048bb= Id376dfa5141402f4d41a8858180ed87e + I74b3c9dd3a8168aacd4369b9ff68fdfd;
            Id76bff2a12cf792e52ccc463647334c0    = I0aa6569579526ac14e0d55caa4cef2a7;

            I3112e793c6e79e1f5da2776e69a34e3c= Id376dfa5141402f4d41a8858180ed87e + I39f9e8430db114991bfb27cc46ef3e39;
            I92ffa890ed6d83d4fc543504e4d421c1    = I87c99b1e08ca19dea7ffbfa15ecc2db9;

            I79152f32b45ed5b4a5302f6460707b01= I98a384bc62ee03f5ad7df20ef2d9af95 + I7095040b38bf9d6b5229c11d2a0d7c57;
            Ifc4a65edeaf630b3d29437bcd6c20121    = I40ba1533f32b981c4e937b2e48f38ea0;

            I3d16e7d6b190639b88a217f19ac63233= I98a384bc62ee03f5ad7df20ef2d9af95 + Ibec442c099da091afcf75a7c970bf8ea;
            Id57a11f56fc223501a9b68b8b05ebd3e    = I83483243e11dd867b1eea10b6ef0dbd2;

            Ia1be780c686163cea54b62d6ede72dc6= I98a384bc62ee03f5ad7df20ef2d9af95 + I56aa548618a4a15e9a35e04f5eeb823f;
            I522ba8bfc1949337e8befe82cc1e86e6    = I8265d9994495dbe871b565be6710b428;

            Ic398c31a2a6ca89d0236534589a5919b= Icfed259ca2bb2732d8e0c26ef67cd4cf + I2c487770d606451440eecf358202db32;
            I7153e27c44ebbc2f04e9ba03cf09b5e1    = I3d4ee0ad8461c2ac5128adc9c231f465;

            Ie91c3202bc957b350d1915000564392f= Icfed259ca2bb2732d8e0c26ef67cd4cf + I143f5e324716a94d24ada126886bf895;
            Id15e4b4f186ec863f12a54acd8ef8963    = Ib609900664dc10ef97873cccb161c320;

            I687957f5300b0d4f50d6893cc556bf25= Icfed259ca2bb2732d8e0c26ef67cd4cf + I1908897b529ca04df7e7da395be4a8ce;
            I95c77eec7575cd7aa93a36f31ea635a2    = If8b44d90a4ef1715e9144255d606a27e;

            I7816b368e8e8b8dd69383b2c9327120d= I20861535c450d6e6bf11c45dac120454 + Ib1f1aef6c0a9291553b62fd555feb2e7;
            I3c8114dbe0658cc2889c787f1366abfa    = I06715db3159c94a5913c05e9827cddd1;

            I5f021f4a664205afbe0761af4c8914f1= I20861535c450d6e6bf11c45dac120454 + I1ea33707e40a2e41513fdb3118371437;
            Ieacf971e9e10fb73c7df9f1da8372f30    = Ia295ba836438cd4e7c1b03b4261949ed;

            I69728004b59b5206a03a8e2087834f7d= I20861535c450d6e6bf11c45dac120454 + Ib2bbd59cd6098608ed53ac556036534f;
            I35de1b03ea865f2c6381ce73e03dc220    = I5f9c502cdffe77bb7e298a9bfdd325b1;

            Ibbe1d623f8f5f3aa7fc70197acc6df5e= I013929385ad819ddfcfcc59c22902ee3 + I118726375ca9381e45f001965fcefc5b;
            Idec12e02904ea98c7580919584f2dba1    = I3f13e4887f4982583fe615807c42d121;

            I4cb9f74288811592fd97fdff52bd6fe7= I013929385ad819ddfcfcc59c22902ee3 + Ia7520053a7c4a94437c6a780b03a28a5;
            Ia370c83631a2c1bbf39c7264deafafb5    = Ie1a491c10dad8dfd4b0fe42977d625b6;

            Ibb471dbccd39d41e951e98348812e343= I013929385ad819ddfcfcc59c22902ee3 + I42455e7e4d0c63f97702d204d18a446e;
            I05b4a07dfc0d2695eae34bea4c1c6565    = Id2334d193c70ad43e5b7cdcd923e364a;

            I7f37d68f8ddcf8b4d5e99fb51eada873= I013929385ad819ddfcfcc59c22902ee3 + If004552b2047ab1cf23bb50375460b01;
            If1ecdc27e3419dd1434e403f237c2b58    = I621999a98b66cc50cf7732668af444e0;

            I72ded7153883418a712ef967439d2159= I34fffcb07fe82f11fe142f7c37f39155 + I88bd8012c93dd9e2ed52ea5e9b8b0004;
            I039c552777d0fb40bebcdd2d4a3394c2    = I8c5fe32c1860a2beb9c14634c62a95aa;

            Ie071e08299bff6bbdbe1f84703aaec08= I34fffcb07fe82f11fe142f7c37f39155 + I7e685b06df8a8c2ac351fa9f9b76a81d;
            Iaa52fb63184514b6d754bcc896235150    = I5cc33aeefc2bbf0d777b4b59bcba7ec4;

            I1b79aa38a39ccfc839260af89aa78e7a= I34fffcb07fe82f11fe142f7c37f39155 + I2603e0b8b93f6680e44c9c8883f6512c;
            Ied9781e625c1fa8741853dd6b8b3a9e7    = I5a2f74df4050f2898061471586f3fb63;

            I7384296e4190d83fb9d9a92cf965125b= I34fffcb07fe82f11fe142f7c37f39155 + If97092e1e2147de199c94a23831cf6b9;
            I767272262e9d2e85dba1aa93f578f25c    = I54c68d66f2692522fdd982a31ff0b3a8;

            Ie03034ce6233ca24effe53a2c0c8f6f3= I61ca60fde05ed88cce714dcd8c13b827 + I0f6cb7a5a31d6f2f6178632c0c898bc6;
            Ib3b4cd6d8ab17869a2278552c02635c8    = I98b0bc583105e551a5c1c7a8b6de61e1;

            Ic298f77f42fc1d41cce684790036ecfe= I61ca60fde05ed88cce714dcd8c13b827 + I4c6d3d6fc2d10066a744fdd9405a7902;
            Ie7a5cb2ecb3fce35825785b9bca6b3bd    = I3ca304e8b6c5440935c6944b64ddde65;

            I805269f95afbeb6b93182f68868d08eb= I61ca60fde05ed88cce714dcd8c13b827 + I716ee53e79883f69aa045380a357e913;
            Ib9a0f8efd3dad427f247ce90fdfb94a4    = I33c7b994472de0942347e9b06ed9f59c;

            I881328804c45b06767af51e11182b27b= I61ca60fde05ed88cce714dcd8c13b827 + Ibf74a4dfaab7f7f538d2b5fac7394b63;
            I69a221a1bd95a588aa74b9bed0357762    = Id5395616ea942f63477bffe5c17560e3;

            I958993626e6e44e12f7c1e8026914680= I4907dd45c158dc7e0041c64f1fb388f6 + Ifbe479e5cab3cba43444bec1e12e72a0;
            I64f125cf2ca6a6da8a9cdae9e246c24a    = If90e3127bcb3ed51a225ce72afb0a793;

            If31528d1fc3a083ebc364e75cdd9c71f= I4907dd45c158dc7e0041c64f1fb388f6 + I62fdc8936121a2707d94cf3bd6e660ac;
            Ifac9dd60dd6c543aa94b39c599f0819a    = Ia6ff80807e320ef75fbdad7c86add89d;

            I4703b8d5a9033027889bfa8685e09e4f= I4907dd45c158dc7e0041c64f1fb388f6 + I42c1d469ff97913cbf15e3ebee6fdfa8;
            Icf062382a1e462571569ccee75b0a3ee    = If8a6eb502f55f58090ffd901b27086c2;

            I22d8e84d2db4b07111b7fdc6eef34cc8= I4907dd45c158dc7e0041c64f1fb388f6 + I991a7a7d562eb0a8b4b8d8f008ef2225;
            Ieed8b94295bed265961c4f52c3379914    = If10a93a95dd1f3e7117e64ae2915bcd5;

            I8b7c6df3b5ea575caab7820c95974608= I2c8f6a9b9f655b317bb0af4d60fdbc4b + I8c2e0c83a8204d6b21e0e3e458d56f05;
            I165eabcdde76821fdc308ff7a8c6d2ea    = Id86eeb13a357d077460584e1941e74a7;

            Ia8aa76bccf7eb310a9356e8b7ea1609d= I2c8f6a9b9f655b317bb0af4d60fdbc4b + Id435b68afb53bef4afc7b70a9512e955;
            I8b3542a6d64d6a7ebba4124bc6702f3e    = I5d7e70c0e768f5868bf9fa07111036e7;

            If9de547bf469b8424f1625e990f72b04= I2c8f6a9b9f655b317bb0af4d60fdbc4b + I56d1025271f1f7704a40dd7f0df02b0b;
            I7b68afec199be705d766c169f1ece981    = I48f780aaedbd67e6342d9e0232635ac8;

            I27d51b2015ea9af9bc345adabdb07b6f= I2c8f6a9b9f655b317bb0af4d60fdbc4b + I64c3d7be41abaa17d6992f9af8e72789;
            I4b6c8226ef2bc20dbd31d242bdb98b8c    = Ia9a47dd6aa0313a806147f2c4a91df0b;

            I93dddce2a0dc01ecb3039fac5cf04011= Ic7dff631559304ec59f0696c66436d62 + Ia1499972c4995268acd828c1289f353d;
            Ic3b4a86f22caf5b6103d52b6c9d2a991    = Id0a9c8069c91546ee6dcdcca1dbddd61;

            I746da2c1d5a620eb7e749f72f0f04a06= Ic7dff631559304ec59f0696c66436d62 + I0071f2168787bd42ab7f2370aed9d0f5;
            Ia37592b207086f63e2d94e3d7d26c740    = I3e30cc2747c9a7dd9c4fcd144f640552;

            I1e15f8d6fdb4ac732768d0cf73af829e= Ic7dff631559304ec59f0696c66436d62 + I4600963866dcb9bbea2515c805f885cb;
            Id0d786026e3ab0ddbffbc20e4d409857    = Ia4433ae2b484d7bfff269cb336831628;

            Ib719e667d7ba857f4f7432a245f4a30f= Ic7dff631559304ec59f0696c66436d62 + Icb91e63ebabc7a75a54eb7c731df4fa0;
            I333837f976cfc7f90ab0a6dcd8c1ce79    = I7aef236fed5567b77c8a3f5c22e3bff3;

            I4c6eec4a0c46e4f5d7c9734df48a16bb= I6a239d3e55b4a9a3be9989a85bbec545 + I3d1dd8b9c7c6d3913f7ac369ad7e625c;
            Id115b4708a49dcfd167e79ef6993e371    = Iff3859ddd94ff25ba5a08a367baf602b;

            I95623ec1fd5516040a9492aae0fc2b70= I6a239d3e55b4a9a3be9989a85bbec545 + I6261e0d339762cb2364421e6b87086cb;
            I666da645400344644e848ee6f7592d3c    = I4c0c110a6f362969bce6db69cb1c0bfc;

            I69017b49c11de463fe6d881e5c96a1aa= I6a239d3e55b4a9a3be9989a85bbec545 + Ib235af5b28d56f24372d3f0af816f2c2;
            Ibafeadd691eee03f855ed657c01022c9    = I51225282195bed9916ae55ae7887c1d2;

            I4fb9ed32471aa614ce6923f6a2279b36= I6a239d3e55b4a9a3be9989a85bbec545 + I673d1d0d0daab99bd940c46cc14ef55a;
            I10ec5c43a3fb65273053063001307280    = I58380b8eb6332c81366215b1dd60cea5;

            I2f0bc217c8a39d71adc1fc45c10b81c3= I630f905e55f08e7d1569a08e937ad216 + I79fe46308b93fbb24245fe1c75edf4a5;
            I05c778eb3588bdaccf714ba456f534c2    = I55df86c0751564116c4f1a65de2ac9fa;

            I0f1c6bb577ea2b8b2ab636e64378544b= I630f905e55f08e7d1569a08e937ad216 + I31e5b2cdc3dc571eafa37510076bcc64;
            Icd11e8d97a6ac6c0a73e8adee1f98c4e    = I0bc0390d7c9b369ebc92e9547b87b9df;

            I7a248af9d606c566e03977e985c280e0= I630f905e55f08e7d1569a08e937ad216 + Ia9e102d8679943c079f16c0228f0f0d1;
            If07c2223d4262e22cca9b77c3ed5ee01    = Icfe3de1a8dc46c883a65345392921c50;

            I0bf9d47bff47277de1e72518e8d88362= I630f905e55f08e7d1569a08e937ad216 + I62cadbd70b07a6a7a2974c7c392696b3;
            If0c8ce0ff66fe2806448f1c819d58ec8    = I4c0e5a2ba1c2b42970f41699d5ddcb9a;

            I24b6f4f68f291dc50caf03dc902282cf= I8d13eb3669785c4279c685763d4f3fad + Ia8d3667adc34b2b50acf7edb970538d8;
            Iccdc2371dfd9fda3e506adc2b1681ba3    = Ib81161d68b741b2656196d7284209d58;

            I79335b28eea15735f760b7a8b803e93a= I8d13eb3669785c4279c685763d4f3fad + If9f2a53dbf6e9b9a335a7657b7a2b468;
            I26e61dca9d045c4661b97afe346152c8    = Ib98bf53c446dcc7920b842d29191fe0a;

            I0b14b34b06cfa90539c2abca5639abec= I8d13eb3669785c4279c685763d4f3fad + I68c85727adecde0aa8aa66ed08c4b502;
            Id488d650b86f5def0668f4a1ef841b6a    = I31c34cf26a3890305171a6beca791fa3;

            I26878777354945712f834740b17dabcb= I8d13eb3669785c4279c685763d4f3fad + Icd8257d7f53d93db989eb56eaeb7e593;
            I479365266255d2228ecd86c350e8d38b    = Idc436d6b98d48c479d762c31bb55e071;

            I6cc5daed4de5950c02c0a57b993e22fc= I25a6f3de9a9a01cbbdd32ed848561aa4 + I03bea609a189246a2375b355df47cf81;
            I08d9c488fd85db45344e649699196263    = I49300b5a8d4f2ce3ef7238f75a2800a9;

            I52c382d5b0c4829127c011fae402ce04= I25a6f3de9a9a01cbbdd32ed848561aa4 + Iaec2f15665e83416bc140890f3cdde9a;
            Icde86d0ead44385b07e9a29057417417    = I4c1b051c518c4fa2e042e11cae60de02;

            I46ea9871e867034daa2d0501038f15e0= I25a6f3de9a9a01cbbdd32ed848561aa4 + Ia7046faae1ab05978e4b32bd44049fb9;
            I21feecd24d912ef3d0aec0e375958f3f    = I3ccb0a4c235cd79c6c11271aa1aeb8af;

            Ibb8a202599550e87831647a93a14181a= I25a6f3de9a9a01cbbdd32ed848561aa4 + I05931ceae6eff26e5a66a44a54d628ae;
            I59f419b3bc183a5fe743be3878fac587    = I8a2e9aba30b284e87bdbb6e91a30d9a6;

            Ibb79f2ce0b6028ebb638fc6661444cf1= Iba3dd4b2c2c85c4cfe770d9b52ef4634 + Ia784f35a5a46837b69eb048dabf84052;
            Ib0804d8bdda49ecd0024300eed52be53    = I29d269323cfbc900f3868dde96e8da48;

            I0d0c07d65eda2eee01df9c330c0d6f4a= Iba3dd4b2c2c85c4cfe770d9b52ef4634 + Iab354cc9ac1173335c0efeef694f3567;
            I37b0efdee34647a5111d698a5a80f367    = I39a53ef95ccd9c8b1b85e3214af441f3;

            Ie6940736944bac9be609b8d58b2cb13c= Iba3dd4b2c2c85c4cfe770d9b52ef4634 + If3a79ede332c39a8d2a276de833242f6;
            Id382a04e94d0749d0858041bdc5861be    = Id64ff7aeff6f73342f863be760a32a16;

            I472a71363435cb3ec054e00f9123ae64= Iba3dd4b2c2c85c4cfe770d9b52ef4634 + I306fec0aa68a0396053a6e0fa1cda38f;
            I368be992a21201268c41506396dcdcf6    = I083900fbd062835b505165f1da19e228;

            I553223e9166dcbddd1a51d0f92d68f28= Ie1b744387b5200a504e4874e14d2f282 + Ic8d47ff5d6c31601a57df868da78c2d4;
            I603a008893b5196d9f273b47a9d63144    = I7cf9dee91f849e28b2b2b38d2df00dfd;

            I495309d795905a53b0a3d3daa4f1f9d0= Ie1b744387b5200a504e4874e14d2f282 + I25c324feaca84e80f58075597e8c448f;
            Ie70d3a768bc09ddff6ac68aaba7d9f2c    = If54b33370dcdf69c464c92dab1248828;

            I21d358fd7673c4392f4e4b3d3a858b2c= Ie1b744387b5200a504e4874e14d2f282 + If64aa8c220b9ab6652e081da7e404e80;
            Ifb8bd837ada3d8ed5116db29da82d2a9    = I79c5230097571dcdf6ec2a15d633cdba;

            Ia1a60175112362f015c5531f7c48b90b= Ie1b744387b5200a504e4874e14d2f282 + Idee8c8144207d676d1f2f9064bbdff45;
            I978b93d46e20cb3eda70e5a976d62348    = I71efb4b4bb9b37a4e9b717282c5fbb03;

            I5644ece811bddcec04c9e3559c86109d= Icf76cb69aedf4db01cd3444f4c4ba471 + Ib504b808f724ca6032e7c746517cd4fd;
            Ib404040d4fb58f47f245184c3be01789    = I0cc336baadd473b40a866cb2944eb719;

            I37d2f9d3f05cb90e2d45bd578299885c= Icf76cb69aedf4db01cd3444f4c4ba471 + Ic308a5413f38b96d244cac3b0bc9462c;
            I9c664265c53ebffaad097b70ff3cbbce    = I42d8c11aefc92acf389d12e26217e867;

            Ie7d10f3c0f8b0add66d2cdd4435ccc88= Icf76cb69aedf4db01cd3444f4c4ba471 + Ia4131464996aabab8aae1db85f6a50e4;
            I781306c6b1ce0741d9c2fa06865f7a19    = I40412ee4da7bae7c7745064488928be1;

            I3c37396a1cef2f9e42b8ccc126db6eda= Icf76cb69aedf4db01cd3444f4c4ba471 + I5855124d566af739caa6511f8598f2c5;
            I16fa2e3dc0b3eddbc72811b51d6ac8ed    = I7f6fc13ef5b20f9f1646a608b63f6f77;

            I2f82390734079b8d289d48a6682cc624= I4857b5b50556c8e7fff4b2d3e08e4b28 + I8edbe77bacf1975e014faeee6b861980;
            Ia6f232495726806d01b702b0e248b2f2    = Iddd6e6676bf1c96936bb1dbecf6fd805;

            I9061728c3163ae684e8c5aec3e807868= I4857b5b50556c8e7fff4b2d3e08e4b28 + I1338d211b5d2d409bfe0df76d2ca2701;
            I66b3734060600caa45d699508c5083d2    = Id0a701ba3adbf20de140020b675cc363;

            I672d7ecc28a788c2602aff76187aa568= I4857b5b50556c8e7fff4b2d3e08e4b28 + I75838ca09e301b8e1301cbf603a1f8c2;
            I85fae6b23d086235a94a0162e2fb5310    = I7e8db4d3310c345d7ada4c2fe05cf9b6;

            I660b2fe99cd0bcaac34e9540118b54bc= I4857b5b50556c8e7fff4b2d3e08e4b28 + I50729db4a8e04f18979707df14cb2419;
            I8d6443d1be42203cb834345ae7e5aff5    = I3fba42f5d091f0b7a5d8b4d099f72284;

            I6aa263fc2a061d2c4059b08309f860f4= I0a1e9cf99f1d4725327615f50fcc3ad0 + I675ab6c4fb93b006f3fcafc985fbc405;
            I717332b7f76e9caf9351f1aa69b72a12    = Ia12c6ec292c6e9fdf58fe58a2af18a53;

            If3aef2d755013d195fd44f734365d7dc= I0a1e9cf99f1d4725327615f50fcc3ad0 + Ia9c043c5e8873fd13e39cf6bd8136c51;
            Ieebd34db071409288f489129b70ab599    = I37448ddc452e005ec974628ade793433;

            I3ad2e0bbff17683824f575deff82c6bc= I0a1e9cf99f1d4725327615f50fcc3ad0 + I566221060f06e724676ec9bec861d7de;
            I917c874137d64a9a495335c8f8ef5374    = I4dee5017c9b71edda82d50b867879afd;

            I5087dc4b32d29bfd7bad49026fa58a5d= I0a1e9cf99f1d4725327615f50fcc3ad0 + Ia3cb3ea64576a3e7332e1fb55953aa3e;
            I15fb4fb838d4a614c468f7d49261bda3    = I2115d9af1cbecde8b5e89c70e582de00;

            I8a7d893f3ef6d6a93ba552320d901599= Ie844f4c446983ce381b0bc4c0e8ef7d7 + I082aa8c413d7ef8f054b1c2857cbe39f;
            I2eb093d2a38ba8cf4be47d1d7f54ecc4    = I0e2c6c08e1bcd629678ff57f6bf23be5;

            Ic057537712e09fa794918e5cde87e084= Ie844f4c446983ce381b0bc4c0e8ef7d7 + Ia0932b3fd6a5ae6da2bacd2b86ba3a43;
            I8f9affdc5cda0fecc35dd15fc5aeb244    = I00a3c15421af76c65865ff21d2598055;

            I0cbab5173052c450504e3a7d15ffda52= Ie844f4c446983ce381b0bc4c0e8ef7d7 + Id682e531735437bc24abbf3d3d51e18b;
            I615a443d49d1479338d033d2a2cab51f    = I9fa21fd04ffc0a7dc281717e599fd443;

            I81ee40feb7abd0fec3faee653f778f5f= Ie844f4c446983ce381b0bc4c0e8ef7d7 + I3cb1f233951d49f985b0deac6e052bfd;
            I0635a3270a9653ca0f23c116fd5b2f97    = I66231fd914db4a60705f1d6de751077d;

            Ia344347a85d4e6afafa2ee3487e65def= I6067f47cccceea96ac46ff0d457b25f2 + If56555b7cf539750706cf678030ccdb2;
            I93a7c75ebce8fbf4c613b4d11dc98b72    = I1142cf230d2632a5972a95316f2fa15f;

            I038fce1597157a3d95bd9579cc2dcbc6= I6067f47cccceea96ac46ff0d457b25f2 + I097722547450582dc5776bdaff914741;
            I39334aa9d55bcc001ece37ce2a6c329c    = Ibe1b4cc79b063aafddadcfdb5bc4a694;

            I546585b819c289d855cd098818792e90= I6067f47cccceea96ac46ff0d457b25f2 + I0e2f746715b901feb69f6b3c94f3a828;
            I07e328d23da9383a296ecb03679ec74b    = I5371e6575d8bdc6f72cb08beca627fec;

            Ibc3a6609765818327e79519f3e348494= I6067f47cccceea96ac46ff0d457b25f2 + I7015def91103398e54f446ce3e43af01;
            I8a6e1eace6152af5c98c415804cb60fa    = I5e78e43fbf13f79a885bb3cee615d926;

            Id1c71a2a34f9e6239559d28fe2780907= Ifd6fd1f3cbf8884ca7f64bc42278e4fa + I8d0f440df332ea96e2d56eec490fbd51;
            I6ed4d6c350e8691b3a12ab51419cfa65    = I735298e3ea4442615df21b3699c94a7d;

            I1cd6cf5f8119d5e6b4ca40694399b1c2= Ifd6fd1f3cbf8884ca7f64bc42278e4fa + I3bfcd63e92f1949234ab1d2701dbb499;
            Ie2b9ed680dac51ac866cb830ca17ef84    = I1f2f072bb15b57b5437572b156499e12;

            I15e2a1b4356785d73e2ab5d51f1f5ec0= Ifd6fd1f3cbf8884ca7f64bc42278e4fa + Ia8849f78971a45ed0daa2489e7d27dd7;
            Ie439b520bbb0c8b29a5ecea167acb1c9    = I0344e18f3a5fe97467ba8e6641562f92;

            I803aeb29e66384bfc62744a841bcc83e= Ifd6fd1f3cbf8884ca7f64bc42278e4fa + I04874bd1bf257f205b5189c8c20e5a12;
            I9f8ef3295578acf5b0a42d074a15a70b    = I8aedaf42a56212b44d820d704945cb99;

            Ib6e220dd4f54410239dd0c791d84a700= Iaec9fd9e79371676bfa8ff14b4feae52 + I7cdc5ada6fc68ee31fd4062e2ff004d3;
            Ief01b06341d489e36ee344fd52084ccf    = If267b8451ce8bfd1c33273a9c5d08233;

            I8a009007fec23f4d492b0da1b6b404fa= Iaec9fd9e79371676bfa8ff14b4feae52 + Ie0622ff815747e4a9f368c74787026ec;
            I3b72a085b104e17dca3d8b2824f84e97    = Ie90356409910181f0ffbfdbfea6a47b2;

            I5f89adcb1ba235a74639eca119fb2655= Iaec9fd9e79371676bfa8ff14b4feae52 + I0cf5cb4cd472502b84dbf6fe1af0be78;
            I5e1f41e23887493db1d723e1e2cbd996    = I43a2d55679515c4766a6e7c19c3ba1e0;

            I8fd2b001ff154e4760ead2df355c80da= Iaec9fd9e79371676bfa8ff14b4feae52 + I937e3a8ede2305ea7c1750283224a870;
            I0e6f4c7bdc39bd22833f3d9fcfa55f1d    = I2b1e17eeb208749a9c320187e98f3c50;

            I581569cc2e63bc68a8466b07ca471b25= I500757c4eda5d3d899aee47b87da585b + I3f0bba472e912f11dea8e788fbc1cb63;
            Ie346802a8898b4b075be289e062b462c    = Ib9c8fc92cd361858e4fb1ddc6dcab191;

            Ia9cfdea21a65b0270de42cef7ebbf822= I500757c4eda5d3d899aee47b87da585b + Ie559401a3a913400dc5e3e5641297fa6;
            I82ea6f21706a97166ef11af548e80392    = I7ef5a40bcc9976da690ae85ee866b2d0;

            Id66a233d2e312aff939549dfa96a8cf0= I500757c4eda5d3d899aee47b87da585b + I4936f823841b0ffe32f801f5134c0211;
            I5f38764f6ecc2dcd1fdd5316102f1f82    = Ia52b8e11416781165d713f38018047d6;

            Ie479c12c25a1964c3804936d45725bdc= I500757c4eda5d3d899aee47b87da585b + Ia7206430a739a11af4d860096eedd6c3;
            Id4034bf7a0e92a6c92d0187e00d3df99    = Ibb05d1616c4b57cdf6a268fe16bb9ef9;

            Ie30d8770ab7e6643fcb67463f6999125= I47bf091b0fa74ad511a760bad9d2506c + I72c2256ba47cf03f95143df8f741fd83;
            I44692fd63388c57268ea9035a7e4c3ef    = I3be04ed5b262f461ad65b860adc6c601;

            I4a17ff532c9341e80f7ed0626f728054= I47bf091b0fa74ad511a760bad9d2506c + I1092325b801600fa7ec85fa640167da9;
            I0c2892a34e5236f1366959eadfd83825    = I0bcc8dd8d2adfb33dace6c005377ef97;

            I597bc1ec224007a78c25f7eea24c2c3e= I47bf091b0fa74ad511a760bad9d2506c + Ibf4c2c00f8e012e9498361bfd3c5b06e;
            Iccef2754044e7066e191bc5e1a3805f1    = Iad8fd338d5a105b6fe3a3a021f96f317;

            If198ec15fcf66e97e69f88f718979c2b= Ia4c3d0cd9957f678880de5775de76e0d + If26d90629e70c5a871e6f5b14471b8cf;
            I8ace46f1c56cfb3f4773324e0f8cae58    = I46f7c02eeea9f5a0058da869a84e57d4;

            I6aa13ef29cf7e86ec83affca4fa11e42= Ia4c3d0cd9957f678880de5775de76e0d + Iebd050e29044153d5881ef80b2db8c28;
            I94ec0139bd827ef5dce2c5ee9eb9aded    = Ie8e3dd32f3ccf581400d8dd0fd5daea7;

            Ide136b08f4b6211bca8cccf494a0baa5= Ia4c3d0cd9957f678880de5775de76e0d + I899e5f03cd1d52d11f898959559aaeea;
            Ied62b116607c549ff5918d5b95e2118f    = Ic23bbefb8e8e80ac5df4ef8a50aa5c83;

            Ieeab247764c23256749776b0a164314d= If5f957fa2f055b1c2c28e8d7cfe3e9ad + I4c03a6569d1b954d088053e38827e811;
            I9efa5796297bc922bc5fe17f8319a515    = I7c56e54d472bc2301521ecb93aed0ea2;

            I210e9ff7f4588185bd712915954543ce= If5f957fa2f055b1c2c28e8d7cfe3e9ad + I0c5250aaca86185fed5978438c8861b6;
            Ifa6908d8fda29713d7c1bbaa69b72b53    = I4979d09a4bf88992a280e598841f5e50;

            I59186d5219833d6dd2e813a2910a61f5= If5f957fa2f055b1c2c28e8d7cfe3e9ad + I59c80c7ec26f43308b1a646c47160568;
            Ieb46857229186ce0391cddb2d30f434e    = I15264bbbe49fff9c53b8066414264010;

            I0c8b2bb61a9c3a67ac7e03e40be2b98e= I3608378a5da8c66bef58528d56192530 + Ibf1c9d86665f696d91c554db748ff42b;
            I67fa03f808026b38ca5b4e71e21588bf    = I32293d41086053c7055fa40ce224631e;

            Ide24c1f9033e7057262da1bc4762b840= I3608378a5da8c66bef58528d56192530 + I49ccb3e14fe61618806e791ecb4f4eae;
            I70938dfe09b0da9d87dafed6af3fa05c    = I4bd0008f9e9598e9f60a0aa8c2aa2da5;

            I4677558b9faf190e7960cfa9b8ee00fd= I3608378a5da8c66bef58528d56192530 + I8a954a331d36266465a0813d2e8b319b;
            Iff30a4e14b6282e9ef92e7f58230b516    = I584861d31ee7ff0efc61b192c64bca32;

            Ie38ab94215851e531d2100b6602d5fa5= Ie6dead855e00ea0a8e6a9b7503aaebb8 + I239a992ebb62899120a74b1c9e6cc4b4;
            I43e0faf8070869ab0528a7a4a5cdc103    = I64f092a873fee78a333072d8c5bbddf8;

            I3f5119e8fac99376aa38e4765b8b0f99= Ie6dead855e00ea0a8e6a9b7503aaebb8 + I2e802c75c6ce34b05943b678ecbfacb1;
            Ib2f0333fac7701ae4a5589d54005b8f3    = Idd6f95a4386cbea3c1533683854a4c75;

            Ie8040301d224f78c1fd18bfe9e29e5ba= Ie6dead855e00ea0a8e6a9b7503aaebb8 + I05ecce409cca00ea5b0df25de5a50cf2;
            Ie4e1491da700923e81b2c1a246e528b1    = I32710d1855b18d6c70f6e23a0a440a69;

            Ied989966cebf0d730633606c5182a249= Ie6dead855e00ea0a8e6a9b7503aaebb8 + Ib49e53ca8efd9564ee9572eb3089bb51;
            Ie8602467de2ece2013878a6b8d3129a1    = I32cc6023f28c6dee2b4b097f1fe890d6;

            Ib8818bc4ca106ae38cacd5c20083aa08= I3bae5e6862e003a8b9a476f72cc6858b + I420e2c5a8745133f6263a71b458f1e2f;
            I85c93c62f79b1703cb6928f96737cf27    = Id91b5daa1685f0e3d492f0c3c8306f8e;

            Ibf08556fc39044222321912e84a4436b= I3bae5e6862e003a8b9a476f72cc6858b + I9fce6091885f1bb97d29fb1f543b1a38;
            I3dc816ee6c2a818b32f6d4e1228704bf    = Icfdd224aa430648d4afe7b224340b91d;

            I985e2740ac0f656da8f9dd973bca99e6= I3bae5e6862e003a8b9a476f72cc6858b + I2de1ca2c390bdd3011fff4a359bb5332;
            Id34d83701e815c01359bc5cd1b9c993c    = Icbcaa7780b1ad02e07cbbc871b0c2729;

            I73012d2d9f6f237bc50bbffc199e012b= I3bae5e6862e003a8b9a476f72cc6858b + Icbde2c6230e9cc67ef12031e38bb344f;
            I0a20e3e26261ba558d681346649cf0b3    = I587b0b57b4f95e8533842965674d1416;

            Iefd0d59e58623b14437b17297fdbf4ff= I4431adecba8be9e5f21bc6b3e1f8cb10 + Ia47f7fb27f2d965cfd2989569c257356;
            I331c6e8dbe2ea1e2232f82766926d0e6    = I1188961bb659f61f0749a27f4ee5c62d;

            I68d2443e98f2fd3fa3baf96f98e1f4bc= I4431adecba8be9e5f21bc6b3e1f8cb10 + I034fb3850485fae2d1358041a1c41888;
            Ie27046fd2751357e4a81dc62086f00be    = I4ed124c919ba9e29d61a5f771b554ead;

            Ia2d1b6833cd8ed02f05281e508e4d716= I4431adecba8be9e5f21bc6b3e1f8cb10 + Id968b34075e351ab01d65abcb4ed8cca;
            I0897ceba8201bc14a49ab30318183875    = I735b52f16a8beb195d3e7332f39a1c86;

            I512e2251bef73108eb0f3e01e79ca3fb= I4431adecba8be9e5f21bc6b3e1f8cb10 + I2e22e867f6f84a7807b82f64a147022e;
            Ie7b15aa8ce2492bfb433894efeb967f3    = I626977a5bbbdb2da503472e8fe6c9569;

            I9bf64811d14ca8b4c633342ad22669a3= I21c7a2885126d532d00484376588a469 + I174fcbc2ee01fc55edbc8238e5da7f0c;
            I255add08e982f701508a98db221e617d    = I8f2450ac5c97afe557d068ee5760b527;

            I45a910acd40d5b9417bdfdc50cddf241= I21c7a2885126d532d00484376588a469 + Ia40dad546d9c852e2fa8942c62a1c1f8;
            If7ca4919fa1449f38777f742ee1fb875    = I13834193a9eb2706cdc680b303efbcf4;

            Ibbcf5c5f4528b03508b506c43e4511c4= I21c7a2885126d532d00484376588a469 + Icd9a876a0feb16ea62bcad5be2004dac;
            I24cafcb5b9825321c54e84827a662fdc    = I798a185688b52e59c92b42161b3da7e7;

            I2b8b54048e164ef2f1c072517fdfe400= I21c7a2885126d532d00484376588a469 + Id9704e1d8096cd28577c5c357d30b7a4;
            I3ede71cb7cb39774aedb9889240a2462    = Ib695cf55b921ed43db22362a28761714;

            Ia48d8883fe4f685477da6b4b05ecd387= I2c4d7339ff2fe68d060dd8d961dcab8c + I6dc671e73b4e9c70cabfdeaac2e5c40b;
            I24da9598a6840d3ba7b12fe4f638219b    = I1dd0afb6f1a979176d01ab7d37f39bed;

            I276395da1f3f1ae246b082408be2cb80= I2c4d7339ff2fe68d060dd8d961dcab8c + Iacf6340a29a5592b61ea875304a2de48;
            I0358ca8833007cec4ce5047db32ab7a3    = I559878eee7f3bee345a0f0e891dd2c05;

            I4d0e2e01d9abf9ce839fe650abfaaddd= I2c4d7339ff2fe68d060dd8d961dcab8c + I487391402b6aa27bf212724a37ea9c33;
            I85b5354463c1c15f91ed67292da912c1    = I6c688b7c6f01ae353117029f80487ec4;

            I7e4e7909094f762c54137cbee99255e5= I2c4d7339ff2fe68d060dd8d961dcab8c + I4b8554cab486a4fc1e14884a6495016e;
            Ie93731739ace44811198d0fd95b04a6a    = I62ad8f36d1e0b80d0d04a326d80e1729;

            I761255e100d161b25645ca3a5187e82a= Iee518b15b067eec58cccfa37f7432ea5 + I94e89b3a841f9760e3967c97e86d7160;
            I464926faf4e005ad491b0bf93a365e07    = Icf1eb32cfc4a48f7e53c180aa94f5833;

            Icc2ce1fa3cde69256378ec3f4a07b0fc= Iee518b15b067eec58cccfa37f7432ea5 + I5975ef8f6cf53cf2132cdd9d707e7912;
            Icdaaccfead6f2d5ac2ce19caf1104d57    = I8bdfadcfa5cb308e6e254d42997340fd;

            Idd99afa80ca23644675d3edd60e74fe4= Iee518b15b067eec58cccfa37f7432ea5 + I6c19936ca2edeb0e261e880a1055e964;
            I916d6f9429f2b0cc1bd6fb900484cde5    = I6ceae370fa59e601566286b127dec684;

            I486bcb4fb0af80c98c2ea21ac64f7a90= Iee518b15b067eec58cccfa37f7432ea5 + Iaa235d085a5916a3b0814c3ed2a9026f;
            I0142f9b3d361a0d88522f1c5f54aca84    = Ifcf5bef8ae2998f0bd3d270e98acc1c5;

            I759cca2c0003fc2c2af7709c5ebc59f7= I42145be9c2a80288ba4a2edd91f661a3 + I8d431a0524241fa54cf6dd1e79de4c74;
            Ie6871983b4f81b5321519647e628bd0e    = Ic1c8e5992501f0e04191fe6dadd2d56c;

            I1d5ce9f132cd1f46e96b511c77234e21= I42145be9c2a80288ba4a2edd91f661a3 + I7b8da162c08f8aa2ae90522ee1526cf6;
            I17d7be125df22153fc1ed051d4e0770a    = I3f88a35a94c77ca32f3b58c4b509b21c;

            I032e26ea05e88c6d325a810b67e82306= I42145be9c2a80288ba4a2edd91f661a3 + I7fc190647082a3d71614f46f670167bc;
            I50b13959e06243e54fad2088eaf65aa7    = Ib875be40a1b73b1583cfc9cfec760e31;

            I0f72df5225a1fec2f276fd3c9138e8c3= I42145be9c2a80288ba4a2edd91f661a3 + I5d86ce0b58c0b281d747116a9069ef33;
            I7a423d609b492f73d5a322849b4b1cce    = I15eae5f35300569305dc03e24d1cdd7f;

            I0d18cf087b2335f1b9e1a621acd5379f= I9dc297ad41fafcda77f5347f331cfc25 + I59547aacdcfde31dc016ec2acbb2f4b4;
            Iefec67e214d1868670a34a7297d4a1c8    = Idffbcb47f4a04fc71d1406e46f4ab6c4;

            I7684fc23c57105e856050a45640f2bfd= I9dc297ad41fafcda77f5347f331cfc25 + Ie4749f8e9ad2b370f9f9814b5a463c43;
            Iae7da7fdc002b635ce4285d6916d8156    = Ifaf09d72a75fd4f9948e997b8a8388f4;

            If778767ab80e59e940deeaa8a0dac99a= I9dc297ad41fafcda77f5347f331cfc25 + I495f8be463b15db906474c518e0741e2;
            Ic561e44b2caeae84df6720f1afa3e8f6    = I661c1624e4d13ba49efc3fb608ba84ed;

            Idaf86833beb8c334f99291db9302ed29= I9dc297ad41fafcda77f5347f331cfc25 + Id20394136fb036435bb4680aac64581f;
            I5be062f5b52e104ca67e615ce75a7c80    = Iaa8bf572a01757f5e9321e6ff7364d7e;

            I6610e8d41cea10498d95850440ce388b= I846700c79f30ca954cc2933fc94d355b + I5ffed139764d90825b9f2eddacd0eddc;
            Iecdde23e34c34ee0055be41f44959a19    = I7ef389b5ce4bdcca7fab9e9ec2bfa3a9;

            Ibc653e701eb995e828c8180efaa122c9= I846700c79f30ca954cc2933fc94d355b + I733c3fa4d84e5680792b16a70bb1a51d;
            Ibe09be9cad0e56d5403868d072d7d628    = I4e7823ff42f8f44a21778dc4b3633a67;

            I21d36c49c9c766139b4b01df7c00a8f3= I846700c79f30ca954cc2933fc94d355b + I3c057d64cf4fca0238a874f0ced99c76;
            I464e1f3c13acaf466afb354a9b35ba0a    = Icf5823b64f3a9b7d2656656b61724bcd;

            I0e4ffded936d7ccfc32b410aec617df8= I846700c79f30ca954cc2933fc94d355b + I8a16afac6e470ca69634d7fe9656387a;
            I160a465c22073a53510e8a4c489c3321    = If77f93c61b38d10360f7dd382686d91c;

            I1a5745021323efb5327d0b893962e852= I8af96a91457316e49e3f7dd5e57c82da + Ie0667fbe76244eaec0b155d69dcc9447;
            I9e86d3e49827861b24f4fbeb308ad3a4    = Iede699ff40abf5838b54678df24ff29d;

            I65547afdcd7fedb7b44bd51358eec4d2= I8af96a91457316e49e3f7dd5e57c82da + Iedb9bb14951bf67bc8865b0983490c14;
            Ib96b7d796e20967e89a47e01bf424e59    = Ia1c9e86b6112a18e7aa613315343e696;

            Iada3eb71e94ff6a6f4e5c702e83036ed= I8af96a91457316e49e3f7dd5e57c82da + Ic78949e07e643f571f23df7e8f15d9fb;
            I565e666f6ba14b4c25e0dd402a3266e1    = Iad94272a2a302f4b6b963e71ccd64ccb;

            I077404a911da16d707a326f18717dc7a= I8af96a91457316e49e3f7dd5e57c82da + Ic4e7f690bc050f1d1f84eae7ca193e1c;
            I97e8bac5becd5128bc70f3bb48f73e6c    = If4d54d2b483d85b0c4f31db721b14323;

            I6da1e92759c96aab8b9207a9acb244ab= I7d1c247500d7d32e406b2a5f7e2b745b + Id4a213e494f9c9be0fd1a307e87c756a;
            Iced39475c6e5e3d8f36d2a5c5a80f146    = Ia3b12887d984da936d88d657090f8972;

            If7110182720ffa279b1cec1305cf9889= I7d1c247500d7d32e406b2a5f7e2b745b + Idda26504e422367082caeafbb29871f9;
            Idcbd423c2b963c1f693dea2ddf428195    = Ib23dbfa64e4a9364e0c1dbbc6b2ff001;

            If0e20ea1696ff84329b9928d7f9e3381= I7d1c247500d7d32e406b2a5f7e2b745b + I461ebbf3a02ae63e2eb27531b1370f24;
            If1640e294bdcc51ee12fca5b3a33be6d    = Ic8d47dcabda3b23d4451e609395c4698;

            I4e69ae6e73a856d4e26203fb9acf3565= I7d1c247500d7d32e406b2a5f7e2b745b + Ia60421aa427236540b4d0d08d52ff507;
            I4754c6c355e632d2ed1336b5a88c3b46    = I5d4903ecdf83967c7f60d876bcd0b215;

            I64c939aa568669b4567c21be09ad0e94= I66d85c030a8864505298919046056305 + I5e2331edf6e881e9f3a8c47eebda0ac4;
            I1634d703ad5d6e58a97b13ef957bdbec    = Ief11c4434035425db82902c38e47be48;

            Ia88eb16f68265e322509d541eb457993= I66d85c030a8864505298919046056305 + Ieb0336a1974a2aec0966f4f59f460802;
            I804e1e6a01edeb780b0159ecae707b71    = I1c3a6173bb59263a31998a5a69aaa38c;

            I916f75e5a3858a420ab5cd4c43b13921= I66d85c030a8864505298919046056305 + Ib028686da9c849e827cf249a744b7db3;
            Iea3c0f3c3c3017fe87a3b01647189fe0    = I2d77f481539c1258b61c2a6ca7208455;

            Id076f99460a8f73a9fd43467216e8f8e= I66d85c030a8864505298919046056305 + Icace650ee3865bd7bbddd2d9435c5561;
            I756b7d7e6bd3e71afa472e7e4727264a    = Ie88dbc3340cd953d819e7fa12d1fe3fb;

            Ib4d7aeb8544fbdc36575a55b9f67f2dc= I4841257ae596d9d3e4eb1e6f886956b0 + If2b17f9e9186542117f43d0dd342326e;
            Ifbeae0a2acf80eda6ffd050d3bb07eb3    = Icad54aaa6f380f2808749db56b76a959;

            If65d2514892fb7ee64fa4dc37fc0fed3= I4841257ae596d9d3e4eb1e6f886956b0 + I0b0dd019d8bd24684403a29aed668b6d;
            I990ab4dcb70ee860c2c40f306ef314d3    = If41dd08de4b2e28dae0404832fa0edd4;

            Ibef07e48768252e9b41baf067bb1ff5d= I4841257ae596d9d3e4eb1e6f886956b0 + I831d214dcb4f8d534b5ddaaeaeeb81ce;
            Ib131087ea9ccc4bd161c3f9ac2c72303    = I161c799aa59a0d82ca4db2b7b0293fdc;

            Ib8fb61fa9cb8e92bc57c53a567891895= I4841257ae596d9d3e4eb1e6f886956b0 + I7d27d070b96b7810f667e1d1845342d3;
            I9a967ac9d11583faaa783984229aeb2c    = I911555064a463cd6a7ebdb4de801b8fb;

            Id8f5f32cd0757b4d6861d17fcbd6e8d0= Icd6f7ec117f9ab4eda8c5eba41386ffa + Id4dc304aef5f35f6ceb91796c278e716;
            Ib9921dfcf121e5f4ac4d8be83a868210    = Ib2fce59707fcc6d804b748678d3fa03a;

            I8be241f29e7eb258e9b3501430820b0d= Icd6f7ec117f9ab4eda8c5eba41386ffa + Ieb3f28762410fb40a0c8a8556b4b3ca0;
            If22d8fd45caed08b2c7cee8b7349700f    = I5d40a4f6c096b4962285bee680a366c0;

            Ica8a188ea43e2f28e70b8ea4e2431dc3= Icd6f7ec117f9ab4eda8c5eba41386ffa + I6fb55222b69475b7168874423226ec9c;
            Iabf029e67c7f827faf17b6518cd1bfa3    = I692db6abe25b064802b76618cfd8d151;

            I83ceb726e57d52698b57dc39ce585897= Icd6f7ec117f9ab4eda8c5eba41386ffa + Ida7ec09c913caa0e78a2c4cbaae517c8;
            Iaeab83001c6285630e3404ae67227f46    = I396539ceb8b33c1dfe096f71954586e7;

            Ic88e7e05d83ff800b4a941ae4b424557= Ibc0498839d1d9b6dc853b8e5d7a88fa3 + I927c870d09285dcb47e6d399f319471e;
            I53ac6d02d2bfc9aca9469148753070a7    = I4335c153299e851249a1492c14987447;

            I7de81aaac1e5776dfb60eed2d12d4f6d= Ibc0498839d1d9b6dc853b8e5d7a88fa3 + Ib402cdbfaa9900820b85bd625415c547;
            I61992979f60b26d313efd1dc23bb54ab    = I5d81087b001624992357f909d2d7e9e2;

            I37058036bd9f4331387ee4a9348541e2= Ibc0498839d1d9b6dc853b8e5d7a88fa3 + I84da4ce7441e132e775167c1cd81dbe5;
            I8b46b3f0835310114208963de7ac8e97    = I2b8539d21de88ded1152a26741003b99;

            I570f85838c418d8501c8ccdc38a53f00= Ibc0498839d1d9b6dc853b8e5d7a88fa3 + Ic5eba898858be1f768841ead792d6d86;
            Icda26ba6f5c7f77a80776b2c1bbc975d    = Ib5f0b838019cb6c583e7aae384a7ffba;

            I4aa6f0c0f5163b944f11328888af73e0= I142ebca7f155e287e38ddf45423ab0fd + I4b8d520ee88fd39d83a16432e962f731;
            I0863565b3ae88137a2384750436f9e19    = Iee7fb9e4ff68c15395c13083bb14e8af;

            Ic7fc1f38ad4e9b2cb472ae75bc3c100c= I142ebca7f155e287e38ddf45423ab0fd + I0e7079db66c15210046b997f319ece89;
            Id646110f8d09cd47dc7695e05f73efc6    = I18176a5b74de8d98a21cbbbfd35b0bdd;

            Ibace8d2fba25834c83b1e57195c81086= I142ebca7f155e287e38ddf45423ab0fd + I8f8273c4cb2a9ace8a09847efd4bdec7;
            I5999eef2304e579a3d47e4f15ba336e1    = I033c58d2361a232bcfa2eda4ac665761;

            Iefc1488e3eb60b99ae08d904a15c5242= I142ebca7f155e287e38ddf45423ab0fd + I72197797a307c611fa8952533e63d7bf;
            Idd302bdc6ff8368a6b73d53bbc8f8425    = I0ddecbd9a2e867e3bf8a447434f626a1;
end

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
              Ifc045af19c3f10d92d2b0dfb4fbbde38 <= {(SUM_LEN){1'b0}};
       end else begin
           if (I65e382d77592c7d1af308d171b27ff3c) begin
              if (Ib325dab091dfc3a1a269adb3ea9c75cd <= HamDist_sum_mm) begin
                  Ifc045af19c3f10d92d2b0dfb4fbbde38 <= Ifc045af19c3f10d92d2b0dfb4fbbde38 + 1;
              end
           end
           else if (start_dec) begin
                  Ifc045af19c3f10d92d2b0dfb4fbbde38 <= {(SUM_LEN){1'b0}};
           end
       end
   end

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
                 Ieb085b219090cde5da2190093ce43730 <= 'h0;
       end else begin
          if (I65e382d77592c7d1af308d171b27ff3c) begin
             if (HamDist_loop == 0)
                 Ieb085b219090cde5da2190093ce43730 <= HamDist_sum_mm;
             else
                 Ieb085b219090cde5da2190093ce43730 <= Ib79e305e6f44a4a6ebef1db5c70246ea;
          end
       end
   end

   always_comb Ib79e305e6f44a4a6ebef1db5c70246ea = ((Ieb085b219090cde5da2190093ce43730 * HamDist_iir1 + HamDist_sum_mm *HamDist_iir2 + HamDist_iir3));



   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= {(SUM_LEN){1'b0}};
       end else begin
          if (I65e382d77592c7d1af308d171b27ff3c) begin
             if (HamDist_loop == 0)
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= {(SUM_LEN){1'b0}};
             else
                 Ib325dab091dfc3a1a269adb3ea9c75cd <= HamDist_sum_mm;
          end
       end
   end





   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin
          converged_loops_ended <= 1'b0;
          converged_pass_fail <= 1'b0;
       end else begin
          if (start_dec) begin
               converged_loops_ended <= 1'b0;
               converged_pass_fail <= 1'b0;
          end else begin
               if (I7d4dc5e91ba3d952184d90de12f67bd3) begin
                       if (
                         (HamDist_sum_mm*100 > Ieb085b219090cde5da2190093ce43730 * HamDist_loop_percentage) ||
                         (Ifc045af19c3f10d92d2b0dfb4fbbde38 > HamDist_loop_max)
                         ) begin
                         converged_loops_ended <= 1'b1;
                         converged_pass_fail <= 1'b0;
                       end else if (HamDist_sum_mm == 0) begin
                         converged_loops_ended <= 1'b1;
                         converged_pass_fail <= 1'b1;
                       end

               end  //I65e382d77592c7d1af308d171b27ff3c
               else begin // else I8bf8854bebe108183caeb845c7676ae4 I65e382d77592c7d1af308d171b27ff3c
                    //wait for I8fc42c6ddf9966db3b09e84365034357 start_dec to I01bc6f8efa4202821e95f4fdf6298b30 I0d149b90e7394297301c90191ae775f0 I3262d48df5d75e3452f0f16b313b7808
                    //converged_loops_ended <= 1'b0;
                    //converged_pass_fail <= 1'b0;
               end


          end  //start_dec
       end  //rstn
   end

//tmp_bit valid Ied2b5c0139cec8ad2873829dc1117d50 Ibd047e2643dc68affb5b4f25b82ded31
// I7fa3b767c460b54a2be4d49030b349c7 I9a4c07402cc2f3740fb5849a16920e13 I7243f8be75253afbadf7477867021f8b I13b5bfe96f3e2fe411c9f66f4a582adf I724a00e315992b82d662231ea0dcbe50 or I190ebdd6b6c2b422296a6ee2cce59699 I0aa6f4210bf373c95eda00232e93cd98
always_comb HamDist_cntr_inc_converged_valid = I6d3acefe6d7dfb94a5d66dcaa1bbbb76;

assign I204375b1fcd1f62621b32a06a9dd0bb6 = I748f85f6680918a2e992df339b4b6558[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[0] = I204375b1fcd1f62621b32a06a9dd0bb6;
assign Ic0ae28dd2fa2d9e0b2a9edaaffd88aff = Ib0f57837099e3fdf1b908d78bcda4a43[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[1] = Ic0ae28dd2fa2d9e0b2a9edaaffd88aff;
assign I63323f8807804f4534429d8aeafc7d23 = If75e99660e3997f53f7b903bc366f47f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[2] = I63323f8807804f4534429d8aeafc7d23;
assign Ie8554592e62dd20a36ef79e06af24a22 = I3253481bee7dbfc0f3eac94c3252ee4e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[3] = Ie8554592e62dd20a36ef79e06af24a22;
assign I67458f3b57d906d3626d4e7656049538 = Ia80693da8182ee2c3708b6ec21d397d2[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[4] = I67458f3b57d906d3626d4e7656049538;
assign I523d96cce3a523da8ca8e065aa5d8f64 = I7fa3f2648baacebf9e4b59c179601fa6[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[5] = I523d96cce3a523da8ca8e065aa5d8f64;
assign I3fad2338742a91d05694c9bbe0584126 = Id7699f8f89380c315303644fdebacb32[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[6] = I3fad2338742a91d05694c9bbe0584126;
assign Id30ee39232f016f983f45208ed802126 = Ibf3e1ead3776901898d4b154aeb61267[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[7] = Id30ee39232f016f983f45208ed802126;
assign I149dbd0f3f68786fc3a842bb0064f0d4 = Ie486617fc1d6354c7f347692cdbd894d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[8] = I149dbd0f3f68786fc3a842bb0064f0d4;
assign Ib383a8f851cd16df009c975ec7efb305 = I7ba403c6745e7d026282ad704e065702[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[9] = Ib383a8f851cd16df009c975ec7efb305;
assign Ia2227bb2140f18af451ea4c397262178 = I93cb3974b8594665b2e7ce5593fde69b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[10] = Ia2227bb2140f18af451ea4c397262178;
assign Idf0b6d7bfa5a9a38e1362c4b3b0d5b99 = Id6a9ab06d58c3a01e1fe04fcf61406fd[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[11] = Idf0b6d7bfa5a9a38e1362c4b3b0d5b99;
assign Iaa15139339207505f231f71669ce022a = I261bd53528b82128acabd405389c8d60[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[12] = Iaa15139339207505f231f71669ce022a;
assign Idc30dece6bd74ad2ff6c0822347a800d = If7fa833bf1b1438e7a5bc783ee745252[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[13] = Idc30dece6bd74ad2ff6c0822347a800d;
assign I7492572ef50294af38fc778e173a60fc = Ibb103853fc21f8f3d466ca16557ccd3e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[14] = I7492572ef50294af38fc778e173a60fc;
assign I4c6718b74573391494789da2e33c1e2d = I37446eb66ccfd268cb418655b8160fe1[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[15] = I4c6718b74573391494789da2e33c1e2d;
assign I03659b77af3e47129d9206af314ec521 = Id17f6250f8c7f1d7f75fd27f92698da3[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[16] = I03659b77af3e47129d9206af314ec521;
assign If0fbb2a55965bb66cfaad70fd9241456 = I9957b02e8d0d888e6950eb553d9084d7[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[17] = If0fbb2a55965bb66cfaad70fd9241456;
assign I4f8bea1f3f8cb9ff1b6d1388c6377861 = Ic71258b745437bc8463fb4f847c55e27[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[18] = I4f8bea1f3f8cb9ff1b6d1388c6377861;
assign I765559024522a12448e338401c10f800 = I24bb5c315eacf0f4e8c86f6582389e39[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[19] = I765559024522a12448e338401c10f800;
assign I815daf68a1ed9f91b02ede68298cc5f3 = I607f203694ff76930cfee4103cb73c30[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[20] = I815daf68a1ed9f91b02ede68298cc5f3;
assign If0e526189886cb9e8af7be4797d8a637 = Ica8e4c56ebb37e189ca8e6b3daafdb80[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[21] = If0e526189886cb9e8af7be4797d8a637;
assign Ic8dfeb5746649e88e59887cda08fb62a = I7089386c94261e0febf3b4f7dc1aec30[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[22] = Ic8dfeb5746649e88e59887cda08fb62a;
assign I0bd3e1beb510558b20c2b4f0f8f20e76 = Ia1e4f20f32f7371cb0078d6e80fe8b7e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[23] = I0bd3e1beb510558b20c2b4f0f8f20e76;
assign I647c8a9b1fd2281c8e129d2cebdd597e = I790cbca796af58b1726d0a4680cc164f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[24] = I647c8a9b1fd2281c8e129d2cebdd597e;
assign I6a803347e6d25dbd012caf725e35c256 = I0a93f095f9efb1542116a295c0db9c8b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[25] = I6a803347e6d25dbd012caf725e35c256;
assign Icf6deff8d81d69b92659b257bbdb53c7 = I989ba39f188a44475a83e65a4960d2af[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[26] = Icf6deff8d81d69b92659b257bbdb53c7;
assign If282e264f908747340e4e4d2022a66fc = I9bcc1d9b3dd258fa7b6042f0185d48cb[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[27] = If282e264f908747340e4e4d2022a66fc;
assign Ib5ca6dc87c214c3d73b265fa0e242452 = I9ba14715d9f33ef45681ad52f5be9593[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[28] = Ib5ca6dc87c214c3d73b265fa0e242452;
assign I3b8dd3a8e7b21202977c976ba687cb7c = I396a897f79b519f4fa02af39d0274f64[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[29] = I3b8dd3a8e7b21202977c976ba687cb7c;
assign I4e1743e1634bdb7ad6e8d072e19f0abd = I197c0cd576e16ee2197a28c86397f801[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[30] = I4e1743e1634bdb7ad6e8d072e19f0abd;
assign I4ccbbd7d8e03a7c7410acaf35ef87608 = I094a178e55425f27ac1ff6195217396b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[31] = I4ccbbd7d8e03a7c7410acaf35ef87608;
assign I1848d733a31c474bcb2d3e4b9b736e94 = I3177408f7d08b431be99297fb10586e6[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[32] = I1848d733a31c474bcb2d3e4b9b736e94;
assign I6fb841a6fe0ad7d433f1a182706d6ad6 = Id4948c876d48bdbf317d32f135e645b4[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[33] = I6fb841a6fe0ad7d433f1a182706d6ad6;
assign Iddb16107d5ce4ef65024a1cd5387dcd1 = Ice5ff01d4fb4583898498651a0ac0171[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[34] = Iddb16107d5ce4ef65024a1cd5387dcd1;
assign I8eb4596c73d1cb6ae5a783a6582cbffe = I0fb33a5ced3d15622c9aefa188052e24[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[35] = I8eb4596c73d1cb6ae5a783a6582cbffe;
assign I014c1931d012f79e954a12e10178f1d9 = I0074e1c3ca0ff903a9201ac5fe7ca841[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[36] = I014c1931d012f79e954a12e10178f1d9;
assign I8ad79c41a8896712d7c26d29c0b1e7cf = If65f587e987a51c093e8dd4df532e26c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[37] = I8ad79c41a8896712d7c26d29c0b1e7cf;
assign I1b16bbdd1e23bbe571bc7769731a03d8 = I33d7e77d08590f0dfb1867e741dd8b6b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[38] = I1b16bbdd1e23bbe571bc7769731a03d8;
assign Ib0cea939898e64f9ec4ee41aa3f062fb = I678c22563e0273403b046df4261f21cf[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[39] = Ib0cea939898e64f9ec4ee41aa3f062fb;
assign Ief16fc889b2326a53224b3b60ecc8955 = Icca700c12ae2e8155ca6b41e692e8a8c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[40] = Ief16fc889b2326a53224b3b60ecc8955;
assign I774b99eb9e3c3c98ce6dd3c60df7eff5 = I5ed74e81d2497681af5a0ca13fe23088[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[41] = I774b99eb9e3c3c98ce6dd3c60df7eff5;
assign Ide90044338620a38b90b5877ce0eb52b = Ic7fa6b8cdfcf7d83d4e101d9c8b7b34f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[42] = Ide90044338620a38b90b5877ce0eb52b;
assign I2271e9b3a663941eed3b939bf80ed2a1 = I26010e26e22d8a2ea831e86fae34a24e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[43] = I2271e9b3a663941eed3b939bf80ed2a1;
assign Ifc1b458539905b3557d79c94954747c0 = I578efe5c2c504f12c8f2466a7f734215[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[44] = Ifc1b458539905b3557d79c94954747c0;
assign Ibe27dea48dd30331b9723a1aec226f0f = Ida86d05f907d23ff9fed06927c2ec9d9[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[45] = Ibe27dea48dd30331b9723a1aec226f0f;
assign Ic214eae29f89949c797816779332aef2 = I9d9f8c7a23d9750ec44e706bf763df76[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[46] = Ic214eae29f89949c797816779332aef2;
assign Icd48fe364089e0250b4fee636590fe28 = I0b41b002a32b8e9e2fe68e819f228fb7[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[47] = Icd48fe364089e0250b4fee636590fe28;
assign I15d7c9e33bce9e3ee1059f73832bb9ad = I0e872d4c07169cac84549178fa144274[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[48] = I15d7c9e33bce9e3ee1059f73832bb9ad;
assign I9514bd70ebe24af7d8bf346ae09219f7 = I6f4ef0f404ae046519b8436171d51e09[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[49] = I9514bd70ebe24af7d8bf346ae09219f7;
assign If987109479436b8d51629513310a948d = I4d04e66ad9103a685fbe088b74517452[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[50] = If987109479436b8d51629513310a948d;
assign I6a91c509b367469511d65174ad4e3b44 = I988e525020c1e43d238fad41dab4e6ea[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[51] = I6a91c509b367469511d65174ad4e3b44;
assign Ib0fc75acbd769930a34393612c6f4fca = I90d92887cb2526a2956d5e8c9fad760c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[52] = Ib0fc75acbd769930a34393612c6f4fca;
assign Ie9ac51d5e0f07e135eb10651d94829d4 = I00fe3792cde1eeab36e576fd6634c4fa[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[53] = Ie9ac51d5e0f07e135eb10651d94829d4;
assign I6faf08de30d6ba38e76cbf7c868a6f73 = I6e586c5ac59a28b30c377e51287bf04d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[54] = I6faf08de30d6ba38e76cbf7c868a6f73;
assign I6a5a58a73d0557e080e6327ee386020b = Ib5dc74106d8841d25a793010fdac599a[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[55] = I6a5a58a73d0557e080e6327ee386020b;
assign I3704ac8ccceb7a319344229dc2db6693 = I3eaf142d2734d2d0decef084dc037b50[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[56] = I3704ac8ccceb7a319344229dc2db6693;
assign Iebedd8e3b4af888431e0a294d56c5c9f = I2d171ad83e27a3745d204849a6f46954[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[57] = Iebedd8e3b4af888431e0a294d56c5c9f;
assign I7bc366f56c020144390350e85747a6f6 = I977f1083f5e4f6f8ac38e2c5aecf1b79[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[58] = I7bc366f56c020144390350e85747a6f6;
assign Ia3252e7c4f3897ef6637bd063b00d3c6 = I9bcd673a4293e14fd20b48fa20492df7[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[59] = Ia3252e7c4f3897ef6637bd063b00d3c6;
assign Id135567b50e17e28d140be2906bfe185 = Icb7422ea46b22b9330c123b40fe343fe[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[60] = Id135567b50e17e28d140be2906bfe185;
assign I3e5c9230c5b091b31ec13fddaea37a8f = Ic414cdba230d7ea73972b0eda1ec6b1b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[61] = I3e5c9230c5b091b31ec13fddaea37a8f;
assign I1c3a83518d660eb2549b1b8d2a2f6186 = Ie4e1e00503dba189b0f871c3c0810d76[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[62] = I1c3a83518d660eb2549b1b8d2a2f6186;
assign I86e509fc0160543f825aefa4dea4eaf4 = I721c43ab62b42a18c3f5228fc0a73262[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[63] = I86e509fc0160543f825aefa4dea4eaf4;
assign I6cb732a94dbf7bed4e70f4b6a1c393f1 = I1f7cb03cf806b247be1cace4d75de942[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[64] = I6cb732a94dbf7bed4e70f4b6a1c393f1;
assign I0d3ce639167582d0b25085ff5b98f7c4 = I775cc766b069022bc00220050feee4e4[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[65] = I0d3ce639167582d0b25085ff5b98f7c4;
assign I7f786778e022e1cba9aa7032c0d43db9 = I08b78f774ed494fa7f119977bd92679e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[66] = I7f786778e022e1cba9aa7032c0d43db9;
assign I4722e6750746bbe43018b591688ac3e9 = Ic7dc7f94af108ca7c8003a2d07e1e168[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[67] = I4722e6750746bbe43018b591688ac3e9;
assign Ie320d1535571a2af4ec61057258a60b6 = Ibe1327961152cc2d26b3f19476a6e2c9[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[68] = Ie320d1535571a2af4ec61057258a60b6;
assign I69c88d14b5244f55911e23f7685f37d0 = I5ba97de444af4e8c9744c3b707502edc[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[69] = I69c88d14b5244f55911e23f7685f37d0;
assign Icbb724c2e16e099c0820935ac4fe21e7 = I3e4f1314042010b5d7384693b580da7b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[70] = Icbb724c2e16e099c0820935ac4fe21e7;
assign I01b9e488ff0277a2e1e8b52004e4cbd3 = I4a47ce6e21c1a274578397e480c184c9[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[71] = I01b9e488ff0277a2e1e8b52004e4cbd3;
assign If329f0c1b6d206280da518bedeb1b5c3 = Id184731beb200ad6a53ce273b963bb3e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[72] = If329f0c1b6d206280da518bedeb1b5c3;
assign I47e322cc161d674131f11ca70479c538 = I3317f2f6eef9a8ef1fe1ff68b47c5d03[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[73] = I47e322cc161d674131f11ca70479c538;
assign Ib343e5b8ebe704ab55692f487b06c156 = Ia6b9fa10c79e6f3847f89b35afb4cc59[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[74] = Ib343e5b8ebe704ab55692f487b06c156;
assign I1a6bc8e0684efd6ea5f73651688f9cc6 = I91e98b804ef82eea53c5e8eccfec827f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[75] = I1a6bc8e0684efd6ea5f73651688f9cc6;
assign Ief7890423e793f41bf2b9f27ff47b4a3 = I5f1e0d0c6b50f70a6f5584124e095501[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[76] = Ief7890423e793f41bf2b9f27ff47b4a3;
assign I145a313064c4d2c5c30fd9458bd32d56 = Id61fcc605b4b581f5d42024c2610c8b7[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[77] = I145a313064c4d2c5c30fd9458bd32d56;
assign I2dfaa00d2d1869026f6c8651ad8cfde9 = Id64738b7668931553151dbadd5605b71[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[78] = I2dfaa00d2d1869026f6c8651ad8cfde9;
assign Ief703cb630f99bc2d59ae0e27bfb3572 = I3bdfb451eb96d256da542864d39024df[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[79] = Ief703cb630f99bc2d59ae0e27bfb3572;
assign I3c5c01afc7096f90c8c6f875dd9686b0 = Ia740d8ccd8230b28d078b2ea3e58d6ba[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[80] = I3c5c01afc7096f90c8c6f875dd9686b0;
assign I5ec91f70ba0346f55caacb7e78f714d4 = I574050722f82569d34bc2cfae1eedaa9[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[81] = I5ec91f70ba0346f55caacb7e78f714d4;
assign Iccf8ad1402095a65a32897af9d8ce23b = Ic8f7ec6ee09fb9ee2467e3cea30a44a3[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[82] = Iccf8ad1402095a65a32897af9d8ce23b;
assign I18950ce49f50b9fd4aa6b1d69b162fe6 = I2b77d922a74fdcef0d57debc789bd539[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[83] = I18950ce49f50b9fd4aa6b1d69b162fe6;
assign I6ad8cf59d777a2e6832471a2cb713eb3 = Ia1d8127af4944b23475bd7deac91d60e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[84] = I6ad8cf59d777a2e6832471a2cb713eb3;
assign I8d24e40d6e2c96260bb58024eb57765d = I247abcede9914633c0a33fc402bf58ae[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[85] = I8d24e40d6e2c96260bb58024eb57765d;
assign I7ebb24e284f0aeb792723e15024fdd7b = I1f413d3e081c6aea012b122fc94f73d5[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[86] = I7ebb24e284f0aeb792723e15024fdd7b;
assign I717cc8e9bb50878c67c3cef72088f279 = I1b812fb764d3b48511c0d15a7efaea29[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[87] = I717cc8e9bb50878c67c3cef72088f279;
assign I9140c28397eaeffd7a3446096bbb8419 = I88882bd8a9f8718411564221ad85b223[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[88] = I9140c28397eaeffd7a3446096bbb8419;
assign I1563ae311393b429f4fe42180f1c61a4 = I232f24e2798488ee66003f3b8cc294c0[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[89] = I1563ae311393b429f4fe42180f1c61a4;
assign I068dc4e9969e691dec22979b38ee588e = I856284e951773518eb6c4232ea7f3d40[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[90] = I068dc4e9969e691dec22979b38ee588e;
assign I9820fcf4305469c0390cf04be00ddf1b = I82cbeaf5b3e4796b2aaf33dcbd119f4f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[91] = I9820fcf4305469c0390cf04be00ddf1b;
assign I24a3a82a62c3c1348663e84e1d80de10 = Iaa7791bbc193412e5fe25000ceec23d6[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[92] = I24a3a82a62c3c1348663e84e1d80de10;
assign I10b2505a209c84c3468bf8c5564ff7b2 = I44bdc0baed3d51ef54ce2728618ad339[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[93] = I10b2505a209c84c3468bf8c5564ff7b2;
assign Iac33806e51f5fcf8e571bfa02272151e = Ib6bc7e75ce750a26113cbb8895c2f024[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[94] = Iac33806e51f5fcf8e571bfa02272151e;
assign Ib0f7718835e96a6b3ce6e7eacc5ae37b = Ib4188380f7e96d5afb99f5045674193d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[95] = Ib0f7718835e96a6b3ce6e7eacc5ae37b;
assign I68bcde39ac1f26fa5c8daa7e616b7924 = I5bba219c5024301e420e9a5acbdc5845[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[96] = I68bcde39ac1f26fa5c8daa7e616b7924;
assign Ia320bdbc669ece554e4dcac16a650551 = I1bb52988c9ba03e16b1b69335d3d7e7c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[97] = Ia320bdbc669ece554e4dcac16a650551;
assign Ic31b8782fe7655bf0dbbbc034acaf00c = I1b9990aaeae716f66b0f89fb02be0a74[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[98] = Ic31b8782fe7655bf0dbbbc034acaf00c;
assign I7f1175afac88a045954988d97e6c014a = Iceec2cf6aba9138648a3340390f39fe9[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[99] = I7f1175afac88a045954988d97e6c014a;
assign I2aec42e2d6c3389d51b99855f4b31413 = Iad7842f3d4672f42c1064c28d4c8ec4e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[100] = I2aec42e2d6c3389d51b99855f4b31413;
assign If6053e257420db5a04d9864730adcb98 = Ie5a53cf9343fdcdb5788667c45fadc83[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[101] = If6053e257420db5a04d9864730adcb98;
assign I107da1e40d1217df6353e403066bacc2 = I30e06d190906bc9eb6f1c3156c47f9f1[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[102] = I107da1e40d1217df6353e403066bacc2;
assign Idb29269890e208fbac5a370a883f180d = Ieaaaced47e22029ad2945eac9cc45e6c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[103] = Idb29269890e208fbac5a370a883f180d;
assign I5ca6297084710e3fc6d343511e4c8e42 = I08dc6f8e837b1f6b80bd3fc742290dab[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[104] = I5ca6297084710e3fc6d343511e4c8e42;
assign I586b30878699ef8f0d09e922262a19d4 = I8eb6a9c907c5909dad6cda98022d70b8[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[105] = I586b30878699ef8f0d09e922262a19d4;
assign I2a833dfb485a2a420a799ef5854b1dee = Ia5067b1b458af82c3c2cd50653099854[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[106] = I2a833dfb485a2a420a799ef5854b1dee;
assign I598ba40aca3b048d684323016e46c777 = I198c6753cf12d423c709d1512e66fa9b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[107] = I598ba40aca3b048d684323016e46c777;
assign Idfe3a41188b5115db103d16bf7b4417b = Ib600dd8a39fda48d28e1289d44d49a84[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[108] = Idfe3a41188b5115db103d16bf7b4417b;
assign I7679c765ab544db47fae6a7867974d61 = Iabf09191227584c76d7fbc634b706d12[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[109] = I7679c765ab544db47fae6a7867974d61;
assign I30afde55f450fcb898f5854004d618e9 = I4869ba08cab90a6dcbc454b0001a7a20[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[110] = I30afde55f450fcb898f5854004d618e9;
assign Ic216abe8348824570dce569f4ff9d186 = If97974406672507f8c9a1c507c4b6951[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[111] = Ic216abe8348824570dce569f4ff9d186;
assign Ieb0dc034a1be9a5d3f2919b4d00d0960 = I4210341f99ac7cb08245137999739114[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[112] = Ieb0dc034a1be9a5d3f2919b4d00d0960;
assign Ia4a51f9d6b4d72bc7edc29acc1938b67 = Ic24f4dbd99c8f4d88c8450d4fef762b8[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[113] = Ia4a51f9d6b4d72bc7edc29acc1938b67;
assign I83757c2cdf0e4516bdafb5f6b4760aa3 = I68dffa1a13eb6ab54615347729c1d6af[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[114] = I83757c2cdf0e4516bdafb5f6b4760aa3;
assign I949a414f7676d024a216b21e3d1a9cac = I10153d5548b184b9ac2cecdba4ec4b1a[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[115] = I949a414f7676d024a216b21e3d1a9cac;
assign Ifa3590aff64fc8ef90046c547e6e6f88 = I104b7f0512440cffc0fcce25e477f537[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[116] = Ifa3590aff64fc8ef90046c547e6e6f88;
assign I133c6136e389a5bee5a3006d939a0a6c = I18b6758319272eebbe76e1eee5ae55b2[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[117] = I133c6136e389a5bee5a3006d939a0a6c;
assign I4b615d38e855bc21d809e3e5b24732b7 = I780263b10b98f9bb0eaf66c045d8d37c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[118] = I4b615d38e855bc21d809e3e5b24732b7;
assign Ib8e420738c31144696b4cf90eb99e270 = I37b772442e55cbcd44ba892a0608d662[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[119] = Ib8e420738c31144696b4cf90eb99e270;
assign I09a993ba748562fb5ca4df9f36f683e6 = I0ac256a6659ff5c6673fd110a8bf578f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[120] = I09a993ba748562fb5ca4df9f36f683e6;
assign Ida3263e09545600a85caf500b5cba32d = If134e1d27e736005e5a390e7a2ea1f4b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[121] = Ida3263e09545600a85caf500b5cba32d;
assign I55f6d7a4bbd8422555543abe0171d576 = I7b37b8f908cd82683832536e02faab0d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[122] = I55f6d7a4bbd8422555543abe0171d576;
assign I9fa0e35a8ecacfa315845aeb73ccbab3 = I08b4bf60c9c7e7229bd1952cc88bc7b3[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[123] = I9fa0e35a8ecacfa315845aeb73ccbab3;
assign Ifdcee23865377289dc0e9986c92325be = I267d637eb63fef9f4723f7978fad88f0[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[124] = Ifdcee23865377289dc0e9986c92325be;
assign Ic8ccb35ab31c6d17b98e5f63c022d187 = I4fb56a70e5ffa71f58f715da36368e04[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[125] = Ic8ccb35ab31c6d17b98e5f63c022d187;
assign Ibfaf924a5a317dbcc967127e153d56ba = I5e9e2acb258baf96ac4b525bba54a462[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[126] = Ibfaf924a5a317dbcc967127e153d56ba;
assign Iedabfd30e25648ea4e62808e1922f016 = Ic40f61443a4d8f87769067fc39381cb3[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[127] = Iedabfd30e25648ea4e62808e1922f016;
assign I437ac9b58f5e248aebec968c948c4125 = Ieb36710c9a3726f33407436d62639c8d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[128] = I437ac9b58f5e248aebec968c948c4125;
assign I0cef2090a761574041a230f80dfce8f9 = Ic804af393da2e4b9c8ef25d4a3b4e8d5[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[129] = I0cef2090a761574041a230f80dfce8f9;
assign Ie25a0d7f0c4b7b25ecffa8af65866f60 = I52e4c446693c29a42bb3b665f72d382d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[130] = Ie25a0d7f0c4b7b25ecffa8af65866f60;
assign Id33e269cf9da206ef2c24e1eb4a1184a = Idbf02cf10add496d30fa44bbb18458c6[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[131] = Id33e269cf9da206ef2c24e1eb4a1184a;
assign I9d21b9384524b55c2eb70826c045052f = Ida095585ad26e215f1c1bf989912da89[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[132] = I9d21b9384524b55c2eb70826c045052f;
assign I1332e87f7d43cae554ff461d3957edb9 = I19f1ffa05c7c9a0df5e7014044024c7b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[133] = I1332e87f7d43cae554ff461d3957edb9;
assign Ie11bc6b5b26c889cf8d2236c17f9ca98 = I4d68a2fe778fa93faac38b138138291f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[134] = Ie11bc6b5b26c889cf8d2236c17f9ca98;
assign If1cf7892a4b06f5e88f3831ba6bcecc8 = I54393ada6f76ac82c31f2668e228e29d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[135] = If1cf7892a4b06f5e88f3831ba6bcecc8;
assign I76a07c1dc9d6d51fe3a31ea3a58ef916 = If5b9ef84f09680f3593250b13a852c1c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[136] = I76a07c1dc9d6d51fe3a31ea3a58ef916;
assign Ia51886b7fca8fc0eda0b93c40d8ccc64 = Ibb759bc4179e5b7aa759d850c7cfa467[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[137] = Ia51886b7fca8fc0eda0b93c40d8ccc64;
assign I48c3c239dfc925169c61fae6fcd16eba = I05e8b5f8b83f07b609b5ebf272bb2229[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[138] = I48c3c239dfc925169c61fae6fcd16eba;
assign I87a5898180c3b4934fa6d4832b6507d5 = If6ac15373ec1146d38e7aeb71c3ece64[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[139] = I87a5898180c3b4934fa6d4832b6507d5;
assign I18279e41940f794e7bfcca8062c42ee1 = I2ab3675e1eede757af80716ba980a4e6[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[140] = I18279e41940f794e7bfcca8062c42ee1;
assign I04cc6e9d889d548aed3e517b1c7a98a4 = I388c271687ab31b57421ad57192273ed[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[141] = I04cc6e9d889d548aed3e517b1c7a98a4;
assign I5b319b9f50e43a7c850594b015d24ef8 = I6121679cec8caa51dc5ff0d1a61f9821[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[142] = I5b319b9f50e43a7c850594b015d24ef8;
assign Idad08f7167bd930530e12f9180bd576a = Ia0649b990bf5716cfab230127cd5d47f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[143] = Idad08f7167bd930530e12f9180bd576a;
assign I044b9326d592e52c74056c2385d9a07b = I867a0626ca22108b16267d95c0aadf4f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[144] = I044b9326d592e52c74056c2385d9a07b;
assign I838a7c657b5ddc47cce2b9fcbd433548 = I1af54bcb73d7c6b93e55450871207976[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[145] = I838a7c657b5ddc47cce2b9fcbd433548;
assign Icf019d30479d47cec2a9508e6ac4882e = I91883553543d0425e9c6dd726dce3d27[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[146] = Icf019d30479d47cec2a9508e6ac4882e;
assign I344dd9d785b1ec8f6c3a0d8fc1f400f5 = Ie95405659701278e3f87bf1f823a037b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[147] = I344dd9d785b1ec8f6c3a0d8fc1f400f5;
assign I380dd5278a22dbf0fd4b86985f91dd6b = Ia42392e2104b50c0908aad82738a5ee7[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[148] = I380dd5278a22dbf0fd4b86985f91dd6b;
assign I5feb2a46a916f5ed44638712d5ecc3a6 = I68ad63230a51b9b9e3daffb307ea970d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[149] = I5feb2a46a916f5ed44638712d5ecc3a6;
assign Ib184353aaeae5ef036ff36d0bd35a27f = I7a052d63944ccf42e598efe3a95b88f8[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[150] = Ib184353aaeae5ef036ff36d0bd35a27f;
assign I53729ddbc242ad9a8724d93648868db6 = I2b3c6d69f79c8d51e4d1614c62c44fcc[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[151] = I53729ddbc242ad9a8724d93648868db6;
assign I6429512833e3251e949ad734bfb1dbfa = Ifcef0e92f50e3920bf1208af5d64c632[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[152] = I6429512833e3251e949ad734bfb1dbfa;
assign I96babc82431ae1d3713786eb68c2e372 = I111340a19625901a3c1b95fd0bd1570e[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[153] = I96babc82431ae1d3713786eb68c2e372;
assign Id76e3859fce7aab300a173587243b0a9 = I11aec4fa85c30f6fe1fd9fa72542ef6c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[154] = Id76e3859fce7aab300a173587243b0a9;
assign Ie607dd51fbd545d298488a6e9c9430c6 = I80cc333c181c16a96b7bd6501c27c2b3[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[155] = Ie607dd51fbd545d298488a6e9c9430c6;
assign I00e222e2e16487cfbac6206d913ebc21 = Idc6354325a6280ae9890da33c06c33ec[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[156] = I00e222e2e16487cfbac6206d913ebc21;
assign I400dac72f25c87765a07e72c3d04240e = Ibb04cf82acc4ac16599ad3ddb0c2ada2[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[157] = I400dac72f25c87765a07e72c3d04240e;
assign Ib0b26ab3c5d3109999c55b41e8399c4e = I3ed096dfd8a14f4acb4d53a70cf8aceb[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[158] = Ib0b26ab3c5d3109999c55b41e8399c4e;
assign Ibd55c6f55d6481b76591e2c565217e4c = I0fa07f95e96326cb0599c0c3f76e2b48[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[159] = Ibd55c6f55d6481b76591e2c565217e4c;
assign Ie5764d99afa00cd108404de18693c4c9 = I87d98fbc97d9a78c2e7d6a6280e7a49a[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[160] = Ie5764d99afa00cd108404de18693c4c9;
assign I5234341950ae6353868b35e84b0d837b = Ib7ddc4dca877f7cf5697a02c3d1915ba[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[161] = I5234341950ae6353868b35e84b0d837b;
assign Ice8048703f0f8018353d8666516e2b7d = I3612ef280891f6017fad205d0484bde7[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[162] = Ice8048703f0f8018353d8666516e2b7d;
assign If4ab153a2932d079ae16480dd788d298 = I561547649aeb5b4c3f10d9506db1f3cf[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[163] = If4ab153a2932d079ae16480dd788d298;
assign Iffdd32b08a1072206b9b83981560b341 = I84cc76c0079b86da7b994844c3ccb875[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[164] = Iffdd32b08a1072206b9b83981560b341;
assign Id328a2bf60eddb0da7bc9fe44eb81163 = Iec013c508d0c6401d7eb856e7eb60446[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[165] = Id328a2bf60eddb0da7bc9fe44eb81163;
assign If39c82e97c07c30522a1b489ec896577 = Ifd8979aac6b6b24aa560b46b18240e92[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[166] = If39c82e97c07c30522a1b489ec896577;
assign Id78ace2bd65545c4add80a2720338443 = If12394e78dc913b01890b56650856a44[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[167] = Id78ace2bd65545c4add80a2720338443;
assign I26cd0e322d30abad73493e57d4157954 = I94d18aa10695f3f22b23246884b72822[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[168] = I26cd0e322d30abad73493e57d4157954;
assign I6d27a778e8595666903f4d20d47dc053 = Ic90b38835dd7e760dd54067b196f8470[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[169] = I6d27a778e8595666903f4d20d47dc053;
assign Ic220ac5d53b5c26985e5c7de2d95d896 = If3691ea51f6efe9b165a31964854d2fe[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[170] = Ic220ac5d53b5c26985e5c7de2d95d896;
assign I9793ca0ff4f0324792cbb1da51d60904 = Ic2ce582555add38a14f5006d3c87eb15[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[171] = I9793ca0ff4f0324792cbb1da51d60904;
assign I76b19931a9589b4658dda1384f13f30f = I58cc950ee2cbe56b7c5a619be3792511[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[172] = I76b19931a9589b4658dda1384f13f30f;
assign I0726346b2914d4aeb149e512d31af95f = I0d8e329ec5873db96df1ec309445a096[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[173] = I0726346b2914d4aeb149e512d31af95f;
assign I399c5a08f19fda00d218b1fe4376eb5b = I106325488e2ecfdba1cf9e5201e6bc8c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[174] = I399c5a08f19fda00d218b1fe4376eb5b;
assign I7c3e36e47bc35c16a8420d88b356e9e1 = Iff73a0085541a511d3912b64686a82c5[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[175] = I7c3e36e47bc35c16a8420d88b356e9e1;
assign Ia0bc5e9d76d19f62b221c666f533d959 = Icdab59de68f2870504598c9ea18f1d2c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[176] = Ia0bc5e9d76d19f62b221c666f533d959;
assign I366301d215cb0f4bc390aa6a5726d86b = I75604d727e82c977741f90113719183a[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[177] = I366301d215cb0f4bc390aa6a5726d86b;
assign Id039bdeb594da7428838b1dc4d6af8c2 = I6f50c4d0d2639857b2dcca300c2d7b04[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[178] = Id039bdeb594da7428838b1dc4d6af8c2;
assign I2df05059b08aa3babba9542b51367c83 = I5cd013a2be2e761c10c6a957632517de[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[179] = I2df05059b08aa3babba9542b51367c83;
assign Ia0a811eaed4d73f4012e1fb6217cbda2 = Iafeedddd02428bd2610c576e68d4ae25[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[180] = Ia0a811eaed4d73f4012e1fb6217cbda2;
assign I43333dfaf1cd037fd6bc16d290e0ea86 = I912d6325e34180e0f668f0f024e63581[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[181] = I43333dfaf1cd037fd6bc16d290e0ea86;
assign I4a7337b53c190d757d250223ede3daf3 = Id1e05294dfd02df499ad0c08bb5c191b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[182] = I4a7337b53c190d757d250223ede3daf3;
assign I49d3d7a17c12933457f26c5232277395 = Id3bb9b100ee4302473b49ac14615e9b0[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[183] = I49d3d7a17c12933457f26c5232277395;
assign Ife2b1721d683a43be53c43e49d96e0f5 = Ief32db1cfc443119b6202b0cc7bf70a2[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[184] = Ife2b1721d683a43be53c43e49d96e0f5;
assign Iecf2a3bbabca3f1ee3c9bbc3ea3d2083 = Iad7dbe9909b5eed3261adf92d3813acc[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[185] = Iecf2a3bbabca3f1ee3c9bbc3ea3d2083;
assign I388f3758e343ea6ee2ca6c14a6a8afac = Ie7daf0789c35caaadbba06cafabd2b70[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[186] = I388f3758e343ea6ee2ca6c14a6a8afac;
assign I70754064855cd8d49164f5a24c2087e7 = I2bd1f9b75d9ab94af9ddceb7528935e8[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[187] = I70754064855cd8d49164f5a24c2087e7;
assign I9443c16fdec0687f97a3fe287787e4b9 = Ic3d9f5c6677758810e4865779ec303e3[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[188] = I9443c16fdec0687f97a3fe287787e4b9;
assign I5d871bf470d68cb1651c695f14a2dcb7 = I00af04882a25e2832d913a67d4d86d7b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[189] = I5d871bf470d68cb1651c695f14a2dcb7;
assign I30a21066d0f7ad97b21dfdcc42fe3aee = Ic9db631df0a1a9108c10c3e0eca7bf15[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[190] = I30a21066d0f7ad97b21dfdcc42fe3aee;
assign If0cb066c4e37fd6772da2ee943543829 = I749f9ed1fb2dddd40ebc28f638e02935[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[191] = If0cb066c4e37fd6772da2ee943543829;
assign Idf3132bae12e52ed9560eac88e2ead65 = Ia45b2a24df24bd5e3c95885c8928686c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[192] = Idf3132bae12e52ed9560eac88e2ead65;
assign If092511da36f3f493f7e3f34a35cb9eb = I7427464fde340780aba7f9847b4ad564[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[193] = If092511da36f3f493f7e3f34a35cb9eb;
assign Ice07207e1867f71dbb58dc0b3d28f5d1 = I33fd1ae225e2b881b2b41e0358675e22[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[194] = Ice07207e1867f71dbb58dc0b3d28f5d1;
assign Id1c6ccb54bf2d0d03f296cbd502fac6a = I2e21a35d1cf560936fd19b944a208b6b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[195] = Id1c6ccb54bf2d0d03f296cbd502fac6a;
assign I7a2b0491133ed6a2daafb889ff46d271 = I249522a3d42cc75d7a6b9ede1222ee76[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[196] = I7a2b0491133ed6a2daafb889ff46d271;
assign I4fabd40b7afb192a9c2a255512fd0852 = I68b4c43d9f40ae4bfd70d2983594392c[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[197] = I4fabd40b7afb192a9c2a255512fd0852;
assign I7b39e709a6939751b11bb3ba6fc42bde = I63145e0fec15c7e7c0de105f348bfd31[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[198] = I7b39e709a6939751b11bb3ba6fc42bde;
assign I3a7a76b3ca144951bb6edeba1650c35a = I8af625de86c04016c3424d116fddab5b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[199] = I3a7a76b3ca144951bb6edeba1650c35a;
assign I3c023a3a1a2ce2fb54b2292401df0019 = I54c9c10527f83b4ee4e1e22f1e4044ed[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[200] = I3c023a3a1a2ce2fb54b2292401df0019;
assign I804cf7b8b79a124cbee51fe473e664a3 = I972559e47c7f83bd9000ca1cfc14d8e0[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[201] = I804cf7b8b79a124cbee51fe473e664a3;
assign I33be2a0d4c64f50472091a4503281558 = Ib97a7f941eb7ce2a867503a04ff86a67[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[202] = I33be2a0d4c64f50472091a4503281558;
assign Ie5f94955ed10ae50d92d3dd0e43c8088 = I5979b55f607c71017537f2b48b40cbea[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[203] = Ie5f94955ed10ae50d92d3dd0e43c8088;
assign Ide6f35e8581e1bec17ec974448b6beed = I6a56760b621f238843b091279c69897f[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[204] = Ide6f35e8581e1bec17ec974448b6beed;
assign I57b47b934005413e4c400a33e7ddc20c = Icec45bf76c241d37c9a50a5cd092da9d[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[205] = I57b47b934005413e4c400a33e7ddc20c;
assign Id4e7f9a0c100dfc591e7693d76a496d9 = I2f6d3f61f2890e584d3063a09587e99b[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[206] = Id4e7f9a0c100dfc591e7693d76a496d9;
assign Ieda30691eb70678f7535eed71e9ee031 = I7c396ea2e959d84fd9a6964617cb29c6[SGN_MAX_SUM_WDTH_P1]; //valid Ied2b5c0139cec8ad2873829dc1117d50 d7
assign final_y_nr_dec[207] = Ieda30691eb70678f7535eed71e9ee031;

   always @(posedge clk or negedge rstn)
   begin
       if (!rstn) begin

// Ie4894ca167b08880bfc35862f18575eb Ied2b5c0139cec8ad2873829dc1117d50 I05531b19bb846b18c09f979eeb429ad3 Ibd047e2643dc68affb5b4f25b82ded31 valid Ied2b5c0139cec8ad2873829dc1117d50 Ibd047e2643dc68affb5b4f25b82ded31
          tmp_bit[0]  <=   0;
          tmp_bit[1]  <=   0;
          tmp_bit[2]  <=   0;
          tmp_bit[3]  <=   0;
          tmp_bit[4]  <=   0;
          tmp_bit[5]  <=   0;
          tmp_bit[6]  <=   0;
          tmp_bit[7]  <=   0;
          tmp_bit[8]  <=   0;
          tmp_bit[9]  <=   0;
          tmp_bit[10]  <=   0;
          tmp_bit[11]  <=   0;
          tmp_bit[12]  <=   0;
          tmp_bit[13]  <=   0;
          tmp_bit[14]  <=   0;
          tmp_bit[15]  <=   0;
          tmp_bit[16]  <=   0;
          tmp_bit[17]  <=   0;
          tmp_bit[18]  <=   0;
          tmp_bit[19]  <=   0;
          tmp_bit[20]  <=   0;
          tmp_bit[21]  <=   0;
          tmp_bit[22]  <=   0;
          tmp_bit[23]  <=   0;
          tmp_bit[24]  <=   0;
          tmp_bit[25]  <=   0;
          tmp_bit[26]  <=   0;
          tmp_bit[27]  <=   0;
          tmp_bit[28]  <=   0;
          tmp_bit[29]  <=   0;
          tmp_bit[30]  <=   0;
          tmp_bit[31]  <=   0;
          tmp_bit[32]  <=   0;
          tmp_bit[33]  <=   0;
          tmp_bit[34]  <=   0;
          tmp_bit[35]  <=   0;
          tmp_bit[36]  <=   0;
          tmp_bit[37]  <=   0;
          tmp_bit[38]  <=   0;
          tmp_bit[39]  <=   0;
          tmp_bit[40]  <=   0;
          tmp_bit[41]  <=   0;
          tmp_bit[42]  <=   0;
          tmp_bit[43]  <=   0;
          tmp_bit[44]  <=   0;
          tmp_bit[45]  <=   0;
          tmp_bit[46]  <=   0;
          tmp_bit[47]  <=   0;
          tmp_bit[48]  <=   0;
          tmp_bit[49]  <=   0;
          tmp_bit[50]  <=   0;
          tmp_bit[51]  <=   0;
          tmp_bit[52]  <=   0;
          tmp_bit[53]  <=   0;
          tmp_bit[54]  <=   0;
          tmp_bit[55]  <=   0;
          tmp_bit[56]  <=   0;
          tmp_bit[57]  <=   0;
          tmp_bit[58]  <=   0;
          tmp_bit[59]  <=   0;
          tmp_bit[60]  <=   0;
          tmp_bit[61]  <=   0;
          tmp_bit[62]  <=   0;
          tmp_bit[63]  <=   0;
          tmp_bit[64]  <=   0;
          tmp_bit[65]  <=   0;
          tmp_bit[66]  <=   0;
          tmp_bit[67]  <=   0;
          tmp_bit[68]  <=   0;
          tmp_bit[69]  <=   0;
          tmp_bit[70]  <=   0;
          tmp_bit[71]  <=   0;
          tmp_bit[72]  <=   0;
          tmp_bit[73]  <=   0;
          tmp_bit[74]  <=   0;
          tmp_bit[75]  <=   0;
          tmp_bit[76]  <=   0;
          tmp_bit[77]  <=   0;
          tmp_bit[78]  <=   0;
          tmp_bit[79]  <=   0;
          tmp_bit[80]  <=   0;
          tmp_bit[81]  <=   0;
          tmp_bit[82]  <=   0;
          tmp_bit[83]  <=   0;
          tmp_bit[84]  <=   0;
          tmp_bit[85]  <=   0;
          tmp_bit[86]  <=   0;
          tmp_bit[87]  <=   0;
          tmp_bit[88]  <=   0;
          tmp_bit[89]  <=   0;
          tmp_bit[90]  <=   0;
          tmp_bit[91]  <=   0;
          tmp_bit[92]  <=   0;
          tmp_bit[93]  <=   0;
          tmp_bit[94]  <=   0;
          tmp_bit[95]  <=   0;
          tmp_bit[96]  <=   0;
          tmp_bit[97]  <=   0;
          tmp_bit[98]  <=   0;
          tmp_bit[99]  <=   0;
          tmp_bit[100]  <=   0;
          tmp_bit[101]  <=   0;
          tmp_bit[102]  <=   0;
          tmp_bit[103]  <=   0;
          tmp_bit[104]  <=   0;
          tmp_bit[105]  <=   0;
          tmp_bit[106]  <=   0;
          tmp_bit[107]  <=   0;
          tmp_bit[108]  <=   0;
          tmp_bit[109]  <=   0;
          tmp_bit[110]  <=   0;
          tmp_bit[111]  <=   0;
          tmp_bit[112]  <=   0;
          tmp_bit[113]  <=   0;
          tmp_bit[114]  <=   0;
          tmp_bit[115]  <=   0;
          tmp_bit[116]  <=   0;
          tmp_bit[117]  <=   0;
          tmp_bit[118]  <=   0;
          tmp_bit[119]  <=   0;
          tmp_bit[120]  <=   0;
          tmp_bit[121]  <=   0;
          tmp_bit[122]  <=   0;
          tmp_bit[123]  <=   0;
          tmp_bit[124]  <=   0;
          tmp_bit[125]  <=   0;
          tmp_bit[126]  <=   0;
          tmp_bit[127]  <=   0;
          tmp_bit[128]  <=   0;
          tmp_bit[129]  <=   0;
          tmp_bit[130]  <=   0;
          tmp_bit[131]  <=   0;
          tmp_bit[132]  <=   0;
          tmp_bit[133]  <=   0;
          tmp_bit[134]  <=   0;
          tmp_bit[135]  <=   0;
          tmp_bit[136]  <=   0;
          tmp_bit[137]  <=   0;
          tmp_bit[138]  <=   0;
          tmp_bit[139]  <=   0;
          tmp_bit[140]  <=   0;
          tmp_bit[141]  <=   0;
          tmp_bit[142]  <=   0;
          tmp_bit[143]  <=   0;
          tmp_bit[144]  <=   0;
          tmp_bit[145]  <=   0;
          tmp_bit[146]  <=   0;
          tmp_bit[147]  <=   0;
          tmp_bit[148]  <=   0;
          tmp_bit[149]  <=   0;
          tmp_bit[150]  <=   0;
          tmp_bit[151]  <=   0;
          tmp_bit[152]  <=   0;
          tmp_bit[153]  <=   0;
          tmp_bit[154]  <=   0;
          tmp_bit[155]  <=   0;
          tmp_bit[156]  <=   0;
          tmp_bit[157]  <=   0;
          tmp_bit[158]  <=   0;
          tmp_bit[159]  <=   0;
          tmp_bit[160]  <=   0;
          tmp_bit[161]  <=   0;
          tmp_bit[162]  <=   0;
          tmp_bit[163]  <=   0;
          tmp_bit[164]  <=   0;
          tmp_bit[165]  <=   0;
          tmp_bit[166]  <=   0;
          tmp_bit[167]  <=   0;
          tmp_bit[168]  <=   0;
          tmp_bit[169]  <=   0;
          tmp_bit[170]  <=   0;
          tmp_bit[171]  <=   0;
          tmp_bit[172]  <=   0;
          tmp_bit[173]  <=   0;
          tmp_bit[174]  <=   0;
          tmp_bit[175]  <=   0;
          tmp_bit[176]  <=   0;
          tmp_bit[177]  <=   0;
          tmp_bit[178]  <=   0;
          tmp_bit[179]  <=   0;
          tmp_bit[180]  <=   0;
          tmp_bit[181]  <=   0;
          tmp_bit[182]  <=   0;
          tmp_bit[183]  <=   0;
          tmp_bit[184]  <=   0;
          tmp_bit[185]  <=   0;
          tmp_bit[186]  <=   0;
          tmp_bit[187]  <=   0;
          tmp_bit[188]  <=   0;
          tmp_bit[189]  <=   0;
          tmp_bit[190]  <=   0;
          tmp_bit[191]  <=   0;
          tmp_bit[192]  <=   0;
          tmp_bit[193]  <=   0;
          tmp_bit[194]  <=   0;
          tmp_bit[195]  <=   0;
          tmp_bit[196]  <=   0;
          tmp_bit[197]  <=   0;
          tmp_bit[198]  <=   0;
          tmp_bit[199]  <=   0;
          tmp_bit[200]  <=   0;
          tmp_bit[201]  <=   0;
          tmp_bit[202]  <=   0;
          tmp_bit[203]  <=   0;
          tmp_bit[204]  <=   0;
          tmp_bit[205]  <=   0;
          tmp_bit[206]  <=   0;
          tmp_bit[207]  <=   0;

       end else begin

// Ie4894ca167b08880bfc35862f18575eb Ied2b5c0139cec8ad2873829dc1117d50 I05531b19bb846b18c09f979eeb429ad3 Ibd047e2643dc68affb5b4f25b82ded31 valid Ied2b5c0139cec8ad2873829dc1117d50 Ibd047e2643dc68affb5b4f25b82ded31
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[0]  <=   I204375b1fcd1f62621b32a06a9dd0bb6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[1]  <=   Ic0ae28dd2fa2d9e0b2a9edaaffd88aff;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[2]  <=   I63323f8807804f4534429d8aeafc7d23;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[3]  <=   Ie8554592e62dd20a36ef79e06af24a22;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[4]  <=   I67458f3b57d906d3626d4e7656049538;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[5]  <=   I523d96cce3a523da8ca8e065aa5d8f64;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[6]  <=   I3fad2338742a91d05694c9bbe0584126;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[7]  <=   Id30ee39232f016f983f45208ed802126;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[8]  <=   I149dbd0f3f68786fc3a842bb0064f0d4;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[9]  <=   Ib383a8f851cd16df009c975ec7efb305;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[10]  <=   Ia2227bb2140f18af451ea4c397262178;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[11]  <=   Idf0b6d7bfa5a9a38e1362c4b3b0d5b99;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[12]  <=   Iaa15139339207505f231f71669ce022a;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[13]  <=   Idc30dece6bd74ad2ff6c0822347a800d;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[14]  <=   I7492572ef50294af38fc778e173a60fc;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[15]  <=   I4c6718b74573391494789da2e33c1e2d;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[16]  <=   I03659b77af3e47129d9206af314ec521;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[17]  <=   If0fbb2a55965bb66cfaad70fd9241456;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[18]  <=   I4f8bea1f3f8cb9ff1b6d1388c6377861;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[19]  <=   I765559024522a12448e338401c10f800;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[20]  <=   I815daf68a1ed9f91b02ede68298cc5f3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[21]  <=   If0e526189886cb9e8af7be4797d8a637;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[22]  <=   Ic8dfeb5746649e88e59887cda08fb62a;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[23]  <=   I0bd3e1beb510558b20c2b4f0f8f20e76;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[24]  <=   I647c8a9b1fd2281c8e129d2cebdd597e;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[25]  <=   I6a803347e6d25dbd012caf725e35c256;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[26]  <=   Icf6deff8d81d69b92659b257bbdb53c7;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[27]  <=   If282e264f908747340e4e4d2022a66fc;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[28]  <=   Ib5ca6dc87c214c3d73b265fa0e242452;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[29]  <=   I3b8dd3a8e7b21202977c976ba687cb7c;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[30]  <=   I4e1743e1634bdb7ad6e8d072e19f0abd;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[31]  <=   I4ccbbd7d8e03a7c7410acaf35ef87608;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[32]  <=   I1848d733a31c474bcb2d3e4b9b736e94;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[33]  <=   I6fb841a6fe0ad7d433f1a182706d6ad6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[34]  <=   Iddb16107d5ce4ef65024a1cd5387dcd1;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[35]  <=   I8eb4596c73d1cb6ae5a783a6582cbffe;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[36]  <=   I014c1931d012f79e954a12e10178f1d9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[37]  <=   I8ad79c41a8896712d7c26d29c0b1e7cf;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[38]  <=   I1b16bbdd1e23bbe571bc7769731a03d8;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[39]  <=   Ib0cea939898e64f9ec4ee41aa3f062fb;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[40]  <=   Ief16fc889b2326a53224b3b60ecc8955;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[41]  <=   I774b99eb9e3c3c98ce6dd3c60df7eff5;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[42]  <=   Ide90044338620a38b90b5877ce0eb52b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[43]  <=   I2271e9b3a663941eed3b939bf80ed2a1;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[44]  <=   Ifc1b458539905b3557d79c94954747c0;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[45]  <=   Ibe27dea48dd30331b9723a1aec226f0f;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[46]  <=   Ic214eae29f89949c797816779332aef2;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[47]  <=   Icd48fe364089e0250b4fee636590fe28;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[48]  <=   I15d7c9e33bce9e3ee1059f73832bb9ad;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[49]  <=   I9514bd70ebe24af7d8bf346ae09219f7;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[50]  <=   If987109479436b8d51629513310a948d;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[51]  <=   I6a91c509b367469511d65174ad4e3b44;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[52]  <=   Ib0fc75acbd769930a34393612c6f4fca;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[53]  <=   Ie9ac51d5e0f07e135eb10651d94829d4;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[54]  <=   I6faf08de30d6ba38e76cbf7c868a6f73;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[55]  <=   I6a5a58a73d0557e080e6327ee386020b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[56]  <=   I3704ac8ccceb7a319344229dc2db6693;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[57]  <=   Iebedd8e3b4af888431e0a294d56c5c9f;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[58]  <=   I7bc366f56c020144390350e85747a6f6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[59]  <=   Ia3252e7c4f3897ef6637bd063b00d3c6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[60]  <=   Id135567b50e17e28d140be2906bfe185;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[61]  <=   I3e5c9230c5b091b31ec13fddaea37a8f;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[62]  <=   I1c3a83518d660eb2549b1b8d2a2f6186;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[63]  <=   I86e509fc0160543f825aefa4dea4eaf4;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[64]  <=   I6cb732a94dbf7bed4e70f4b6a1c393f1;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[65]  <=   I0d3ce639167582d0b25085ff5b98f7c4;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[66]  <=   I7f786778e022e1cba9aa7032c0d43db9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[67]  <=   I4722e6750746bbe43018b591688ac3e9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[68]  <=   Ie320d1535571a2af4ec61057258a60b6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[69]  <=   I69c88d14b5244f55911e23f7685f37d0;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[70]  <=   Icbb724c2e16e099c0820935ac4fe21e7;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[71]  <=   I01b9e488ff0277a2e1e8b52004e4cbd3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[72]  <=   If329f0c1b6d206280da518bedeb1b5c3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[73]  <=   I47e322cc161d674131f11ca70479c538;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[74]  <=   Ib343e5b8ebe704ab55692f487b06c156;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[75]  <=   I1a6bc8e0684efd6ea5f73651688f9cc6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[76]  <=   Ief7890423e793f41bf2b9f27ff47b4a3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[77]  <=   I145a313064c4d2c5c30fd9458bd32d56;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[78]  <=   I2dfaa00d2d1869026f6c8651ad8cfde9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[79]  <=   Ief703cb630f99bc2d59ae0e27bfb3572;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[80]  <=   I3c5c01afc7096f90c8c6f875dd9686b0;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[81]  <=   I5ec91f70ba0346f55caacb7e78f714d4;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[82]  <=   Iccf8ad1402095a65a32897af9d8ce23b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[83]  <=   I18950ce49f50b9fd4aa6b1d69b162fe6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[84]  <=   I6ad8cf59d777a2e6832471a2cb713eb3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[85]  <=   I8d24e40d6e2c96260bb58024eb57765d;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[86]  <=   I7ebb24e284f0aeb792723e15024fdd7b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[87]  <=   I717cc8e9bb50878c67c3cef72088f279;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[88]  <=   I9140c28397eaeffd7a3446096bbb8419;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[89]  <=   I1563ae311393b429f4fe42180f1c61a4;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[90]  <=   I068dc4e9969e691dec22979b38ee588e;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[91]  <=   I9820fcf4305469c0390cf04be00ddf1b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[92]  <=   I24a3a82a62c3c1348663e84e1d80de10;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[93]  <=   I10b2505a209c84c3468bf8c5564ff7b2;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[94]  <=   Iac33806e51f5fcf8e571bfa02272151e;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[95]  <=   Ib0f7718835e96a6b3ce6e7eacc5ae37b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[96]  <=   I68bcde39ac1f26fa5c8daa7e616b7924;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[97]  <=   Ia320bdbc669ece554e4dcac16a650551;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[98]  <=   Ic31b8782fe7655bf0dbbbc034acaf00c;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[99]  <=   I7f1175afac88a045954988d97e6c014a;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[100]  <=   I2aec42e2d6c3389d51b99855f4b31413;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[101]  <=   If6053e257420db5a04d9864730adcb98;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[102]  <=   I107da1e40d1217df6353e403066bacc2;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[103]  <=   Idb29269890e208fbac5a370a883f180d;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[104]  <=   I5ca6297084710e3fc6d343511e4c8e42;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[105]  <=   I586b30878699ef8f0d09e922262a19d4;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[106]  <=   I2a833dfb485a2a420a799ef5854b1dee;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[107]  <=   I598ba40aca3b048d684323016e46c777;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[108]  <=   Idfe3a41188b5115db103d16bf7b4417b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[109]  <=   I7679c765ab544db47fae6a7867974d61;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[110]  <=   I30afde55f450fcb898f5854004d618e9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[111]  <=   Ic216abe8348824570dce569f4ff9d186;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[112]  <=   Ieb0dc034a1be9a5d3f2919b4d00d0960;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[113]  <=   Ia4a51f9d6b4d72bc7edc29acc1938b67;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[114]  <=   I83757c2cdf0e4516bdafb5f6b4760aa3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[115]  <=   I949a414f7676d024a216b21e3d1a9cac;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[116]  <=   Ifa3590aff64fc8ef90046c547e6e6f88;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[117]  <=   I133c6136e389a5bee5a3006d939a0a6c;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[118]  <=   I4b615d38e855bc21d809e3e5b24732b7;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[119]  <=   Ib8e420738c31144696b4cf90eb99e270;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[120]  <=   I09a993ba748562fb5ca4df9f36f683e6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[121]  <=   Ida3263e09545600a85caf500b5cba32d;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[122]  <=   I55f6d7a4bbd8422555543abe0171d576;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[123]  <=   I9fa0e35a8ecacfa315845aeb73ccbab3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[124]  <=   Ifdcee23865377289dc0e9986c92325be;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[125]  <=   Ic8ccb35ab31c6d17b98e5f63c022d187;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[126]  <=   Ibfaf924a5a317dbcc967127e153d56ba;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[127]  <=   Iedabfd30e25648ea4e62808e1922f016;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[128]  <=   I437ac9b58f5e248aebec968c948c4125;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[129]  <=   I0cef2090a761574041a230f80dfce8f9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[130]  <=   Ie25a0d7f0c4b7b25ecffa8af65866f60;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[131]  <=   Id33e269cf9da206ef2c24e1eb4a1184a;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[132]  <=   I9d21b9384524b55c2eb70826c045052f;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[133]  <=   I1332e87f7d43cae554ff461d3957edb9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[134]  <=   Ie11bc6b5b26c889cf8d2236c17f9ca98;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[135]  <=   If1cf7892a4b06f5e88f3831ba6bcecc8;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[136]  <=   I76a07c1dc9d6d51fe3a31ea3a58ef916;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[137]  <=   Ia51886b7fca8fc0eda0b93c40d8ccc64;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[138]  <=   I48c3c239dfc925169c61fae6fcd16eba;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[139]  <=   I87a5898180c3b4934fa6d4832b6507d5;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[140]  <=   I18279e41940f794e7bfcca8062c42ee1;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[141]  <=   I04cc6e9d889d548aed3e517b1c7a98a4;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[142]  <=   I5b319b9f50e43a7c850594b015d24ef8;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[143]  <=   Idad08f7167bd930530e12f9180bd576a;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[144]  <=   I044b9326d592e52c74056c2385d9a07b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[145]  <=   I838a7c657b5ddc47cce2b9fcbd433548;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[146]  <=   Icf019d30479d47cec2a9508e6ac4882e;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[147]  <=   I344dd9d785b1ec8f6c3a0d8fc1f400f5;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[148]  <=   I380dd5278a22dbf0fd4b86985f91dd6b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[149]  <=   I5feb2a46a916f5ed44638712d5ecc3a6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[150]  <=   Ib184353aaeae5ef036ff36d0bd35a27f;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[151]  <=   I53729ddbc242ad9a8724d93648868db6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[152]  <=   I6429512833e3251e949ad734bfb1dbfa;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[153]  <=   I96babc82431ae1d3713786eb68c2e372;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[154]  <=   Id76e3859fce7aab300a173587243b0a9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[155]  <=   Ie607dd51fbd545d298488a6e9c9430c6;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[156]  <=   I00e222e2e16487cfbac6206d913ebc21;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[157]  <=   I400dac72f25c87765a07e72c3d04240e;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[158]  <=   Ib0b26ab3c5d3109999c55b41e8399c4e;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[159]  <=   Ibd55c6f55d6481b76591e2c565217e4c;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[160]  <=   Ie5764d99afa00cd108404de18693c4c9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[161]  <=   I5234341950ae6353868b35e84b0d837b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[162]  <=   Ice8048703f0f8018353d8666516e2b7d;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[163]  <=   If4ab153a2932d079ae16480dd788d298;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[164]  <=   Iffdd32b08a1072206b9b83981560b341;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[165]  <=   Id328a2bf60eddb0da7bc9fe44eb81163;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[166]  <=   If39c82e97c07c30522a1b489ec896577;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[167]  <=   Id78ace2bd65545c4add80a2720338443;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[168]  <=   I26cd0e322d30abad73493e57d4157954;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[169]  <=   I6d27a778e8595666903f4d20d47dc053;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[170]  <=   Ic220ac5d53b5c26985e5c7de2d95d896;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[171]  <=   I9793ca0ff4f0324792cbb1da51d60904;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[172]  <=   I76b19931a9589b4658dda1384f13f30f;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[173]  <=   I0726346b2914d4aeb149e512d31af95f;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[174]  <=   I399c5a08f19fda00d218b1fe4376eb5b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[175]  <=   I7c3e36e47bc35c16a8420d88b356e9e1;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[176]  <=   Ia0bc5e9d76d19f62b221c666f533d959;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[177]  <=   I366301d215cb0f4bc390aa6a5726d86b;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[178]  <=   Id039bdeb594da7428838b1dc4d6af8c2;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[179]  <=   I2df05059b08aa3babba9542b51367c83;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[180]  <=   Ia0a811eaed4d73f4012e1fb6217cbda2;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[181]  <=   I43333dfaf1cd037fd6bc16d290e0ea86;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[182]  <=   I4a7337b53c190d757d250223ede3daf3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[183]  <=   I49d3d7a17c12933457f26c5232277395;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[184]  <=   Ife2b1721d683a43be53c43e49d96e0f5;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[185]  <=   Iecf2a3bbabca3f1ee3c9bbc3ea3d2083;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[186]  <=   I388f3758e343ea6ee2ca6c14a6a8afac;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[187]  <=   I70754064855cd8d49164f5a24c2087e7;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[188]  <=   I9443c16fdec0687f97a3fe287787e4b9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[189]  <=   I5d871bf470d68cb1651c695f14a2dcb7;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[190]  <=   I30a21066d0f7ad97b21dfdcc42fe3aee;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[191]  <=   If0cb066c4e37fd6772da2ee943543829;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[192]  <=   Idf3132bae12e52ed9560eac88e2ead65;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[193]  <=   If092511da36f3f493f7e3f34a35cb9eb;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[194]  <=   Ice07207e1867f71dbb58dc0b3d28f5d1;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[195]  <=   Id1c6ccb54bf2d0d03f296cbd502fac6a;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[196]  <=   I7a2b0491133ed6a2daafb889ff46d271;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[197]  <=   I4fabd40b7afb192a9c2a255512fd0852;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[198]  <=   I7b39e709a6939751b11bb3ba6fc42bde;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[199]  <=   I3a7a76b3ca144951bb6edeba1650c35a;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[200]  <=   I3c023a3a1a2ce2fb54b2292401df0019;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[201]  <=   I804cf7b8b79a124cbee51fe473e664a3;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[202]  <=   I33be2a0d4c64f50472091a4503281558;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[203]  <=   Ie5f94955ed10ae50d92d3dd0e43c8088;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[204]  <=   Ide6f35e8581e1bec17ec974448b6beed;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[205]  <=   I57b47b934005413e4c400a33e7ddc20c;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[206]  <=   Id4e7f9a0c100dfc591e7693d76a496d9;
           end
           if (Ibd047e2643dc68affb5b4f25b82ded31) begin
               tmp_bit[207]  <=   Ieda30691eb70678f7535eed71e9ee031;
           end

       end
   end

assign final_y_nr_dec = tmp_bit;


`ifdef ENCRYPT
`endif

endmodule


module Ic9c2f173881d25f8976d723957809f51 #(
`include "NR_2_0_4/fgallag/GF2_LDPC_fgallag_param_inc.sv"

) (

input wire [fgallag_SEL - 1:0]       fgallag_sel ,
output reg [fgallag_WDTH  - 1:0]     fgallag,
input wire                           start_in,
output wire                          start_out,
input wire                           rstn,
input wire                           clk

);

`include "NR_2_0_4/fgallag/GF2_LDPC_fgallag_inc_inc_all.sv"

// fgallag::'h380
`include "NR_2_0_4/fgallag/GF2_LDPC_fgallag_inc_all.sv"

assign start_d_fgallag0x00000 = start_in;
assign start_out = start_d_fgallag0xffffffff_q;

always_comb
begin
     fgallag = fgallag0xffffffff_0_q;
end


endmodule







module Ic3da32f100a43f826b89a492544e7812 #(
`include "NR_2_0_4/flogtanh/GF2_LDPC_flogtanh_param_inc.sv"

) (

input wire [flogtanh_SEL - 1:0]      flogtanh_sel ,
output reg [flogtanh_WDTH  - 1:0]    flogtanh,
input wire                           start_in,
output wire                          start_out,
input wire                           rstn,
input wire                           clk

);

`include "NR_2_0_4/flogtanh/GF2_LDPC_flogtanh_inc_inc_all.sv"

// flogtanh::'h380
`include "NR_2_0_4/flogtanh/GF2_LDPC_flogtanh_inc_all.sv"

assign start_d_flogtanh0x00000 = start_in;
assign start_out = start_d_flogtanh0xffffffff_q;

always_comb
begin
     flogtanh = flogtanh0xffffffff_0_q;
end




endmodule




//C Ia642a85aab89544a289fb1f29eab689d: Ib6f6b4efd9391d1fa207d325ff1bbd60 I83878c91171338902e0fe0fb97a8c47a:0.100000 I7290d6b1f1458098d2f225877e609ba6:2.197225 percent_probability_int:'d141

 //Ic07b0b4d7660314f711a68fc47c4ab38 I48d8d6f5a3efbf52837d6b788a22859a valid Ic13367945d5d4c91047b3b50234aa7ab Ic47d187067c6cf953245f128b5fde62a
//y_int:
 //44010bdd34c9a17a9dc5c9798ef00a0604fe89b67904e634be0b
//Iebc6097498b06421e2759a773c992ed3:
 //0200400200100008100880c0000680200320002200
//C Ia642a85aab89544a289fb1f29eab689d: Ib6f6b4efd9391d1fa207d325ff1bbd60 I83878c91171338902e0fe0fb97a8c47a:0.038462 I7290d6b1f1458098d2f225877e609ba6:3.218876 percent_probability_int:'d206
