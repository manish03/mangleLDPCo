 reg  ['h1ff:0] [$clog2('h7000+1)-1:0] I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c ;
