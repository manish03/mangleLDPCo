//`include "GF2_LDPC_fgallag_0x00010_assign_inc.sv"
//always_comb begin
              I23c1c03fb2d7ef8b2dc0921ddaf652a0['h00000] = 
          (!fgallag_sel['h00010]) ? 
                       Ice223344c1d41676e20d7b2668ccff71['h00000] : //%
                       Ice223344c1d41676e20d7b2668ccff71['h00001] ;
//end
//always_comb begin // 
               I23c1c03fb2d7ef8b2dc0921ddaf652a0['h00001] =  Ice223344c1d41676e20d7b2668ccff71['h00002] ;
//end
//always_comb begin // 
               I23c1c03fb2d7ef8b2dc0921ddaf652a0['h00002] =  Ice223344c1d41676e20d7b2668ccff71['h00004] ;
//end
//always_comb begin // 
               I23c1c03fb2d7ef8b2dc0921ddaf652a0['h00003] =  Ice223344c1d41676e20d7b2668ccff71['h00006] ;
//end
