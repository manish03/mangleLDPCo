`include "GF2_LDPC_flogtanh.sv"
`include "GF2_LDPC_flogtanh_0x00000_assign.sv"
`include "GF2_LDPC_flogtanh_0x00001_assign.sv"
`include "GF2_LDPC_flogtanh_0x00002_assign.sv"
`include "GF2_LDPC_flogtanh_0x00003_assign.sv"
`include "GF2_LDPC_flogtanh_0x00004_assign.sv"
`include "GF2_LDPC_flogtanh_0x00005_assign.sv"
`include "GF2_LDPC_flogtanh_0x00006_assign.sv"
`include "GF2_LDPC_flogtanh_0x00007_assign.sv"
`include "GF2_LDPC_flogtanh_0x00008_assign.sv"
`include "GF2_LDPC_flogtanh_0x00009_assign.sv"
`include "GF2_LDPC_flogtanh_0x0000a_assign.sv"
`include "GF2_LDPC_flogtanh_0x0000b_assign.sv"
`include "GF2_LDPC_flogtanh_0x0000c_assign.sv"
`include "GF2_LDPC_flogtanh_0x0000d_assign.sv"
`include "GF2_LDPC_flogtanh_0x0000e_assign.sv"
`include "GF2_LDPC_flogtanh_0x0000f_assign.sv"
`include "GF2_LDPC_flogtanh_0x00010_assign.sv"
`include "GF2_LDPC_flogtanh_0x00011_assign.sv"
`include "GF2_LDPC_flogtanh_0x00012_assign.sv"
