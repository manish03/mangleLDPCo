 reg  ['hffff:0] [$clog2('h7000+1)-1:0] I8b89f6bc8b4c4e5485f1e82f685bd307d9752d3cb0cc6bcc55a42210c2d367a2 ;
