//`include "GF2_LDPC_flogtanh_0x00009_assign_inc.sv"
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00000] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00000] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00001] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00001] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00002] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00003] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00002] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00004] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00005] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00003] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00006] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00007] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00004] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00008] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00009] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00005] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h0000a] : //%
                       I810764ca41a2b12d686e115c79b0578f['h0000b] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00006] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h0000c] : //%
                       I810764ca41a2b12d686e115c79b0578f['h0000d] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00007] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h0000e] : //%
                       I810764ca41a2b12d686e115c79b0578f['h0000f] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00008] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00010] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00011] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00009] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00012] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00013] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h0000a] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00014] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00015] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h0000b] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00016] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00017] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h0000c] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00018] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00019] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h0000d] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h0001a] : //%
                       I810764ca41a2b12d686e115c79b0578f['h0001b] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h0000e] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h0001c] : //%
                       I810764ca41a2b12d686e115c79b0578f['h0001d] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h0000f] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h0001e] : //%
                       I810764ca41a2b12d686e115c79b0578f['h0001f] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00010] =  I810764ca41a2b12d686e115c79b0578f['h00020] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00011] =  I810764ca41a2b12d686e115c79b0578f['h00022] ;
//end
//always_comb begin
              I986ccea2f9226242e2772b9c3af42d87['h00012] = 
          (!flogtanh_sel['h00009]) ? 
                       I810764ca41a2b12d686e115c79b0578f['h00024] : //%
                       I810764ca41a2b12d686e115c79b0578f['h00025] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00013] =  I810764ca41a2b12d686e115c79b0578f['h00026] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00014] =  I810764ca41a2b12d686e115c79b0578f['h00028] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00015] =  I810764ca41a2b12d686e115c79b0578f['h0002a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00016] =  I810764ca41a2b12d686e115c79b0578f['h0002c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00017] =  I810764ca41a2b12d686e115c79b0578f['h0002e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00018] =  I810764ca41a2b12d686e115c79b0578f['h00030] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00019] =  I810764ca41a2b12d686e115c79b0578f['h00032] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0001a] =  I810764ca41a2b12d686e115c79b0578f['h00034] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0001b] =  I810764ca41a2b12d686e115c79b0578f['h00036] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0001c] =  I810764ca41a2b12d686e115c79b0578f['h00038] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0001d] =  I810764ca41a2b12d686e115c79b0578f['h0003a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0001e] =  I810764ca41a2b12d686e115c79b0578f['h0003c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0001f] =  I810764ca41a2b12d686e115c79b0578f['h0003e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00020] =  I810764ca41a2b12d686e115c79b0578f['h00040] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00021] =  I810764ca41a2b12d686e115c79b0578f['h00042] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00022] =  I810764ca41a2b12d686e115c79b0578f['h00044] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00023] =  I810764ca41a2b12d686e115c79b0578f['h00046] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00024] =  I810764ca41a2b12d686e115c79b0578f['h00048] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00025] =  I810764ca41a2b12d686e115c79b0578f['h0004a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00026] =  I810764ca41a2b12d686e115c79b0578f['h0004c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00027] =  I810764ca41a2b12d686e115c79b0578f['h0004e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00028] =  I810764ca41a2b12d686e115c79b0578f['h00050] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00029] =  I810764ca41a2b12d686e115c79b0578f['h00052] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0002a] =  I810764ca41a2b12d686e115c79b0578f['h00054] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0002b] =  I810764ca41a2b12d686e115c79b0578f['h00056] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0002c] =  I810764ca41a2b12d686e115c79b0578f['h00058] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0002d] =  I810764ca41a2b12d686e115c79b0578f['h0005a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0002e] =  I810764ca41a2b12d686e115c79b0578f['h0005c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0002f] =  I810764ca41a2b12d686e115c79b0578f['h0005e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00030] =  I810764ca41a2b12d686e115c79b0578f['h00060] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00031] =  I810764ca41a2b12d686e115c79b0578f['h00062] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00032] =  I810764ca41a2b12d686e115c79b0578f['h00064] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00033] =  I810764ca41a2b12d686e115c79b0578f['h00066] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00034] =  I810764ca41a2b12d686e115c79b0578f['h00068] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00035] =  I810764ca41a2b12d686e115c79b0578f['h0006a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00036] =  I810764ca41a2b12d686e115c79b0578f['h0006c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00037] =  I810764ca41a2b12d686e115c79b0578f['h0006e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00038] =  I810764ca41a2b12d686e115c79b0578f['h00070] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00039] =  I810764ca41a2b12d686e115c79b0578f['h00072] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0003a] =  I810764ca41a2b12d686e115c79b0578f['h00074] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0003b] =  I810764ca41a2b12d686e115c79b0578f['h00076] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0003c] =  I810764ca41a2b12d686e115c79b0578f['h00078] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0003d] =  I810764ca41a2b12d686e115c79b0578f['h0007a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0003e] =  I810764ca41a2b12d686e115c79b0578f['h0007c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0003f] =  I810764ca41a2b12d686e115c79b0578f['h0007e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00040] =  I810764ca41a2b12d686e115c79b0578f['h00080] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00041] =  I810764ca41a2b12d686e115c79b0578f['h00082] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00042] =  I810764ca41a2b12d686e115c79b0578f['h00084] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00043] =  I810764ca41a2b12d686e115c79b0578f['h00086] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00044] =  I810764ca41a2b12d686e115c79b0578f['h00088] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00045] =  I810764ca41a2b12d686e115c79b0578f['h0008a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00046] =  I810764ca41a2b12d686e115c79b0578f['h0008c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00047] =  I810764ca41a2b12d686e115c79b0578f['h0008e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00048] =  I810764ca41a2b12d686e115c79b0578f['h00090] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00049] =  I810764ca41a2b12d686e115c79b0578f['h00092] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0004a] =  I810764ca41a2b12d686e115c79b0578f['h00094] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0004b] =  I810764ca41a2b12d686e115c79b0578f['h00096] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0004c] =  I810764ca41a2b12d686e115c79b0578f['h00098] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0004d] =  I810764ca41a2b12d686e115c79b0578f['h0009a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0004e] =  I810764ca41a2b12d686e115c79b0578f['h0009c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0004f] =  I810764ca41a2b12d686e115c79b0578f['h0009e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00050] =  I810764ca41a2b12d686e115c79b0578f['h000a0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00051] =  I810764ca41a2b12d686e115c79b0578f['h000a2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00052] =  I810764ca41a2b12d686e115c79b0578f['h000a4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00053] =  I810764ca41a2b12d686e115c79b0578f['h000a6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00054] =  I810764ca41a2b12d686e115c79b0578f['h000a8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00055] =  I810764ca41a2b12d686e115c79b0578f['h000aa] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00056] =  I810764ca41a2b12d686e115c79b0578f['h000ac] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00057] =  I810764ca41a2b12d686e115c79b0578f['h000ae] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00058] =  I810764ca41a2b12d686e115c79b0578f['h000b0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00059] =  I810764ca41a2b12d686e115c79b0578f['h000b2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0005a] =  I810764ca41a2b12d686e115c79b0578f['h000b4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0005b] =  I810764ca41a2b12d686e115c79b0578f['h000b6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0005c] =  I810764ca41a2b12d686e115c79b0578f['h000b8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0005d] =  I810764ca41a2b12d686e115c79b0578f['h000ba] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0005e] =  I810764ca41a2b12d686e115c79b0578f['h000bc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0005f] =  I810764ca41a2b12d686e115c79b0578f['h000be] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00060] =  I810764ca41a2b12d686e115c79b0578f['h000c0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00061] =  I810764ca41a2b12d686e115c79b0578f['h000c2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00062] =  I810764ca41a2b12d686e115c79b0578f['h000c4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00063] =  I810764ca41a2b12d686e115c79b0578f['h000c6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00064] =  I810764ca41a2b12d686e115c79b0578f['h000c8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00065] =  I810764ca41a2b12d686e115c79b0578f['h000ca] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00066] =  I810764ca41a2b12d686e115c79b0578f['h000cc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00067] =  I810764ca41a2b12d686e115c79b0578f['h000ce] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00068] =  I810764ca41a2b12d686e115c79b0578f['h000d0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00069] =  I810764ca41a2b12d686e115c79b0578f['h000d2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0006a] =  I810764ca41a2b12d686e115c79b0578f['h000d4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0006b] =  I810764ca41a2b12d686e115c79b0578f['h000d6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0006c] =  I810764ca41a2b12d686e115c79b0578f['h000d8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0006d] =  I810764ca41a2b12d686e115c79b0578f['h000da] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0006e] =  I810764ca41a2b12d686e115c79b0578f['h000dc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0006f] =  I810764ca41a2b12d686e115c79b0578f['h000de] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00070] =  I810764ca41a2b12d686e115c79b0578f['h000e0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00071] =  I810764ca41a2b12d686e115c79b0578f['h000e2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00072] =  I810764ca41a2b12d686e115c79b0578f['h000e4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00073] =  I810764ca41a2b12d686e115c79b0578f['h000e6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00074] =  I810764ca41a2b12d686e115c79b0578f['h000e8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00075] =  I810764ca41a2b12d686e115c79b0578f['h000ea] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00076] =  I810764ca41a2b12d686e115c79b0578f['h000ec] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00077] =  I810764ca41a2b12d686e115c79b0578f['h000ee] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00078] =  I810764ca41a2b12d686e115c79b0578f['h000f0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00079] =  I810764ca41a2b12d686e115c79b0578f['h000f2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0007a] =  I810764ca41a2b12d686e115c79b0578f['h000f4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0007b] =  I810764ca41a2b12d686e115c79b0578f['h000f6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0007c] =  I810764ca41a2b12d686e115c79b0578f['h000f8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0007d] =  I810764ca41a2b12d686e115c79b0578f['h000fa] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0007e] =  I810764ca41a2b12d686e115c79b0578f['h000fc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0007f] =  I810764ca41a2b12d686e115c79b0578f['h000fe] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00080] =  I810764ca41a2b12d686e115c79b0578f['h00100] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00081] =  I810764ca41a2b12d686e115c79b0578f['h00102] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00082] =  I810764ca41a2b12d686e115c79b0578f['h00104] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00083] =  I810764ca41a2b12d686e115c79b0578f['h00106] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00084] =  I810764ca41a2b12d686e115c79b0578f['h00108] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00085] =  I810764ca41a2b12d686e115c79b0578f['h0010a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00086] =  I810764ca41a2b12d686e115c79b0578f['h0010c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00087] =  I810764ca41a2b12d686e115c79b0578f['h0010e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00088] =  I810764ca41a2b12d686e115c79b0578f['h00110] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00089] =  I810764ca41a2b12d686e115c79b0578f['h00112] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0008a] =  I810764ca41a2b12d686e115c79b0578f['h00114] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0008b] =  I810764ca41a2b12d686e115c79b0578f['h00116] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0008c] =  I810764ca41a2b12d686e115c79b0578f['h00118] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0008d] =  I810764ca41a2b12d686e115c79b0578f['h0011a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0008e] =  I810764ca41a2b12d686e115c79b0578f['h0011c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0008f] =  I810764ca41a2b12d686e115c79b0578f['h0011e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00090] =  I810764ca41a2b12d686e115c79b0578f['h00120] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00091] =  I810764ca41a2b12d686e115c79b0578f['h00122] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00092] =  I810764ca41a2b12d686e115c79b0578f['h00124] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00093] =  I810764ca41a2b12d686e115c79b0578f['h00126] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00094] =  I810764ca41a2b12d686e115c79b0578f['h00128] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00095] =  I810764ca41a2b12d686e115c79b0578f['h0012a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00096] =  I810764ca41a2b12d686e115c79b0578f['h0012c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00097] =  I810764ca41a2b12d686e115c79b0578f['h0012e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00098] =  I810764ca41a2b12d686e115c79b0578f['h00130] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00099] =  I810764ca41a2b12d686e115c79b0578f['h00132] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0009a] =  I810764ca41a2b12d686e115c79b0578f['h00134] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0009b] =  I810764ca41a2b12d686e115c79b0578f['h00136] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0009c] =  I810764ca41a2b12d686e115c79b0578f['h00138] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0009d] =  I810764ca41a2b12d686e115c79b0578f['h0013a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0009e] =  I810764ca41a2b12d686e115c79b0578f['h0013c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0009f] =  I810764ca41a2b12d686e115c79b0578f['h0013e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a0] =  I810764ca41a2b12d686e115c79b0578f['h00140] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a1] =  I810764ca41a2b12d686e115c79b0578f['h00142] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a2] =  I810764ca41a2b12d686e115c79b0578f['h00144] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a3] =  I810764ca41a2b12d686e115c79b0578f['h00146] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a4] =  I810764ca41a2b12d686e115c79b0578f['h00148] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a5] =  I810764ca41a2b12d686e115c79b0578f['h0014a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a6] =  I810764ca41a2b12d686e115c79b0578f['h0014c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a7] =  I810764ca41a2b12d686e115c79b0578f['h0014e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a8] =  I810764ca41a2b12d686e115c79b0578f['h00150] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000a9] =  I810764ca41a2b12d686e115c79b0578f['h00152] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000aa] =  I810764ca41a2b12d686e115c79b0578f['h00154] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ab] =  I810764ca41a2b12d686e115c79b0578f['h00156] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ac] =  I810764ca41a2b12d686e115c79b0578f['h00158] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ad] =  I810764ca41a2b12d686e115c79b0578f['h0015a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ae] =  I810764ca41a2b12d686e115c79b0578f['h0015c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000af] =  I810764ca41a2b12d686e115c79b0578f['h0015e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b0] =  I810764ca41a2b12d686e115c79b0578f['h00160] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b1] =  I810764ca41a2b12d686e115c79b0578f['h00162] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b2] =  I810764ca41a2b12d686e115c79b0578f['h00164] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b3] =  I810764ca41a2b12d686e115c79b0578f['h00166] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b4] =  I810764ca41a2b12d686e115c79b0578f['h00168] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b5] =  I810764ca41a2b12d686e115c79b0578f['h0016a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b6] =  I810764ca41a2b12d686e115c79b0578f['h0016c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b7] =  I810764ca41a2b12d686e115c79b0578f['h0016e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b8] =  I810764ca41a2b12d686e115c79b0578f['h00170] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000b9] =  I810764ca41a2b12d686e115c79b0578f['h00172] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ba] =  I810764ca41a2b12d686e115c79b0578f['h00174] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000bb] =  I810764ca41a2b12d686e115c79b0578f['h00176] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000bc] =  I810764ca41a2b12d686e115c79b0578f['h00178] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000bd] =  I810764ca41a2b12d686e115c79b0578f['h0017a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000be] =  I810764ca41a2b12d686e115c79b0578f['h0017c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000bf] =  I810764ca41a2b12d686e115c79b0578f['h0017e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c0] =  I810764ca41a2b12d686e115c79b0578f['h00180] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c1] =  I810764ca41a2b12d686e115c79b0578f['h00182] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c2] =  I810764ca41a2b12d686e115c79b0578f['h00184] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c3] =  I810764ca41a2b12d686e115c79b0578f['h00186] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c4] =  I810764ca41a2b12d686e115c79b0578f['h00188] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c5] =  I810764ca41a2b12d686e115c79b0578f['h0018a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c6] =  I810764ca41a2b12d686e115c79b0578f['h0018c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c7] =  I810764ca41a2b12d686e115c79b0578f['h0018e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c8] =  I810764ca41a2b12d686e115c79b0578f['h00190] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000c9] =  I810764ca41a2b12d686e115c79b0578f['h00192] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ca] =  I810764ca41a2b12d686e115c79b0578f['h00194] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000cb] =  I810764ca41a2b12d686e115c79b0578f['h00196] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000cc] =  I810764ca41a2b12d686e115c79b0578f['h00198] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000cd] =  I810764ca41a2b12d686e115c79b0578f['h0019a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ce] =  I810764ca41a2b12d686e115c79b0578f['h0019c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000cf] =  I810764ca41a2b12d686e115c79b0578f['h0019e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d0] =  I810764ca41a2b12d686e115c79b0578f['h001a0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d1] =  I810764ca41a2b12d686e115c79b0578f['h001a2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d2] =  I810764ca41a2b12d686e115c79b0578f['h001a4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d3] =  I810764ca41a2b12d686e115c79b0578f['h001a6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d4] =  I810764ca41a2b12d686e115c79b0578f['h001a8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d5] =  I810764ca41a2b12d686e115c79b0578f['h001aa] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d6] =  I810764ca41a2b12d686e115c79b0578f['h001ac] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d7] =  I810764ca41a2b12d686e115c79b0578f['h001ae] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d8] =  I810764ca41a2b12d686e115c79b0578f['h001b0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000d9] =  I810764ca41a2b12d686e115c79b0578f['h001b2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000da] =  I810764ca41a2b12d686e115c79b0578f['h001b4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000db] =  I810764ca41a2b12d686e115c79b0578f['h001b6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000dc] =  I810764ca41a2b12d686e115c79b0578f['h001b8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000dd] =  I810764ca41a2b12d686e115c79b0578f['h001ba] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000de] =  I810764ca41a2b12d686e115c79b0578f['h001bc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000df] =  I810764ca41a2b12d686e115c79b0578f['h001be] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e0] =  I810764ca41a2b12d686e115c79b0578f['h001c0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e1] =  I810764ca41a2b12d686e115c79b0578f['h001c2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e2] =  I810764ca41a2b12d686e115c79b0578f['h001c4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e3] =  I810764ca41a2b12d686e115c79b0578f['h001c6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e4] =  I810764ca41a2b12d686e115c79b0578f['h001c8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e5] =  I810764ca41a2b12d686e115c79b0578f['h001ca] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e6] =  I810764ca41a2b12d686e115c79b0578f['h001cc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e7] =  I810764ca41a2b12d686e115c79b0578f['h001ce] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e8] =  I810764ca41a2b12d686e115c79b0578f['h001d0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000e9] =  I810764ca41a2b12d686e115c79b0578f['h001d2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ea] =  I810764ca41a2b12d686e115c79b0578f['h001d4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000eb] =  I810764ca41a2b12d686e115c79b0578f['h001d6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ec] =  I810764ca41a2b12d686e115c79b0578f['h001d8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ed] =  I810764ca41a2b12d686e115c79b0578f['h001da] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ee] =  I810764ca41a2b12d686e115c79b0578f['h001dc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ef] =  I810764ca41a2b12d686e115c79b0578f['h001de] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f0] =  I810764ca41a2b12d686e115c79b0578f['h001e0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f1] =  I810764ca41a2b12d686e115c79b0578f['h001e2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f2] =  I810764ca41a2b12d686e115c79b0578f['h001e4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f3] =  I810764ca41a2b12d686e115c79b0578f['h001e6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f4] =  I810764ca41a2b12d686e115c79b0578f['h001e8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f5] =  I810764ca41a2b12d686e115c79b0578f['h001ea] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f6] =  I810764ca41a2b12d686e115c79b0578f['h001ec] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f7] =  I810764ca41a2b12d686e115c79b0578f['h001ee] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f8] =  I810764ca41a2b12d686e115c79b0578f['h001f0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000f9] =  I810764ca41a2b12d686e115c79b0578f['h001f2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000fa] =  I810764ca41a2b12d686e115c79b0578f['h001f4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000fb] =  I810764ca41a2b12d686e115c79b0578f['h001f6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000fc] =  I810764ca41a2b12d686e115c79b0578f['h001f8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000fd] =  I810764ca41a2b12d686e115c79b0578f['h001fa] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000fe] =  I810764ca41a2b12d686e115c79b0578f['h001fc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h000ff] =  I810764ca41a2b12d686e115c79b0578f['h001fe] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00100] =  I810764ca41a2b12d686e115c79b0578f['h00200] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00101] =  I810764ca41a2b12d686e115c79b0578f['h00202] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00102] =  I810764ca41a2b12d686e115c79b0578f['h00204] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00103] =  I810764ca41a2b12d686e115c79b0578f['h00206] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00104] =  I810764ca41a2b12d686e115c79b0578f['h00208] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00105] =  I810764ca41a2b12d686e115c79b0578f['h0020a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00106] =  I810764ca41a2b12d686e115c79b0578f['h0020c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00107] =  I810764ca41a2b12d686e115c79b0578f['h0020e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00108] =  I810764ca41a2b12d686e115c79b0578f['h00210] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00109] =  I810764ca41a2b12d686e115c79b0578f['h00212] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0010a] =  I810764ca41a2b12d686e115c79b0578f['h00214] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0010b] =  I810764ca41a2b12d686e115c79b0578f['h00216] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0010c] =  I810764ca41a2b12d686e115c79b0578f['h00218] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0010d] =  I810764ca41a2b12d686e115c79b0578f['h0021a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0010e] =  I810764ca41a2b12d686e115c79b0578f['h0021c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0010f] =  I810764ca41a2b12d686e115c79b0578f['h0021e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00110] =  I810764ca41a2b12d686e115c79b0578f['h00220] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00111] =  I810764ca41a2b12d686e115c79b0578f['h00222] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00112] =  I810764ca41a2b12d686e115c79b0578f['h00224] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00113] =  I810764ca41a2b12d686e115c79b0578f['h00226] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00114] =  I810764ca41a2b12d686e115c79b0578f['h00228] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00115] =  I810764ca41a2b12d686e115c79b0578f['h0022a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00116] =  I810764ca41a2b12d686e115c79b0578f['h0022c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00117] =  I810764ca41a2b12d686e115c79b0578f['h0022e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00118] =  I810764ca41a2b12d686e115c79b0578f['h00230] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00119] =  I810764ca41a2b12d686e115c79b0578f['h00232] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0011a] =  I810764ca41a2b12d686e115c79b0578f['h00234] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0011b] =  I810764ca41a2b12d686e115c79b0578f['h00236] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0011c] =  I810764ca41a2b12d686e115c79b0578f['h00238] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0011d] =  I810764ca41a2b12d686e115c79b0578f['h0023a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0011e] =  I810764ca41a2b12d686e115c79b0578f['h0023c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0011f] =  I810764ca41a2b12d686e115c79b0578f['h0023e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00120] =  I810764ca41a2b12d686e115c79b0578f['h00240] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00121] =  I810764ca41a2b12d686e115c79b0578f['h00242] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00122] =  I810764ca41a2b12d686e115c79b0578f['h00244] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00123] =  I810764ca41a2b12d686e115c79b0578f['h00246] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00124] =  I810764ca41a2b12d686e115c79b0578f['h00248] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00125] =  I810764ca41a2b12d686e115c79b0578f['h0024a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00126] =  I810764ca41a2b12d686e115c79b0578f['h0024c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00127] =  I810764ca41a2b12d686e115c79b0578f['h0024e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00128] =  I810764ca41a2b12d686e115c79b0578f['h00250] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00129] =  I810764ca41a2b12d686e115c79b0578f['h00252] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0012a] =  I810764ca41a2b12d686e115c79b0578f['h00254] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0012b] =  I810764ca41a2b12d686e115c79b0578f['h00256] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0012c] =  I810764ca41a2b12d686e115c79b0578f['h00258] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0012d] =  I810764ca41a2b12d686e115c79b0578f['h0025a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0012e] =  I810764ca41a2b12d686e115c79b0578f['h0025c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0012f] =  I810764ca41a2b12d686e115c79b0578f['h0025e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00130] =  I810764ca41a2b12d686e115c79b0578f['h00260] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00131] =  I810764ca41a2b12d686e115c79b0578f['h00262] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00132] =  I810764ca41a2b12d686e115c79b0578f['h00264] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00133] =  I810764ca41a2b12d686e115c79b0578f['h00266] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00134] =  I810764ca41a2b12d686e115c79b0578f['h00268] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00135] =  I810764ca41a2b12d686e115c79b0578f['h0026a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00136] =  I810764ca41a2b12d686e115c79b0578f['h0026c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00137] =  I810764ca41a2b12d686e115c79b0578f['h0026e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00138] =  I810764ca41a2b12d686e115c79b0578f['h00270] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00139] =  I810764ca41a2b12d686e115c79b0578f['h00272] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0013a] =  I810764ca41a2b12d686e115c79b0578f['h00274] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0013b] =  I810764ca41a2b12d686e115c79b0578f['h00276] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0013c] =  I810764ca41a2b12d686e115c79b0578f['h00278] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0013d] =  I810764ca41a2b12d686e115c79b0578f['h0027a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0013e] =  I810764ca41a2b12d686e115c79b0578f['h0027c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0013f] =  I810764ca41a2b12d686e115c79b0578f['h0027e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00140] =  I810764ca41a2b12d686e115c79b0578f['h00280] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00141] =  I810764ca41a2b12d686e115c79b0578f['h00282] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00142] =  I810764ca41a2b12d686e115c79b0578f['h00284] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00143] =  I810764ca41a2b12d686e115c79b0578f['h00286] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00144] =  I810764ca41a2b12d686e115c79b0578f['h00288] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00145] =  I810764ca41a2b12d686e115c79b0578f['h0028a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00146] =  I810764ca41a2b12d686e115c79b0578f['h0028c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00147] =  I810764ca41a2b12d686e115c79b0578f['h0028e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00148] =  I810764ca41a2b12d686e115c79b0578f['h00290] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00149] =  I810764ca41a2b12d686e115c79b0578f['h00292] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0014a] =  I810764ca41a2b12d686e115c79b0578f['h00294] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0014b] =  I810764ca41a2b12d686e115c79b0578f['h00296] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0014c] =  I810764ca41a2b12d686e115c79b0578f['h00298] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0014d] =  I810764ca41a2b12d686e115c79b0578f['h0029a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0014e] =  I810764ca41a2b12d686e115c79b0578f['h0029c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0014f] =  I810764ca41a2b12d686e115c79b0578f['h0029e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00150] =  I810764ca41a2b12d686e115c79b0578f['h002a0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00151] =  I810764ca41a2b12d686e115c79b0578f['h002a2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00152] =  I810764ca41a2b12d686e115c79b0578f['h002a4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00153] =  I810764ca41a2b12d686e115c79b0578f['h002a6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00154] =  I810764ca41a2b12d686e115c79b0578f['h002a8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00155] =  I810764ca41a2b12d686e115c79b0578f['h002aa] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00156] =  I810764ca41a2b12d686e115c79b0578f['h002ac] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00157] =  I810764ca41a2b12d686e115c79b0578f['h002ae] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00158] =  I810764ca41a2b12d686e115c79b0578f['h002b0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00159] =  I810764ca41a2b12d686e115c79b0578f['h002b2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0015a] =  I810764ca41a2b12d686e115c79b0578f['h002b4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0015b] =  I810764ca41a2b12d686e115c79b0578f['h002b6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0015c] =  I810764ca41a2b12d686e115c79b0578f['h002b8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0015d] =  I810764ca41a2b12d686e115c79b0578f['h002ba] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0015e] =  I810764ca41a2b12d686e115c79b0578f['h002bc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0015f] =  I810764ca41a2b12d686e115c79b0578f['h002be] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00160] =  I810764ca41a2b12d686e115c79b0578f['h002c0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00161] =  I810764ca41a2b12d686e115c79b0578f['h002c2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00162] =  I810764ca41a2b12d686e115c79b0578f['h002c4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00163] =  I810764ca41a2b12d686e115c79b0578f['h002c6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00164] =  I810764ca41a2b12d686e115c79b0578f['h002c8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00165] =  I810764ca41a2b12d686e115c79b0578f['h002ca] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00166] =  I810764ca41a2b12d686e115c79b0578f['h002cc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00167] =  I810764ca41a2b12d686e115c79b0578f['h002ce] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00168] =  I810764ca41a2b12d686e115c79b0578f['h002d0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00169] =  I810764ca41a2b12d686e115c79b0578f['h002d2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0016a] =  I810764ca41a2b12d686e115c79b0578f['h002d4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0016b] =  I810764ca41a2b12d686e115c79b0578f['h002d6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0016c] =  I810764ca41a2b12d686e115c79b0578f['h002d8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0016d] =  I810764ca41a2b12d686e115c79b0578f['h002da] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0016e] =  I810764ca41a2b12d686e115c79b0578f['h002dc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0016f] =  I810764ca41a2b12d686e115c79b0578f['h002de] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00170] =  I810764ca41a2b12d686e115c79b0578f['h002e0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00171] =  I810764ca41a2b12d686e115c79b0578f['h002e2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00172] =  I810764ca41a2b12d686e115c79b0578f['h002e4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00173] =  I810764ca41a2b12d686e115c79b0578f['h002e6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00174] =  I810764ca41a2b12d686e115c79b0578f['h002e8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00175] =  I810764ca41a2b12d686e115c79b0578f['h002ea] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00176] =  I810764ca41a2b12d686e115c79b0578f['h002ec] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00177] =  I810764ca41a2b12d686e115c79b0578f['h002ee] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00178] =  I810764ca41a2b12d686e115c79b0578f['h002f0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00179] =  I810764ca41a2b12d686e115c79b0578f['h002f2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0017a] =  I810764ca41a2b12d686e115c79b0578f['h002f4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0017b] =  I810764ca41a2b12d686e115c79b0578f['h002f6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0017c] =  I810764ca41a2b12d686e115c79b0578f['h002f8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0017d] =  I810764ca41a2b12d686e115c79b0578f['h002fa] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0017e] =  I810764ca41a2b12d686e115c79b0578f['h002fc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0017f] =  I810764ca41a2b12d686e115c79b0578f['h002fe] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00180] =  I810764ca41a2b12d686e115c79b0578f['h00300] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00181] =  I810764ca41a2b12d686e115c79b0578f['h00302] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00182] =  I810764ca41a2b12d686e115c79b0578f['h00304] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00183] =  I810764ca41a2b12d686e115c79b0578f['h00306] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00184] =  I810764ca41a2b12d686e115c79b0578f['h00308] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00185] =  I810764ca41a2b12d686e115c79b0578f['h0030a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00186] =  I810764ca41a2b12d686e115c79b0578f['h0030c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00187] =  I810764ca41a2b12d686e115c79b0578f['h0030e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00188] =  I810764ca41a2b12d686e115c79b0578f['h00310] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00189] =  I810764ca41a2b12d686e115c79b0578f['h00312] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0018a] =  I810764ca41a2b12d686e115c79b0578f['h00314] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0018b] =  I810764ca41a2b12d686e115c79b0578f['h00316] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0018c] =  I810764ca41a2b12d686e115c79b0578f['h00318] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0018d] =  I810764ca41a2b12d686e115c79b0578f['h0031a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0018e] =  I810764ca41a2b12d686e115c79b0578f['h0031c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0018f] =  I810764ca41a2b12d686e115c79b0578f['h0031e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00190] =  I810764ca41a2b12d686e115c79b0578f['h00320] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00191] =  I810764ca41a2b12d686e115c79b0578f['h00322] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00192] =  I810764ca41a2b12d686e115c79b0578f['h00324] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00193] =  I810764ca41a2b12d686e115c79b0578f['h00326] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00194] =  I810764ca41a2b12d686e115c79b0578f['h00328] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00195] =  I810764ca41a2b12d686e115c79b0578f['h0032a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00196] =  I810764ca41a2b12d686e115c79b0578f['h0032c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00197] =  I810764ca41a2b12d686e115c79b0578f['h0032e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00198] =  I810764ca41a2b12d686e115c79b0578f['h00330] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h00199] =  I810764ca41a2b12d686e115c79b0578f['h00332] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0019a] =  I810764ca41a2b12d686e115c79b0578f['h00334] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0019b] =  I810764ca41a2b12d686e115c79b0578f['h00336] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0019c] =  I810764ca41a2b12d686e115c79b0578f['h00338] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0019d] =  I810764ca41a2b12d686e115c79b0578f['h0033a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0019e] =  I810764ca41a2b12d686e115c79b0578f['h0033c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h0019f] =  I810764ca41a2b12d686e115c79b0578f['h0033e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a0] =  I810764ca41a2b12d686e115c79b0578f['h00340] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a1] =  I810764ca41a2b12d686e115c79b0578f['h00342] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a2] =  I810764ca41a2b12d686e115c79b0578f['h00344] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a3] =  I810764ca41a2b12d686e115c79b0578f['h00346] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a4] =  I810764ca41a2b12d686e115c79b0578f['h00348] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a5] =  I810764ca41a2b12d686e115c79b0578f['h0034a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a6] =  I810764ca41a2b12d686e115c79b0578f['h0034c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a7] =  I810764ca41a2b12d686e115c79b0578f['h0034e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a8] =  I810764ca41a2b12d686e115c79b0578f['h00350] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001a9] =  I810764ca41a2b12d686e115c79b0578f['h00352] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001aa] =  I810764ca41a2b12d686e115c79b0578f['h00354] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ab] =  I810764ca41a2b12d686e115c79b0578f['h00356] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ac] =  I810764ca41a2b12d686e115c79b0578f['h00358] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ad] =  I810764ca41a2b12d686e115c79b0578f['h0035a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ae] =  I810764ca41a2b12d686e115c79b0578f['h0035c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001af] =  I810764ca41a2b12d686e115c79b0578f['h0035e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b0] =  I810764ca41a2b12d686e115c79b0578f['h00360] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b1] =  I810764ca41a2b12d686e115c79b0578f['h00362] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b2] =  I810764ca41a2b12d686e115c79b0578f['h00364] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b3] =  I810764ca41a2b12d686e115c79b0578f['h00366] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b4] =  I810764ca41a2b12d686e115c79b0578f['h00368] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b5] =  I810764ca41a2b12d686e115c79b0578f['h0036a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b6] =  I810764ca41a2b12d686e115c79b0578f['h0036c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b7] =  I810764ca41a2b12d686e115c79b0578f['h0036e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b8] =  I810764ca41a2b12d686e115c79b0578f['h00370] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001b9] =  I810764ca41a2b12d686e115c79b0578f['h00372] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ba] =  I810764ca41a2b12d686e115c79b0578f['h00374] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001bb] =  I810764ca41a2b12d686e115c79b0578f['h00376] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001bc] =  I810764ca41a2b12d686e115c79b0578f['h00378] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001bd] =  I810764ca41a2b12d686e115c79b0578f['h0037a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001be] =  I810764ca41a2b12d686e115c79b0578f['h0037c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001bf] =  I810764ca41a2b12d686e115c79b0578f['h0037e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c0] =  I810764ca41a2b12d686e115c79b0578f['h00380] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c1] =  I810764ca41a2b12d686e115c79b0578f['h00382] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c2] =  I810764ca41a2b12d686e115c79b0578f['h00384] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c3] =  I810764ca41a2b12d686e115c79b0578f['h00386] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c4] =  I810764ca41a2b12d686e115c79b0578f['h00388] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c5] =  I810764ca41a2b12d686e115c79b0578f['h0038a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c6] =  I810764ca41a2b12d686e115c79b0578f['h0038c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c7] =  I810764ca41a2b12d686e115c79b0578f['h0038e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c8] =  I810764ca41a2b12d686e115c79b0578f['h00390] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001c9] =  I810764ca41a2b12d686e115c79b0578f['h00392] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ca] =  I810764ca41a2b12d686e115c79b0578f['h00394] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001cb] =  I810764ca41a2b12d686e115c79b0578f['h00396] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001cc] =  I810764ca41a2b12d686e115c79b0578f['h00398] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001cd] =  I810764ca41a2b12d686e115c79b0578f['h0039a] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ce] =  I810764ca41a2b12d686e115c79b0578f['h0039c] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001cf] =  I810764ca41a2b12d686e115c79b0578f['h0039e] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d0] =  I810764ca41a2b12d686e115c79b0578f['h003a0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d1] =  I810764ca41a2b12d686e115c79b0578f['h003a2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d2] =  I810764ca41a2b12d686e115c79b0578f['h003a4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d3] =  I810764ca41a2b12d686e115c79b0578f['h003a6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d4] =  I810764ca41a2b12d686e115c79b0578f['h003a8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d5] =  I810764ca41a2b12d686e115c79b0578f['h003aa] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d6] =  I810764ca41a2b12d686e115c79b0578f['h003ac] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d7] =  I810764ca41a2b12d686e115c79b0578f['h003ae] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d8] =  I810764ca41a2b12d686e115c79b0578f['h003b0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001d9] =  I810764ca41a2b12d686e115c79b0578f['h003b2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001da] =  I810764ca41a2b12d686e115c79b0578f['h003b4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001db] =  I810764ca41a2b12d686e115c79b0578f['h003b6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001dc] =  I810764ca41a2b12d686e115c79b0578f['h003b8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001dd] =  I810764ca41a2b12d686e115c79b0578f['h003ba] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001de] =  I810764ca41a2b12d686e115c79b0578f['h003bc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001df] =  I810764ca41a2b12d686e115c79b0578f['h003be] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e0] =  I810764ca41a2b12d686e115c79b0578f['h003c0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e1] =  I810764ca41a2b12d686e115c79b0578f['h003c2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e2] =  I810764ca41a2b12d686e115c79b0578f['h003c4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e3] =  I810764ca41a2b12d686e115c79b0578f['h003c6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e4] =  I810764ca41a2b12d686e115c79b0578f['h003c8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e5] =  I810764ca41a2b12d686e115c79b0578f['h003ca] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e6] =  I810764ca41a2b12d686e115c79b0578f['h003cc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e7] =  I810764ca41a2b12d686e115c79b0578f['h003ce] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e8] =  I810764ca41a2b12d686e115c79b0578f['h003d0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001e9] =  I810764ca41a2b12d686e115c79b0578f['h003d2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ea] =  I810764ca41a2b12d686e115c79b0578f['h003d4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001eb] =  I810764ca41a2b12d686e115c79b0578f['h003d6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ec] =  I810764ca41a2b12d686e115c79b0578f['h003d8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ed] =  I810764ca41a2b12d686e115c79b0578f['h003da] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ee] =  I810764ca41a2b12d686e115c79b0578f['h003dc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ef] =  I810764ca41a2b12d686e115c79b0578f['h003de] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f0] =  I810764ca41a2b12d686e115c79b0578f['h003e0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f1] =  I810764ca41a2b12d686e115c79b0578f['h003e2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f2] =  I810764ca41a2b12d686e115c79b0578f['h003e4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f3] =  I810764ca41a2b12d686e115c79b0578f['h003e6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f4] =  I810764ca41a2b12d686e115c79b0578f['h003e8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f5] =  I810764ca41a2b12d686e115c79b0578f['h003ea] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f6] =  I810764ca41a2b12d686e115c79b0578f['h003ec] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f7] =  I810764ca41a2b12d686e115c79b0578f['h003ee] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f8] =  I810764ca41a2b12d686e115c79b0578f['h003f0] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001f9] =  I810764ca41a2b12d686e115c79b0578f['h003f2] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001fa] =  I810764ca41a2b12d686e115c79b0578f['h003f4] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001fb] =  I810764ca41a2b12d686e115c79b0578f['h003f6] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001fc] =  I810764ca41a2b12d686e115c79b0578f['h003f8] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001fd] =  I810764ca41a2b12d686e115c79b0578f['h003fa] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001fe] =  I810764ca41a2b12d686e115c79b0578f['h003fc] ;
//end
//always_comb begin // 
               I986ccea2f9226242e2772b9c3af42d87['h001ff] =  I810764ca41a2b12d686e115c79b0578f['h003fe] ;
//end
