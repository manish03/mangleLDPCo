//`include "GF2_LDPC_flogtanh_0x0000a_assign_inc.sv"
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00000] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00000] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00001] ;
//end
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00001] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00002] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00003] ;
//end
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00002] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00004] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00005] ;
//end
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00003] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00006] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00007] ;
//end
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00004] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00008] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00009] ;
//end
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00005] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000a] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000b] ;
//end
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00006] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000c] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000d] ;
//end
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00007] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000e] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0000f] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00008] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00010] ;
//end
//always_comb begin
              I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00009] = 
          (!flogtanh_sel['h0000a]) ? 
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00012] : //%
                       I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00013] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00014] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00016] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00018] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0000f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0001e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00010] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00020] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00011] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00022] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00012] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00024] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00013] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00026] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00014] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00028] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00015] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00016] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00017] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0002e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00018] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00030] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00019] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00032] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00034] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00036] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00038] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0001f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0003e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00020] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00040] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00021] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00042] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00022] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00044] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00023] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00046] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00024] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00048] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00025] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00026] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00027] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0004e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00028] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00050] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00029] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00052] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00054] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00056] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00058] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0002f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0005e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00030] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00060] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00031] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00062] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00032] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00064] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00033] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00066] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00034] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00068] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00035] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00036] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00037] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0006e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00038] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00070] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00039] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00072] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00074] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00076] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00078] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0003f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0007e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00040] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00080] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00041] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00082] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00042] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00084] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00043] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00086] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00044] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00088] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00045] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00046] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00047] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0008e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00048] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00090] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00049] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00092] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00094] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00096] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00098] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0004f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0009e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00050] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00051] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00052] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00053] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00054] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000a8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00055] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000aa] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00056] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ac] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00057] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ae] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00058] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00059] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000b8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ba] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000bc] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0005f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000be] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00060] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00061] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00062] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00063] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00064] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000c8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00065] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ca] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00066] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000cc] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00067] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ce] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00068] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00069] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000d8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000da] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000dc] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0006f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000de] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00070] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00071] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00072] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00073] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00074] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000e8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00075] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ea] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00076] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ec] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00077] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000ee] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00078] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00079] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000f8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000fa] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000fc] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0007f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h000fe] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00080] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00100] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00081] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00102] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00082] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00104] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00083] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00106] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00084] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00108] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00085] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00086] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00087] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0010e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00088] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00110] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00089] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00112] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00114] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00116] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00118] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0008f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0011e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00090] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00120] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00091] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00122] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00092] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00124] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00093] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00126] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00094] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00128] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00095] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00096] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00097] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0012e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00098] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00130] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h00099] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00132] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009a] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00134] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009b] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00136] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009c] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00138] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009d] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009e] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h0009f] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0013e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a0] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00140] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a1] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00142] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a2] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00144] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a3] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00146] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a4] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00148] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a5] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a6] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a7] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0014e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a8] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00150] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000a9] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00152] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000aa] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00154] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ab] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00156] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ac] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00158] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ad] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ae] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000af] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0015e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b0] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00160] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b1] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00162] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b2] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00164] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b3] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00166] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b4] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00168] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b5] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b6] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b7] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0016e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b8] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00170] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000b9] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00172] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ba] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00174] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000bb] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00176] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000bc] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00178] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000bd] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000be] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000bf] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0017e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c0] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00180] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c1] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00182] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c2] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00184] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c3] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00186] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c4] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00188] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c5] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c6] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c7] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0018e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c8] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00190] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000c9] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00192] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ca] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00194] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000cb] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00196] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000cc] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h00198] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000cd] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019a] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ce] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019c] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000cf] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h0019e] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d0] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d1] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d2] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d3] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d4] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001a8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d5] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001aa] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d6] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ac] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d7] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ae] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d8] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000d9] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000da] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000db] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000dc] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001b8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000dd] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ba] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000de] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001bc] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000df] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001be] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e0] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e1] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e2] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e3] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e4] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001c8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e5] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ca] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e6] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001cc] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e7] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ce] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e8] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000e9] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ea] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000eb] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ec] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001d8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ed] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001da] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ee] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001dc] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ef] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001de] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f0] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f1] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f2] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f3] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f4] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001e8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f5] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ea] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f6] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ec] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f7] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001ee] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f8] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f0] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000f9] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f2] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000fa] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f4] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000fb] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f6] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000fc] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001f8] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000fd] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001fa] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000fe] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001fc] ;
//end
//always_comb begin // 
               I2ecbcc572903aaa9f9e6bfb59957cff826adf9fe96957361e1672bd8af0514dd['h000ff] =  I788dad44cd5e5d97be2f1de201a0d998975cc499b5a5f05f0dc940adc7d56d6c['h001fe] ;
//end
