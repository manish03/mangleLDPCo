reg [fgallag_WDTH -1:0] fgallag0x00000_0,  fgallag0x00000_0_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_1,  fgallag0x00000_1_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_2,  fgallag0x00000_2_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_3,  fgallag0x00000_3_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_4,  fgallag0x00000_4_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_5,  fgallag0x00000_5_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_6,  fgallag0x00000_6_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_7,  fgallag0x00000_7_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_8,  fgallag0x00000_8_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_9,  fgallag0x00000_9_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_10,  fgallag0x00000_10_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_11,  fgallag0x00000_11_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_12,  fgallag0x00000_12_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_13,  fgallag0x00000_13_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_14,  fgallag0x00000_14_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_15,  fgallag0x00000_15_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_16,  fgallag0x00000_16_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_17,  fgallag0x00000_17_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_18,  fgallag0x00000_18_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_19,  fgallag0x00000_19_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_20,  fgallag0x00000_20_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_21,  fgallag0x00000_21_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_22,  fgallag0x00000_22_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_23,  fgallag0x00000_23_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_24,  fgallag0x00000_24_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_25,  fgallag0x00000_25_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_26,  fgallag0x00000_26_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_27,  fgallag0x00000_27_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_28,  fgallag0x00000_28_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_29,  fgallag0x00000_29_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_30,  fgallag0x00000_30_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_31,  fgallag0x00000_31_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_32,  fgallag0x00000_32_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_33,  fgallag0x00000_33_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_34,  fgallag0x00000_34_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_35,  fgallag0x00000_35_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_36,  fgallag0x00000_36_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_37,  fgallag0x00000_37_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_38,  fgallag0x00000_38_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_39,  fgallag0x00000_39_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_40,  fgallag0x00000_40_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_41,  fgallag0x00000_41_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_42,  fgallag0x00000_42_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_43,  fgallag0x00000_43_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_44,  fgallag0x00000_44_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_45,  fgallag0x00000_45_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_46,  fgallag0x00000_46_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_47,  fgallag0x00000_47_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_48,  fgallag0x00000_48_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_49,  fgallag0x00000_49_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_50,  fgallag0x00000_50_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_51,  fgallag0x00000_51_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_52,  fgallag0x00000_52_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_53,  fgallag0x00000_53_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_54,  fgallag0x00000_54_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_55,  fgallag0x00000_55_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_56,  fgallag0x00000_56_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_57,  fgallag0x00000_57_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_58,  fgallag0x00000_58_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_59,  fgallag0x00000_59_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_60,  fgallag0x00000_60_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_61,  fgallag0x00000_61_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_62,  fgallag0x00000_62_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_63,  fgallag0x00000_63_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_64,  fgallag0x00000_64_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_65,  fgallag0x00000_65_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_66,  fgallag0x00000_66_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_67,  fgallag0x00000_67_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_68,  fgallag0x00000_68_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_69,  fgallag0x00000_69_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_70,  fgallag0x00000_70_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_71,  fgallag0x00000_71_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_72,  fgallag0x00000_72_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_73,  fgallag0x00000_73_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_74,  fgallag0x00000_74_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_75,  fgallag0x00000_75_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_76,  fgallag0x00000_76_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_77,  fgallag0x00000_77_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_78,  fgallag0x00000_78_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_79,  fgallag0x00000_79_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_80,  fgallag0x00000_80_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_81,  fgallag0x00000_81_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_82,  fgallag0x00000_82_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_83,  fgallag0x00000_83_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_84,  fgallag0x00000_84_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_85,  fgallag0x00000_85_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_86,  fgallag0x00000_86_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_87,  fgallag0x00000_87_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_88,  fgallag0x00000_88_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_89,  fgallag0x00000_89_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_90,  fgallag0x00000_90_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_91,  fgallag0x00000_91_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_92,  fgallag0x00000_92_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_93,  fgallag0x00000_93_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_94,  fgallag0x00000_94_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_95,  fgallag0x00000_95_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_96,  fgallag0x00000_96_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_97,  fgallag0x00000_97_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_98,  fgallag0x00000_98_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_99,  fgallag0x00000_99_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_100,  fgallag0x00000_100_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_101,  fgallag0x00000_101_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_102,  fgallag0x00000_102_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_103,  fgallag0x00000_103_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_104,  fgallag0x00000_104_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_105,  fgallag0x00000_105_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_106,  fgallag0x00000_106_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_107,  fgallag0x00000_107_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_108,  fgallag0x00000_108_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_109,  fgallag0x00000_109_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_110,  fgallag0x00000_110_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_111,  fgallag0x00000_111_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_112,  fgallag0x00000_112_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_113,  fgallag0x00000_113_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_114,  fgallag0x00000_114_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_115,  fgallag0x00000_115_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_116,  fgallag0x00000_116_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_117,  fgallag0x00000_117_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_118,  fgallag0x00000_118_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_119,  fgallag0x00000_119_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_120,  fgallag0x00000_120_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_121,  fgallag0x00000_121_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_122,  fgallag0x00000_122_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_123,  fgallag0x00000_123_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_124,  fgallag0x00000_124_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_125,  fgallag0x00000_125_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_126,  fgallag0x00000_126_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_127,  fgallag0x00000_127_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_128,  fgallag0x00000_128_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_129,  fgallag0x00000_129_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_130,  fgallag0x00000_130_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_131,  fgallag0x00000_131_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_132,  fgallag0x00000_132_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_133,  fgallag0x00000_133_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_134,  fgallag0x00000_134_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_135,  fgallag0x00000_135_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_136,  fgallag0x00000_136_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_137,  fgallag0x00000_137_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_138,  fgallag0x00000_138_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_139,  fgallag0x00000_139_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_140,  fgallag0x00000_140_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_141,  fgallag0x00000_141_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_142,  fgallag0x00000_142_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_143,  fgallag0x00000_143_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_144,  fgallag0x00000_144_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_145,  fgallag0x00000_145_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_146,  fgallag0x00000_146_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_147,  fgallag0x00000_147_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_148,  fgallag0x00000_148_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_149,  fgallag0x00000_149_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_150,  fgallag0x00000_150_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_151,  fgallag0x00000_151_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_152,  fgallag0x00000_152_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_153,  fgallag0x00000_153_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_154,  fgallag0x00000_154_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_155,  fgallag0x00000_155_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_156,  fgallag0x00000_156_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_157,  fgallag0x00000_157_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_158,  fgallag0x00000_158_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_159,  fgallag0x00000_159_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_160,  fgallag0x00000_160_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_161,  fgallag0x00000_161_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_162,  fgallag0x00000_162_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_163,  fgallag0x00000_163_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_164,  fgallag0x00000_164_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_165,  fgallag0x00000_165_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_166,  fgallag0x00000_166_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_167,  fgallag0x00000_167_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_168,  fgallag0x00000_168_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_169,  fgallag0x00000_169_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_170,  fgallag0x00000_170_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_171,  fgallag0x00000_171_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_172,  fgallag0x00000_172_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_173,  fgallag0x00000_173_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_174,  fgallag0x00000_174_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_175,  fgallag0x00000_175_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_176,  fgallag0x00000_176_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_177,  fgallag0x00000_177_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_178,  fgallag0x00000_178_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_179,  fgallag0x00000_179_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_180,  fgallag0x00000_180_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_181,  fgallag0x00000_181_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_182,  fgallag0x00000_182_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_183,  fgallag0x00000_183_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_184,  fgallag0x00000_184_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_185,  fgallag0x00000_185_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_186,  fgallag0x00000_186_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_187,  fgallag0x00000_187_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_188,  fgallag0x00000_188_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_189,  fgallag0x00000_189_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_190,  fgallag0x00000_190_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_191,  fgallag0x00000_191_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_192,  fgallag0x00000_192_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_193,  fgallag0x00000_193_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_194,  fgallag0x00000_194_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_195,  fgallag0x00000_195_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_196,  fgallag0x00000_196_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_197,  fgallag0x00000_197_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_198,  fgallag0x00000_198_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_199,  fgallag0x00000_199_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_200,  fgallag0x00000_200_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_201,  fgallag0x00000_201_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_202,  fgallag0x00000_202_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_203,  fgallag0x00000_203_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_204,  fgallag0x00000_204_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_205,  fgallag0x00000_205_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_206,  fgallag0x00000_206_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_207,  fgallag0x00000_207_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_208,  fgallag0x00000_208_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_209,  fgallag0x00000_209_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_210,  fgallag0x00000_210_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_211,  fgallag0x00000_211_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_212,  fgallag0x00000_212_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_213,  fgallag0x00000_213_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_214,  fgallag0x00000_214_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_215,  fgallag0x00000_215_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_216,  fgallag0x00000_216_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_217,  fgallag0x00000_217_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_218,  fgallag0x00000_218_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_219,  fgallag0x00000_219_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_220,  fgallag0x00000_220_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_221,  fgallag0x00000_221_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_222,  fgallag0x00000_222_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_223,  fgallag0x00000_223_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_224,  fgallag0x00000_224_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_225,  fgallag0x00000_225_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_226,  fgallag0x00000_226_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_227,  fgallag0x00000_227_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_228,  fgallag0x00000_228_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_229,  fgallag0x00000_229_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_230,  fgallag0x00000_230_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_231,  fgallag0x00000_231_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_232,  fgallag0x00000_232_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_233,  fgallag0x00000_233_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_234,  fgallag0x00000_234_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_235,  fgallag0x00000_235_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_236,  fgallag0x00000_236_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_237,  fgallag0x00000_237_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_238,  fgallag0x00000_238_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_239,  fgallag0x00000_239_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_240,  fgallag0x00000_240_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_241,  fgallag0x00000_241_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_242,  fgallag0x00000_242_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_243,  fgallag0x00000_243_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_244,  fgallag0x00000_244_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_245,  fgallag0x00000_245_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_246,  fgallag0x00000_246_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_247,  fgallag0x00000_247_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_248,  fgallag0x00000_248_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_249,  fgallag0x00000_249_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_250,  fgallag0x00000_250_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_251,  fgallag0x00000_251_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_252,  fgallag0x00000_252_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_253,  fgallag0x00000_253_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_254,  fgallag0x00000_254_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_255,  fgallag0x00000_255_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_256,  fgallag0x00000_256_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_257,  fgallag0x00000_257_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_258,  fgallag0x00000_258_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_259,  fgallag0x00000_259_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_260,  fgallag0x00000_260_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_261,  fgallag0x00000_261_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_262,  fgallag0x00000_262_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_263,  fgallag0x00000_263_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_264,  fgallag0x00000_264_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_265,  fgallag0x00000_265_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_266,  fgallag0x00000_266_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_267,  fgallag0x00000_267_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_268,  fgallag0x00000_268_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_269,  fgallag0x00000_269_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_270,  fgallag0x00000_270_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_271,  fgallag0x00000_271_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_272,  fgallag0x00000_272_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_273,  fgallag0x00000_273_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_274,  fgallag0x00000_274_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_275,  fgallag0x00000_275_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_276,  fgallag0x00000_276_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_277,  fgallag0x00000_277_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_278,  fgallag0x00000_278_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_279,  fgallag0x00000_279_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_280,  fgallag0x00000_280_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_281,  fgallag0x00000_281_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_282,  fgallag0x00000_282_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_283,  fgallag0x00000_283_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_284,  fgallag0x00000_284_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_285,  fgallag0x00000_285_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_286,  fgallag0x00000_286_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_287,  fgallag0x00000_287_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_288,  fgallag0x00000_288_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_289,  fgallag0x00000_289_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_290,  fgallag0x00000_290_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_291,  fgallag0x00000_291_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_292,  fgallag0x00000_292_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_293,  fgallag0x00000_293_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_294,  fgallag0x00000_294_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_295,  fgallag0x00000_295_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_296,  fgallag0x00000_296_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_297,  fgallag0x00000_297_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_298,  fgallag0x00000_298_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_299,  fgallag0x00000_299_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_300,  fgallag0x00000_300_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_301,  fgallag0x00000_301_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_302,  fgallag0x00000_302_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_303,  fgallag0x00000_303_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_304,  fgallag0x00000_304_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_305,  fgallag0x00000_305_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_306,  fgallag0x00000_306_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_307,  fgallag0x00000_307_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_308,  fgallag0x00000_308_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_309,  fgallag0x00000_309_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_310,  fgallag0x00000_310_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_311,  fgallag0x00000_311_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_312,  fgallag0x00000_312_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_313,  fgallag0x00000_313_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_314,  fgallag0x00000_314_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_315,  fgallag0x00000_315_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_316,  fgallag0x00000_316_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_317,  fgallag0x00000_317_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_318,  fgallag0x00000_318_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_319,  fgallag0x00000_319_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_320,  fgallag0x00000_320_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_321,  fgallag0x00000_321_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_322,  fgallag0x00000_322_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_323,  fgallag0x00000_323_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_324,  fgallag0x00000_324_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_325,  fgallag0x00000_325_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_326,  fgallag0x00000_326_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_327,  fgallag0x00000_327_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_328,  fgallag0x00000_328_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_329,  fgallag0x00000_329_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_330,  fgallag0x00000_330_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_331,  fgallag0x00000_331_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_332,  fgallag0x00000_332_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_333,  fgallag0x00000_333_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_334,  fgallag0x00000_334_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_335,  fgallag0x00000_335_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_336,  fgallag0x00000_336_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_337,  fgallag0x00000_337_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_338,  fgallag0x00000_338_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_339,  fgallag0x00000_339_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_340,  fgallag0x00000_340_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_341,  fgallag0x00000_341_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_342,  fgallag0x00000_342_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_343,  fgallag0x00000_343_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_344,  fgallag0x00000_344_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_345,  fgallag0x00000_345_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_346,  fgallag0x00000_346_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_347,  fgallag0x00000_347_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_348,  fgallag0x00000_348_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_349,  fgallag0x00000_349_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_350,  fgallag0x00000_350_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_351,  fgallag0x00000_351_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_352,  fgallag0x00000_352_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_353,  fgallag0x00000_353_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_354,  fgallag0x00000_354_q;
reg [fgallag_WDTH -1:0] fgallag0x00000_355,  fgallag0x00000_355_q;
wire start_d_fgallag0x00000;
reg start_d_fgallag0x00000_q;
always @(posedge clk or negedge rstn)
if (!rstn) begin
 fgallag0x00000_0_q <= 'h0;
 fgallag0x00000_1_q <= 'h0;
 fgallag0x00000_2_q <= 'h0;
 fgallag0x00000_3_q <= 'h0;
 fgallag0x00000_4_q <= 'h0;
 fgallag0x00000_5_q <= 'h0;
 fgallag0x00000_6_q <= 'h0;
 fgallag0x00000_7_q <= 'h0;
 fgallag0x00000_8_q <= 'h0;
 fgallag0x00000_9_q <= 'h0;
 fgallag0x00000_10_q <= 'h0;
 fgallag0x00000_11_q <= 'h0;
 fgallag0x00000_12_q <= 'h0;
 fgallag0x00000_13_q <= 'h0;
 fgallag0x00000_14_q <= 'h0;
 fgallag0x00000_15_q <= 'h0;
 fgallag0x00000_16_q <= 'h0;
 fgallag0x00000_17_q <= 'h0;
 fgallag0x00000_18_q <= 'h0;
 fgallag0x00000_19_q <= 'h0;
 fgallag0x00000_20_q <= 'h0;
 fgallag0x00000_21_q <= 'h0;
 fgallag0x00000_22_q <= 'h0;
 fgallag0x00000_23_q <= 'h0;
 fgallag0x00000_24_q <= 'h0;
 fgallag0x00000_25_q <= 'h0;
 fgallag0x00000_26_q <= 'h0;
 fgallag0x00000_27_q <= 'h0;
 fgallag0x00000_28_q <= 'h0;
 fgallag0x00000_29_q <= 'h0;
 fgallag0x00000_30_q <= 'h0;
 fgallag0x00000_31_q <= 'h0;
 fgallag0x00000_32_q <= 'h0;
 fgallag0x00000_33_q <= 'h0;
 fgallag0x00000_34_q <= 'h0;
 fgallag0x00000_35_q <= 'h0;
 fgallag0x00000_36_q <= 'h0;
 fgallag0x00000_37_q <= 'h0;
 fgallag0x00000_38_q <= 'h0;
 fgallag0x00000_39_q <= 'h0;
 fgallag0x00000_40_q <= 'h0;
 fgallag0x00000_41_q <= 'h0;
 fgallag0x00000_42_q <= 'h0;
 fgallag0x00000_43_q <= 'h0;
 fgallag0x00000_44_q <= 'h0;
 fgallag0x00000_45_q <= 'h0;
 fgallag0x00000_46_q <= 'h0;
 fgallag0x00000_47_q <= 'h0;
 fgallag0x00000_48_q <= 'h0;
 fgallag0x00000_49_q <= 'h0;
 fgallag0x00000_50_q <= 'h0;
 fgallag0x00000_51_q <= 'h0;
 fgallag0x00000_52_q <= 'h0;
 fgallag0x00000_53_q <= 'h0;
 fgallag0x00000_54_q <= 'h0;
 fgallag0x00000_55_q <= 'h0;
 fgallag0x00000_56_q <= 'h0;
 fgallag0x00000_57_q <= 'h0;
 fgallag0x00000_58_q <= 'h0;
 fgallag0x00000_59_q <= 'h0;
 fgallag0x00000_60_q <= 'h0;
 fgallag0x00000_61_q <= 'h0;
 fgallag0x00000_62_q <= 'h0;
 fgallag0x00000_63_q <= 'h0;
 fgallag0x00000_64_q <= 'h0;
 fgallag0x00000_65_q <= 'h0;
 fgallag0x00000_66_q <= 'h0;
 fgallag0x00000_67_q <= 'h0;
 fgallag0x00000_68_q <= 'h0;
 fgallag0x00000_69_q <= 'h0;
 fgallag0x00000_70_q <= 'h0;
 fgallag0x00000_71_q <= 'h0;
 fgallag0x00000_72_q <= 'h0;
 fgallag0x00000_73_q <= 'h0;
 fgallag0x00000_74_q <= 'h0;
 fgallag0x00000_75_q <= 'h0;
 fgallag0x00000_76_q <= 'h0;
 fgallag0x00000_77_q <= 'h0;
 fgallag0x00000_78_q <= 'h0;
 fgallag0x00000_79_q <= 'h0;
 fgallag0x00000_80_q <= 'h0;
 fgallag0x00000_81_q <= 'h0;
 fgallag0x00000_82_q <= 'h0;
 fgallag0x00000_83_q <= 'h0;
 fgallag0x00000_84_q <= 'h0;
 fgallag0x00000_85_q <= 'h0;
 fgallag0x00000_86_q <= 'h0;
 fgallag0x00000_87_q <= 'h0;
 fgallag0x00000_88_q <= 'h0;
 fgallag0x00000_89_q <= 'h0;
 fgallag0x00000_90_q <= 'h0;
 fgallag0x00000_91_q <= 'h0;
 fgallag0x00000_92_q <= 'h0;
 fgallag0x00000_93_q <= 'h0;
 fgallag0x00000_94_q <= 'h0;
 fgallag0x00000_95_q <= 'h0;
 fgallag0x00000_96_q <= 'h0;
 fgallag0x00000_97_q <= 'h0;
 fgallag0x00000_98_q <= 'h0;
 fgallag0x00000_99_q <= 'h0;
 fgallag0x00000_100_q <= 'h0;
 fgallag0x00000_101_q <= 'h0;
 fgallag0x00000_102_q <= 'h0;
 fgallag0x00000_103_q <= 'h0;
 fgallag0x00000_104_q <= 'h0;
 fgallag0x00000_105_q <= 'h0;
 fgallag0x00000_106_q <= 'h0;
 fgallag0x00000_107_q <= 'h0;
 fgallag0x00000_108_q <= 'h0;
 fgallag0x00000_109_q <= 'h0;
 fgallag0x00000_110_q <= 'h0;
 fgallag0x00000_111_q <= 'h0;
 fgallag0x00000_112_q <= 'h0;
 fgallag0x00000_113_q <= 'h0;
 fgallag0x00000_114_q <= 'h0;
 fgallag0x00000_115_q <= 'h0;
 fgallag0x00000_116_q <= 'h0;
 fgallag0x00000_117_q <= 'h0;
 fgallag0x00000_118_q <= 'h0;
 fgallag0x00000_119_q <= 'h0;
 fgallag0x00000_120_q <= 'h0;
 fgallag0x00000_121_q <= 'h0;
 fgallag0x00000_122_q <= 'h0;
 fgallag0x00000_123_q <= 'h0;
 fgallag0x00000_124_q <= 'h0;
 fgallag0x00000_125_q <= 'h0;
 fgallag0x00000_126_q <= 'h0;
 fgallag0x00000_127_q <= 'h0;
 fgallag0x00000_128_q <= 'h0;
 fgallag0x00000_129_q <= 'h0;
 fgallag0x00000_130_q <= 'h0;
 fgallag0x00000_131_q <= 'h0;
 fgallag0x00000_132_q <= 'h0;
 fgallag0x00000_133_q <= 'h0;
 fgallag0x00000_134_q <= 'h0;
 fgallag0x00000_135_q <= 'h0;
 fgallag0x00000_136_q <= 'h0;
 fgallag0x00000_137_q <= 'h0;
 fgallag0x00000_138_q <= 'h0;
 fgallag0x00000_139_q <= 'h0;
 fgallag0x00000_140_q <= 'h0;
 fgallag0x00000_141_q <= 'h0;
 fgallag0x00000_142_q <= 'h0;
 fgallag0x00000_143_q <= 'h0;
 fgallag0x00000_144_q <= 'h0;
 fgallag0x00000_145_q <= 'h0;
 fgallag0x00000_146_q <= 'h0;
 fgallag0x00000_147_q <= 'h0;
 fgallag0x00000_148_q <= 'h0;
 fgallag0x00000_149_q <= 'h0;
 fgallag0x00000_150_q <= 'h0;
 fgallag0x00000_151_q <= 'h0;
 fgallag0x00000_152_q <= 'h0;
 fgallag0x00000_153_q <= 'h0;
 fgallag0x00000_154_q <= 'h0;
 fgallag0x00000_155_q <= 'h0;
 fgallag0x00000_156_q <= 'h0;
 fgallag0x00000_157_q <= 'h0;
 fgallag0x00000_158_q <= 'h0;
 fgallag0x00000_159_q <= 'h0;
 fgallag0x00000_160_q <= 'h0;
 fgallag0x00000_161_q <= 'h0;
 fgallag0x00000_162_q <= 'h0;
 fgallag0x00000_163_q <= 'h0;
 fgallag0x00000_164_q <= 'h0;
 fgallag0x00000_165_q <= 'h0;
 fgallag0x00000_166_q <= 'h0;
 fgallag0x00000_167_q <= 'h0;
 fgallag0x00000_168_q <= 'h0;
 fgallag0x00000_169_q <= 'h0;
 fgallag0x00000_170_q <= 'h0;
 fgallag0x00000_171_q <= 'h0;
 fgallag0x00000_172_q <= 'h0;
 fgallag0x00000_173_q <= 'h0;
 fgallag0x00000_174_q <= 'h0;
 fgallag0x00000_175_q <= 'h0;
 fgallag0x00000_176_q <= 'h0;
 fgallag0x00000_177_q <= 'h0;
 fgallag0x00000_178_q <= 'h0;
 fgallag0x00000_179_q <= 'h0;
 fgallag0x00000_180_q <= 'h0;
 fgallag0x00000_181_q <= 'h0;
 fgallag0x00000_182_q <= 'h0;
 fgallag0x00000_183_q <= 'h0;
 fgallag0x00000_184_q <= 'h0;
 fgallag0x00000_185_q <= 'h0;
 fgallag0x00000_186_q <= 'h0;
 fgallag0x00000_187_q <= 'h0;
 fgallag0x00000_188_q <= 'h0;
 fgallag0x00000_189_q <= 'h0;
 fgallag0x00000_190_q <= 'h0;
 fgallag0x00000_191_q <= 'h0;
 fgallag0x00000_192_q <= 'h0;
 fgallag0x00000_193_q <= 'h0;
 fgallag0x00000_194_q <= 'h0;
 fgallag0x00000_195_q <= 'h0;
 fgallag0x00000_196_q <= 'h0;
 fgallag0x00000_197_q <= 'h0;
 fgallag0x00000_198_q <= 'h0;
 fgallag0x00000_199_q <= 'h0;
 fgallag0x00000_200_q <= 'h0;
 fgallag0x00000_201_q <= 'h0;
 fgallag0x00000_202_q <= 'h0;
 fgallag0x00000_203_q <= 'h0;
 fgallag0x00000_204_q <= 'h0;
 fgallag0x00000_205_q <= 'h0;
 fgallag0x00000_206_q <= 'h0;
 fgallag0x00000_207_q <= 'h0;
 fgallag0x00000_208_q <= 'h0;
 fgallag0x00000_209_q <= 'h0;
 fgallag0x00000_210_q <= 'h0;
 fgallag0x00000_211_q <= 'h0;
 fgallag0x00000_212_q <= 'h0;
 fgallag0x00000_213_q <= 'h0;
 fgallag0x00000_214_q <= 'h0;
 fgallag0x00000_215_q <= 'h0;
 fgallag0x00000_216_q <= 'h0;
 fgallag0x00000_217_q <= 'h0;
 fgallag0x00000_218_q <= 'h0;
 fgallag0x00000_219_q <= 'h0;
 fgallag0x00000_220_q <= 'h0;
 fgallag0x00000_221_q <= 'h0;
 fgallag0x00000_222_q <= 'h0;
 fgallag0x00000_223_q <= 'h0;
 fgallag0x00000_224_q <= 'h0;
 fgallag0x00000_225_q <= 'h0;
 fgallag0x00000_226_q <= 'h0;
 fgallag0x00000_227_q <= 'h0;
 fgallag0x00000_228_q <= 'h0;
 fgallag0x00000_229_q <= 'h0;
 fgallag0x00000_230_q <= 'h0;
 fgallag0x00000_231_q <= 'h0;
 fgallag0x00000_232_q <= 'h0;
 fgallag0x00000_233_q <= 'h0;
 fgallag0x00000_234_q <= 'h0;
 fgallag0x00000_235_q <= 'h0;
 fgallag0x00000_236_q <= 'h0;
 fgallag0x00000_237_q <= 'h0;
 fgallag0x00000_238_q <= 'h0;
 fgallag0x00000_239_q <= 'h0;
 fgallag0x00000_240_q <= 'h0;
 fgallag0x00000_241_q <= 'h0;
 fgallag0x00000_242_q <= 'h0;
 fgallag0x00000_243_q <= 'h0;
 fgallag0x00000_244_q <= 'h0;
 fgallag0x00000_245_q <= 'h0;
 fgallag0x00000_246_q <= 'h0;
 fgallag0x00000_247_q <= 'h0;
 fgallag0x00000_248_q <= 'h0;
 fgallag0x00000_249_q <= 'h0;
 fgallag0x00000_250_q <= 'h0;
 fgallag0x00000_251_q <= 'h0;
 fgallag0x00000_252_q <= 'h0;
 fgallag0x00000_253_q <= 'h0;
 fgallag0x00000_254_q <= 'h0;
 fgallag0x00000_255_q <= 'h0;
 fgallag0x00000_256_q <= 'h0;
 fgallag0x00000_257_q <= 'h0;
 fgallag0x00000_258_q <= 'h0;
 fgallag0x00000_259_q <= 'h0;
 fgallag0x00000_260_q <= 'h0;
 fgallag0x00000_261_q <= 'h0;
 fgallag0x00000_262_q <= 'h0;
 fgallag0x00000_263_q <= 'h0;
 fgallag0x00000_264_q <= 'h0;
 fgallag0x00000_265_q <= 'h0;
 fgallag0x00000_266_q <= 'h0;
 fgallag0x00000_267_q <= 'h0;
 fgallag0x00000_268_q <= 'h0;
 fgallag0x00000_269_q <= 'h0;
 fgallag0x00000_270_q <= 'h0;
 fgallag0x00000_271_q <= 'h0;
 fgallag0x00000_272_q <= 'h0;
 fgallag0x00000_273_q <= 'h0;
 fgallag0x00000_274_q <= 'h0;
 fgallag0x00000_275_q <= 'h0;
 fgallag0x00000_276_q <= 'h0;
 fgallag0x00000_277_q <= 'h0;
 fgallag0x00000_278_q <= 'h0;
 fgallag0x00000_279_q <= 'h0;
 fgallag0x00000_280_q <= 'h0;
 fgallag0x00000_281_q <= 'h0;
 fgallag0x00000_282_q <= 'h0;
 fgallag0x00000_283_q <= 'h0;
 fgallag0x00000_284_q <= 'h0;
 fgallag0x00000_285_q <= 'h0;
 fgallag0x00000_286_q <= 'h0;
 fgallag0x00000_287_q <= 'h0;
 fgallag0x00000_288_q <= 'h0;
 fgallag0x00000_289_q <= 'h0;
 fgallag0x00000_290_q <= 'h0;
 fgallag0x00000_291_q <= 'h0;
 fgallag0x00000_292_q <= 'h0;
 fgallag0x00000_293_q <= 'h0;
 fgallag0x00000_294_q <= 'h0;
 fgallag0x00000_295_q <= 'h0;
 fgallag0x00000_296_q <= 'h0;
 fgallag0x00000_297_q <= 'h0;
 fgallag0x00000_298_q <= 'h0;
 fgallag0x00000_299_q <= 'h0;
 fgallag0x00000_300_q <= 'h0;
 fgallag0x00000_301_q <= 'h0;
 fgallag0x00000_302_q <= 'h0;
 fgallag0x00000_303_q <= 'h0;
 fgallag0x00000_304_q <= 'h0;
 fgallag0x00000_305_q <= 'h0;
 fgallag0x00000_306_q <= 'h0;
 fgallag0x00000_307_q <= 'h0;
 fgallag0x00000_308_q <= 'h0;
 fgallag0x00000_309_q <= 'h0;
 fgallag0x00000_310_q <= 'h0;
 fgallag0x00000_311_q <= 'h0;
 fgallag0x00000_312_q <= 'h0;
 fgallag0x00000_313_q <= 'h0;
 fgallag0x00000_314_q <= 'h0;
 fgallag0x00000_315_q <= 'h0;
 fgallag0x00000_316_q <= 'h0;
 fgallag0x00000_317_q <= 'h0;
 fgallag0x00000_318_q <= 'h0;
 fgallag0x00000_319_q <= 'h0;
 fgallag0x00000_320_q <= 'h0;
 fgallag0x00000_321_q <= 'h0;
 fgallag0x00000_322_q <= 'h0;
 fgallag0x00000_323_q <= 'h0;
 fgallag0x00000_324_q <= 'h0;
 fgallag0x00000_325_q <= 'h0;
 fgallag0x00000_326_q <= 'h0;
 fgallag0x00000_327_q <= 'h0;
 fgallag0x00000_328_q <= 'h0;
 fgallag0x00000_329_q <= 'h0;
 fgallag0x00000_330_q <= 'h0;
 fgallag0x00000_331_q <= 'h0;
 fgallag0x00000_332_q <= 'h0;
 fgallag0x00000_333_q <= 'h0;
 fgallag0x00000_334_q <= 'h0;
 fgallag0x00000_335_q <= 'h0;
 fgallag0x00000_336_q <= 'h0;
 fgallag0x00000_337_q <= 'h0;
 fgallag0x00000_338_q <= 'h0;
 fgallag0x00000_339_q <= 'h0;
 fgallag0x00000_340_q <= 'h0;
 fgallag0x00000_341_q <= 'h0;
 fgallag0x00000_342_q <= 'h0;
 fgallag0x00000_343_q <= 'h0;
 fgallag0x00000_344_q <= 'h0;
 fgallag0x00000_345_q <= 'h0;
 fgallag0x00000_346_q <= 'h0;
 fgallag0x00000_347_q <= 'h0;
 fgallag0x00000_348_q <= 'h0;
 fgallag0x00000_349_q <= 'h0;
 fgallag0x00000_350_q <= 'h0;
 fgallag0x00000_351_q <= 'h0;
 fgallag0x00000_352_q <= 'h0;
 fgallag0x00000_353_q <= 'h0;
 fgallag0x00000_354_q <= 'h0;
 fgallag0x00000_355_q <= 'h0;
 start_d_fgallag0x00000_q <= 'h0;
end
else
begin
 fgallag0x00000_0_q <= fgallag0x00000_0;
 fgallag0x00000_1_q <= fgallag0x00000_1;
 fgallag0x00000_2_q <= fgallag0x00000_2;
 fgallag0x00000_3_q <= fgallag0x00000_3;
 fgallag0x00000_4_q <= fgallag0x00000_4;
 fgallag0x00000_5_q <= fgallag0x00000_5;
 fgallag0x00000_6_q <= fgallag0x00000_6;
 fgallag0x00000_7_q <= fgallag0x00000_7;
 fgallag0x00000_8_q <= fgallag0x00000_8;
 fgallag0x00000_9_q <= fgallag0x00000_9;
 fgallag0x00000_10_q <= fgallag0x00000_10;
 fgallag0x00000_11_q <= fgallag0x00000_11;
 fgallag0x00000_12_q <= fgallag0x00000_12;
 fgallag0x00000_13_q <= fgallag0x00000_13;
 fgallag0x00000_14_q <= fgallag0x00000_14;
 fgallag0x00000_15_q <= fgallag0x00000_15;
 fgallag0x00000_16_q <= fgallag0x00000_16;
 fgallag0x00000_17_q <= fgallag0x00000_17;
 fgallag0x00000_18_q <= fgallag0x00000_18;
 fgallag0x00000_19_q <= fgallag0x00000_19;
 fgallag0x00000_20_q <= fgallag0x00000_20;
 fgallag0x00000_21_q <= fgallag0x00000_21;
 fgallag0x00000_22_q <= fgallag0x00000_22;
 fgallag0x00000_23_q <= fgallag0x00000_23;
 fgallag0x00000_24_q <= fgallag0x00000_24;
 fgallag0x00000_25_q <= fgallag0x00000_25;
 fgallag0x00000_26_q <= fgallag0x00000_26;
 fgallag0x00000_27_q <= fgallag0x00000_27;
 fgallag0x00000_28_q <= fgallag0x00000_28;
 fgallag0x00000_29_q <= fgallag0x00000_29;
 fgallag0x00000_30_q <= fgallag0x00000_30;
 fgallag0x00000_31_q <= fgallag0x00000_31;
 fgallag0x00000_32_q <= fgallag0x00000_32;
 fgallag0x00000_33_q <= fgallag0x00000_33;
 fgallag0x00000_34_q <= fgallag0x00000_34;
 fgallag0x00000_35_q <= fgallag0x00000_35;
 fgallag0x00000_36_q <= fgallag0x00000_36;
 fgallag0x00000_37_q <= fgallag0x00000_37;
 fgallag0x00000_38_q <= fgallag0x00000_38;
 fgallag0x00000_39_q <= fgallag0x00000_39;
 fgallag0x00000_40_q <= fgallag0x00000_40;
 fgallag0x00000_41_q <= fgallag0x00000_41;
 fgallag0x00000_42_q <= fgallag0x00000_42;
 fgallag0x00000_43_q <= fgallag0x00000_43;
 fgallag0x00000_44_q <= fgallag0x00000_44;
 fgallag0x00000_45_q <= fgallag0x00000_45;
 fgallag0x00000_46_q <= fgallag0x00000_46;
 fgallag0x00000_47_q <= fgallag0x00000_47;
 fgallag0x00000_48_q <= fgallag0x00000_48;
 fgallag0x00000_49_q <= fgallag0x00000_49;
 fgallag0x00000_50_q <= fgallag0x00000_50;
 fgallag0x00000_51_q <= fgallag0x00000_51;
 fgallag0x00000_52_q <= fgallag0x00000_52;
 fgallag0x00000_53_q <= fgallag0x00000_53;
 fgallag0x00000_54_q <= fgallag0x00000_54;
 fgallag0x00000_55_q <= fgallag0x00000_55;
 fgallag0x00000_56_q <= fgallag0x00000_56;
 fgallag0x00000_57_q <= fgallag0x00000_57;
 fgallag0x00000_58_q <= fgallag0x00000_58;
 fgallag0x00000_59_q <= fgallag0x00000_59;
 fgallag0x00000_60_q <= fgallag0x00000_60;
 fgallag0x00000_61_q <= fgallag0x00000_61;
 fgallag0x00000_62_q <= fgallag0x00000_62;
 fgallag0x00000_63_q <= fgallag0x00000_63;
 fgallag0x00000_64_q <= fgallag0x00000_64;
 fgallag0x00000_65_q <= fgallag0x00000_65;
 fgallag0x00000_66_q <= fgallag0x00000_66;
 fgallag0x00000_67_q <= fgallag0x00000_67;
 fgallag0x00000_68_q <= fgallag0x00000_68;
 fgallag0x00000_69_q <= fgallag0x00000_69;
 fgallag0x00000_70_q <= fgallag0x00000_70;
 fgallag0x00000_71_q <= fgallag0x00000_71;
 fgallag0x00000_72_q <= fgallag0x00000_72;
 fgallag0x00000_73_q <= fgallag0x00000_73;
 fgallag0x00000_74_q <= fgallag0x00000_74;
 fgallag0x00000_75_q <= fgallag0x00000_75;
 fgallag0x00000_76_q <= fgallag0x00000_76;
 fgallag0x00000_77_q <= fgallag0x00000_77;
 fgallag0x00000_78_q <= fgallag0x00000_78;
 fgallag0x00000_79_q <= fgallag0x00000_79;
 fgallag0x00000_80_q <= fgallag0x00000_80;
 fgallag0x00000_81_q <= fgallag0x00000_81;
 fgallag0x00000_82_q <= fgallag0x00000_82;
 fgallag0x00000_83_q <= fgallag0x00000_83;
 fgallag0x00000_84_q <= fgallag0x00000_84;
 fgallag0x00000_85_q <= fgallag0x00000_85;
 fgallag0x00000_86_q <= fgallag0x00000_86;
 fgallag0x00000_87_q <= fgallag0x00000_87;
 fgallag0x00000_88_q <= fgallag0x00000_88;
 fgallag0x00000_89_q <= fgallag0x00000_89;
 fgallag0x00000_90_q <= fgallag0x00000_90;
 fgallag0x00000_91_q <= fgallag0x00000_91;
 fgallag0x00000_92_q <= fgallag0x00000_92;
 fgallag0x00000_93_q <= fgallag0x00000_93;
 fgallag0x00000_94_q <= fgallag0x00000_94;
 fgallag0x00000_95_q <= fgallag0x00000_95;
 fgallag0x00000_96_q <= fgallag0x00000_96;
 fgallag0x00000_97_q <= fgallag0x00000_97;
 fgallag0x00000_98_q <= fgallag0x00000_98;
 fgallag0x00000_99_q <= fgallag0x00000_99;
 fgallag0x00000_100_q <= fgallag0x00000_100;
 fgallag0x00000_101_q <= fgallag0x00000_101;
 fgallag0x00000_102_q <= fgallag0x00000_102;
 fgallag0x00000_103_q <= fgallag0x00000_103;
 fgallag0x00000_104_q <= fgallag0x00000_104;
 fgallag0x00000_105_q <= fgallag0x00000_105;
 fgallag0x00000_106_q <= fgallag0x00000_106;
 fgallag0x00000_107_q <= fgallag0x00000_107;
 fgallag0x00000_108_q <= fgallag0x00000_108;
 fgallag0x00000_109_q <= fgallag0x00000_109;
 fgallag0x00000_110_q <= fgallag0x00000_110;
 fgallag0x00000_111_q <= fgallag0x00000_111;
 fgallag0x00000_112_q <= fgallag0x00000_112;
 fgallag0x00000_113_q <= fgallag0x00000_113;
 fgallag0x00000_114_q <= fgallag0x00000_114;
 fgallag0x00000_115_q <= fgallag0x00000_115;
 fgallag0x00000_116_q <= fgallag0x00000_116;
 fgallag0x00000_117_q <= fgallag0x00000_117;
 fgallag0x00000_118_q <= fgallag0x00000_118;
 fgallag0x00000_119_q <= fgallag0x00000_119;
 fgallag0x00000_120_q <= fgallag0x00000_120;
 fgallag0x00000_121_q <= fgallag0x00000_121;
 fgallag0x00000_122_q <= fgallag0x00000_122;
 fgallag0x00000_123_q <= fgallag0x00000_123;
 fgallag0x00000_124_q <= fgallag0x00000_124;
 fgallag0x00000_125_q <= fgallag0x00000_125;
 fgallag0x00000_126_q <= fgallag0x00000_126;
 fgallag0x00000_127_q <= fgallag0x00000_127;
 fgallag0x00000_128_q <= fgallag0x00000_128;
 fgallag0x00000_129_q <= fgallag0x00000_129;
 fgallag0x00000_130_q <= fgallag0x00000_130;
 fgallag0x00000_131_q <= fgallag0x00000_131;
 fgallag0x00000_132_q <= fgallag0x00000_132;
 fgallag0x00000_133_q <= fgallag0x00000_133;
 fgallag0x00000_134_q <= fgallag0x00000_134;
 fgallag0x00000_135_q <= fgallag0x00000_135;
 fgallag0x00000_136_q <= fgallag0x00000_136;
 fgallag0x00000_137_q <= fgallag0x00000_137;
 fgallag0x00000_138_q <= fgallag0x00000_138;
 fgallag0x00000_139_q <= fgallag0x00000_139;
 fgallag0x00000_140_q <= fgallag0x00000_140;
 fgallag0x00000_141_q <= fgallag0x00000_141;
 fgallag0x00000_142_q <= fgallag0x00000_142;
 fgallag0x00000_143_q <= fgallag0x00000_143;
 fgallag0x00000_144_q <= fgallag0x00000_144;
 fgallag0x00000_145_q <= fgallag0x00000_145;
 fgallag0x00000_146_q <= fgallag0x00000_146;
 fgallag0x00000_147_q <= fgallag0x00000_147;
 fgallag0x00000_148_q <= fgallag0x00000_148;
 fgallag0x00000_149_q <= fgallag0x00000_149;
 fgallag0x00000_150_q <= fgallag0x00000_150;
 fgallag0x00000_151_q <= fgallag0x00000_151;
 fgallag0x00000_152_q <= fgallag0x00000_152;
 fgallag0x00000_153_q <= fgallag0x00000_153;
 fgallag0x00000_154_q <= fgallag0x00000_154;
 fgallag0x00000_155_q <= fgallag0x00000_155;
 fgallag0x00000_156_q <= fgallag0x00000_156;
 fgallag0x00000_157_q <= fgallag0x00000_157;
 fgallag0x00000_158_q <= fgallag0x00000_158;
 fgallag0x00000_159_q <= fgallag0x00000_159;
 fgallag0x00000_160_q <= fgallag0x00000_160;
 fgallag0x00000_161_q <= fgallag0x00000_161;
 fgallag0x00000_162_q <= fgallag0x00000_162;
 fgallag0x00000_163_q <= fgallag0x00000_163;
 fgallag0x00000_164_q <= fgallag0x00000_164;
 fgallag0x00000_165_q <= fgallag0x00000_165;
 fgallag0x00000_166_q <= fgallag0x00000_166;
 fgallag0x00000_167_q <= fgallag0x00000_167;
 fgallag0x00000_168_q <= fgallag0x00000_168;
 fgallag0x00000_169_q <= fgallag0x00000_169;
 fgallag0x00000_170_q <= fgallag0x00000_170;
 fgallag0x00000_171_q <= fgallag0x00000_171;
 fgallag0x00000_172_q <= fgallag0x00000_172;
 fgallag0x00000_173_q <= fgallag0x00000_173;
 fgallag0x00000_174_q <= fgallag0x00000_174;
 fgallag0x00000_175_q <= fgallag0x00000_175;
 fgallag0x00000_176_q <= fgallag0x00000_176;
 fgallag0x00000_177_q <= fgallag0x00000_177;
 fgallag0x00000_178_q <= fgallag0x00000_178;
 fgallag0x00000_179_q <= fgallag0x00000_179;
 fgallag0x00000_180_q <= fgallag0x00000_180;
 fgallag0x00000_181_q <= fgallag0x00000_181;
 fgallag0x00000_182_q <= fgallag0x00000_182;
 fgallag0x00000_183_q <= fgallag0x00000_183;
 fgallag0x00000_184_q <= fgallag0x00000_184;
 fgallag0x00000_185_q <= fgallag0x00000_185;
 fgallag0x00000_186_q <= fgallag0x00000_186;
 fgallag0x00000_187_q <= fgallag0x00000_187;
 fgallag0x00000_188_q <= fgallag0x00000_188;
 fgallag0x00000_189_q <= fgallag0x00000_189;
 fgallag0x00000_190_q <= fgallag0x00000_190;
 fgallag0x00000_191_q <= fgallag0x00000_191;
 fgallag0x00000_192_q <= fgallag0x00000_192;
 fgallag0x00000_193_q <= fgallag0x00000_193;
 fgallag0x00000_194_q <= fgallag0x00000_194;
 fgallag0x00000_195_q <= fgallag0x00000_195;
 fgallag0x00000_196_q <= fgallag0x00000_196;
 fgallag0x00000_197_q <= fgallag0x00000_197;
 fgallag0x00000_198_q <= fgallag0x00000_198;
 fgallag0x00000_199_q <= fgallag0x00000_199;
 fgallag0x00000_200_q <= fgallag0x00000_200;
 fgallag0x00000_201_q <= fgallag0x00000_201;
 fgallag0x00000_202_q <= fgallag0x00000_202;
 fgallag0x00000_203_q <= fgallag0x00000_203;
 fgallag0x00000_204_q <= fgallag0x00000_204;
 fgallag0x00000_205_q <= fgallag0x00000_205;
 fgallag0x00000_206_q <= fgallag0x00000_206;
 fgallag0x00000_207_q <= fgallag0x00000_207;
 fgallag0x00000_208_q <= fgallag0x00000_208;
 fgallag0x00000_209_q <= fgallag0x00000_209;
 fgallag0x00000_210_q <= fgallag0x00000_210;
 fgallag0x00000_211_q <= fgallag0x00000_211;
 fgallag0x00000_212_q <= fgallag0x00000_212;
 fgallag0x00000_213_q <= fgallag0x00000_213;
 fgallag0x00000_214_q <= fgallag0x00000_214;
 fgallag0x00000_215_q <= fgallag0x00000_215;
 fgallag0x00000_216_q <= fgallag0x00000_216;
 fgallag0x00000_217_q <= fgallag0x00000_217;
 fgallag0x00000_218_q <= fgallag0x00000_218;
 fgallag0x00000_219_q <= fgallag0x00000_219;
 fgallag0x00000_220_q <= fgallag0x00000_220;
 fgallag0x00000_221_q <= fgallag0x00000_221;
 fgallag0x00000_222_q <= fgallag0x00000_222;
 fgallag0x00000_223_q <= fgallag0x00000_223;
 fgallag0x00000_224_q <= fgallag0x00000_224;
 fgallag0x00000_225_q <= fgallag0x00000_225;
 fgallag0x00000_226_q <= fgallag0x00000_226;
 fgallag0x00000_227_q <= fgallag0x00000_227;
 fgallag0x00000_228_q <= fgallag0x00000_228;
 fgallag0x00000_229_q <= fgallag0x00000_229;
 fgallag0x00000_230_q <= fgallag0x00000_230;
 fgallag0x00000_231_q <= fgallag0x00000_231;
 fgallag0x00000_232_q <= fgallag0x00000_232;
 fgallag0x00000_233_q <= fgallag0x00000_233;
 fgallag0x00000_234_q <= fgallag0x00000_234;
 fgallag0x00000_235_q <= fgallag0x00000_235;
 fgallag0x00000_236_q <= fgallag0x00000_236;
 fgallag0x00000_237_q <= fgallag0x00000_237;
 fgallag0x00000_238_q <= fgallag0x00000_238;
 fgallag0x00000_239_q <= fgallag0x00000_239;
 fgallag0x00000_240_q <= fgallag0x00000_240;
 fgallag0x00000_241_q <= fgallag0x00000_241;
 fgallag0x00000_242_q <= fgallag0x00000_242;
 fgallag0x00000_243_q <= fgallag0x00000_243;
 fgallag0x00000_244_q <= fgallag0x00000_244;
 fgallag0x00000_245_q <= fgallag0x00000_245;
 fgallag0x00000_246_q <= fgallag0x00000_246;
 fgallag0x00000_247_q <= fgallag0x00000_247;
 fgallag0x00000_248_q <= fgallag0x00000_248;
 fgallag0x00000_249_q <= fgallag0x00000_249;
 fgallag0x00000_250_q <= fgallag0x00000_250;
 fgallag0x00000_251_q <= fgallag0x00000_251;
 fgallag0x00000_252_q <= fgallag0x00000_252;
 fgallag0x00000_253_q <= fgallag0x00000_253;
 fgallag0x00000_254_q <= fgallag0x00000_254;
 fgallag0x00000_255_q <= fgallag0x00000_255;
 fgallag0x00000_256_q <= fgallag0x00000_256;
 fgallag0x00000_257_q <= fgallag0x00000_257;
 fgallag0x00000_258_q <= fgallag0x00000_258;
 fgallag0x00000_259_q <= fgallag0x00000_259;
 fgallag0x00000_260_q <= fgallag0x00000_260;
 fgallag0x00000_261_q <= fgallag0x00000_261;
 fgallag0x00000_262_q <= fgallag0x00000_262;
 fgallag0x00000_263_q <= fgallag0x00000_263;
 fgallag0x00000_264_q <= fgallag0x00000_264;
 fgallag0x00000_265_q <= fgallag0x00000_265;
 fgallag0x00000_266_q <= fgallag0x00000_266;
 fgallag0x00000_267_q <= fgallag0x00000_267;
 fgallag0x00000_268_q <= fgallag0x00000_268;
 fgallag0x00000_269_q <= fgallag0x00000_269;
 fgallag0x00000_270_q <= fgallag0x00000_270;
 fgallag0x00000_271_q <= fgallag0x00000_271;
 fgallag0x00000_272_q <= fgallag0x00000_272;
 fgallag0x00000_273_q <= fgallag0x00000_273;
 fgallag0x00000_274_q <= fgallag0x00000_274;
 fgallag0x00000_275_q <= fgallag0x00000_275;
 fgallag0x00000_276_q <= fgallag0x00000_276;
 fgallag0x00000_277_q <= fgallag0x00000_277;
 fgallag0x00000_278_q <= fgallag0x00000_278;
 fgallag0x00000_279_q <= fgallag0x00000_279;
 fgallag0x00000_280_q <= fgallag0x00000_280;
 fgallag0x00000_281_q <= fgallag0x00000_281;
 fgallag0x00000_282_q <= fgallag0x00000_282;
 fgallag0x00000_283_q <= fgallag0x00000_283;
 fgallag0x00000_284_q <= fgallag0x00000_284;
 fgallag0x00000_285_q <= fgallag0x00000_285;
 fgallag0x00000_286_q <= fgallag0x00000_286;
 fgallag0x00000_287_q <= fgallag0x00000_287;
 fgallag0x00000_288_q <= fgallag0x00000_288;
 fgallag0x00000_289_q <= fgallag0x00000_289;
 fgallag0x00000_290_q <= fgallag0x00000_290;
 fgallag0x00000_291_q <= fgallag0x00000_291;
 fgallag0x00000_292_q <= fgallag0x00000_292;
 fgallag0x00000_293_q <= fgallag0x00000_293;
 fgallag0x00000_294_q <= fgallag0x00000_294;
 fgallag0x00000_295_q <= fgallag0x00000_295;
 fgallag0x00000_296_q <= fgallag0x00000_296;
 fgallag0x00000_297_q <= fgallag0x00000_297;
 fgallag0x00000_298_q <= fgallag0x00000_298;
 fgallag0x00000_299_q <= fgallag0x00000_299;
 fgallag0x00000_300_q <= fgallag0x00000_300;
 fgallag0x00000_301_q <= fgallag0x00000_301;
 fgallag0x00000_302_q <= fgallag0x00000_302;
 fgallag0x00000_303_q <= fgallag0x00000_303;
 fgallag0x00000_304_q <= fgallag0x00000_304;
 fgallag0x00000_305_q <= fgallag0x00000_305;
 fgallag0x00000_306_q <= fgallag0x00000_306;
 fgallag0x00000_307_q <= fgallag0x00000_307;
 fgallag0x00000_308_q <= fgallag0x00000_308;
 fgallag0x00000_309_q <= fgallag0x00000_309;
 fgallag0x00000_310_q <= fgallag0x00000_310;
 fgallag0x00000_311_q <= fgallag0x00000_311;
 fgallag0x00000_312_q <= fgallag0x00000_312;
 fgallag0x00000_313_q <= fgallag0x00000_313;
 fgallag0x00000_314_q <= fgallag0x00000_314;
 fgallag0x00000_315_q <= fgallag0x00000_315;
 fgallag0x00000_316_q <= fgallag0x00000_316;
 fgallag0x00000_317_q <= fgallag0x00000_317;
 fgallag0x00000_318_q <= fgallag0x00000_318;
 fgallag0x00000_319_q <= fgallag0x00000_319;
 fgallag0x00000_320_q <= fgallag0x00000_320;
 fgallag0x00000_321_q <= fgallag0x00000_321;
 fgallag0x00000_322_q <= fgallag0x00000_322;
 fgallag0x00000_323_q <= fgallag0x00000_323;
 fgallag0x00000_324_q <= fgallag0x00000_324;
 fgallag0x00000_325_q <= fgallag0x00000_325;
 fgallag0x00000_326_q <= fgallag0x00000_326;
 fgallag0x00000_327_q <= fgallag0x00000_327;
 fgallag0x00000_328_q <= fgallag0x00000_328;
 fgallag0x00000_329_q <= fgallag0x00000_329;
 fgallag0x00000_330_q <= fgallag0x00000_330;
 fgallag0x00000_331_q <= fgallag0x00000_331;
 fgallag0x00000_332_q <= fgallag0x00000_332;
 fgallag0x00000_333_q <= fgallag0x00000_333;
 fgallag0x00000_334_q <= fgallag0x00000_334;
 fgallag0x00000_335_q <= fgallag0x00000_335;
 fgallag0x00000_336_q <= fgallag0x00000_336;
 fgallag0x00000_337_q <= fgallag0x00000_337;
 fgallag0x00000_338_q <= fgallag0x00000_338;
 fgallag0x00000_339_q <= fgallag0x00000_339;
 fgallag0x00000_340_q <= fgallag0x00000_340;
 fgallag0x00000_341_q <= fgallag0x00000_341;
 fgallag0x00000_342_q <= fgallag0x00000_342;
 fgallag0x00000_343_q <= fgallag0x00000_343;
 fgallag0x00000_344_q <= fgallag0x00000_344;
 fgallag0x00000_345_q <= fgallag0x00000_345;
 fgallag0x00000_346_q <= fgallag0x00000_346;
 fgallag0x00000_347_q <= fgallag0x00000_347;
 fgallag0x00000_348_q <= fgallag0x00000_348;
 fgallag0x00000_349_q <= fgallag0x00000_349;
 fgallag0x00000_350_q <= fgallag0x00000_350;
 fgallag0x00000_351_q <= fgallag0x00000_351;
 fgallag0x00000_352_q <= fgallag0x00000_352;
 fgallag0x00000_353_q <= fgallag0x00000_353;
 fgallag0x00000_354_q <= fgallag0x00000_354;
 fgallag0x00000_355_q <= fgallag0x00000_355;
 start_d_fgallag0x00000_q <=  start_d_fgallag0x00000;
end
