//`include "GF2_LDPC_flogtanh_0x00010_assign_inc.sv"
//always_comb begin
              I3bcb7ea9f76eac891526e809fd382eaceb4a8f0a204c5ca7f391e7ffd9b7808f['h00000] = 
          (!flogtanh_sel['h00010]) ? 
                       Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00000] : //%
                       Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00001] ;
//end
//always_comb begin // 
               I3bcb7ea9f76eac891526e809fd382eaceb4a8f0a204c5ca7f391e7ffd9b7808f['h00001] =  Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00002] ;
//end
//always_comb begin // 
               I3bcb7ea9f76eac891526e809fd382eaceb4a8f0a204c5ca7f391e7ffd9b7808f['h00002] =  Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00004] ;
//end
//always_comb begin // 
               I3bcb7ea9f76eac891526e809fd382eaceb4a8f0a204c5ca7f391e7ffd9b7808f['h00003] =  Iae34f8e78093d5bcc3db929580c94da8015f69b8c6dd2133f36668c2d4b1e0c7['h00006] ;
//end
