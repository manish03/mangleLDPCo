//`include "GF2_LDPC_fgallag_0x00010_assign_inc.sv"
//always_comb begin
              Ia5096e066539b84a69d699a447597782df45e307c461c4dec11d6ed88887b470['h00000] = 
          (!fgallag_sel['h00010]) ? 
                       I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00000] : //%
                       I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00001] ;
//end
//always_comb begin // 
               Ia5096e066539b84a69d699a447597782df45e307c461c4dec11d6ed88887b470['h00001] =  I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00002] ;
//end
//always_comb begin // 
               Ia5096e066539b84a69d699a447597782df45e307c461c4dec11d6ed88887b470['h00002] =  I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00004] ;
//end
//always_comb begin // 
               Ia5096e066539b84a69d699a447597782df45e307c461c4dec11d6ed88887b470['h00003] =  I98107a78f863405ab587091acd4c59b33ef305f66522c9abc368493558d59e6c['h00006] ;
//end
